netcdf gfs_r24_2018072300_f096 {
dimensions: 
 lat = 601; 
 lon = 701; 
variables:  
float lat(lat) ; 
   lat:long_name = "latitude" ;
   lat:units = "degrees_north" ;
   lat:standard_name = "latitude" ;
float lon(lon) ;
   lon:long_name = "longitude" ;
   lon:units = "degrees_east" ;
   lon:standard_name = "longitude" ;
float APCP_24(lat, lon) ;
   APCP_24:name = "APCP_24" ;
   APCP_24:long_name = "Total Precipitation" ;
   APCP_24:level = "A24" ;
   APCP_24:units = "kg/m^2" ;
   APCP_24:_FillValue = -9999.f ;
   APCP_24:init_time = "20180723_000000" ;
   APCP_24:init_time_ut = "1532304000.0" ;
   APCP_24:valid_time = "20180727_000000" ;
   APCP_24:valid_time_ut = "1532649600.0" ;
   APCP_24:accum_time = "240000" ;
   APCP_24:_FillValue = 65535 ;
   APCP_24:accum_time_sec = 86400 ;
 // global attributes: 
 :_NCProperties = "version=1|netcdflibversion=4.4.1.1" ;
	:FileOrigins = "GFS_HR_APCP24" ; 
	:MET_version = "V7.0" ;
	:Projection = "LatLon" ;
	:lat_ll = "0.0 degrees_north" ; 
	:lon_ll = "70.0 degrees_east" ; 
	:delta_lat = "0.10 degrees" ;
	:delta_lon = "0.10 degrees" ;
	:Nlat = "601 grid_points" ; 
	:Nlon = "701 grid_points" ; 
data:
lat = 0.0,0.1,0.2,0.3,0.4,0.5,0.6,0.7,0.8,0.90000004,1.0,1.1,1.2,1.3000001,1.4,1.5,1.6,1.7,1.8000001,1.9,2.0,2.1000001,2.2,2.3,2.4,2.5,2.6000001,2.7,2.8,2.9,3.0,3.1000001,3.2,3.3,3.4,3.5,3.6000001,3.7,3.8,3.9,4.0,4.1,4.2000003,4.3,4.4,4.5,4.6,4.7000003,4.8,4.9,5.0,5.1,5.2000003,5.3,5.4,5.5,5.6,5.7000003,5.8,5.9,6.0,6.1,6.2000003,6.3,6.4,6.5,6.6,6.7000003,6.8,6.9,7.0,7.1,7.2000003,7.3,7.4,7.5,7.6,7.7000003,7.8,7.9,8.0,8.1,8.2,8.3,8.400001,8.5,8.6,8.7,8.8,8.900001,9.0,9.1,9.2,9.3,9.400001,9.5,9.6,9.7,9.8,9.900001,10.0,10.1,10.2,10.3,10.400001,10.5,10.6,10.7,10.8,10.900001,11.0,11.1,11.2,11.3,11.400001,11.5,11.6,11.7,11.8,11.900001,12.0,12.1,12.2,12.3,12.400001,12.5,12.6,12.7,12.8,12.900001,13.0,13.1,13.2,13.3,13.400001,13.5,13.6,13.7,13.8,13.900001,14.0,14.1,14.2,14.3,14.400001,14.5,14.6,14.7,14.8,14.900001,15.0,15.1,15.2,15.3,15.400001,15.5,15.6,15.7,15.8,15.900001,16.0,16.1,16.2,16.300001,16.4,16.5,16.6,16.7,16.800001,16.9,17.0,17.1,17.2,17.300001,17.4,17.5,17.6,17.7,17.800001,17.9,18.0,18.1,18.2,18.300001,18.4,18.5,18.6,18.7,18.800001,18.9,19.0,19.1,19.2,19.300001,19.4,19.5,19.6,19.7,19.800001,19.9,20.0,20.1,20.2,20.300001,20.4,20.5,20.6,20.7,20.800001,20.9,21.0,21.1,21.2,21.300001,21.4,21.5,21.6,21.7,21.800001,21.9,22.0,22.1,22.2,22.300001,22.4,22.5,22.6,22.7,22.800001,22.9,23.0,23.1,23.2,23.300001,23.4,23.5,23.6,23.7,23.800001,23.9,24.0,24.1,24.2,24.300001,24.4,24.5,24.6,24.7,24.800001,24.9,25.0,25.1,25.2,25.300001,25.4,25.5,25.6,25.7,25.800001,25.9,26.0,26.1,26.2,26.300001,26.4,26.5,26.6,26.7,26.800001,26.9,27.0,27.1,27.2,27.300001,27.4,27.5,27.6,27.7,27.800001,27.9,28.0,28.1,28.2,28.300001,28.4,28.5,28.6,28.7,28.800001,28.9,29.0,29.1,29.2,29.300001,29.4,29.5,29.6,29.7,29.800001,29.9,30.0,30.1,30.2,30.300001,30.4,30.5,30.6,30.7,30.800001,30.9,31.0,31.1,31.2,31.300001,31.4,31.5,31.6,31.7,31.800001,31.9,32.0,32.100002,32.2,32.3,32.4,32.5,32.600002,32.7,32.8,32.9,33.0,33.100002,33.2,33.3,33.4,33.5,33.600002,33.7,33.8,33.9,34.0,34.100002,34.2,34.3,34.4,34.5,34.600002,34.7,34.8,34.9,35.0,35.100002,35.2,35.3,35.4,35.5,35.600002,35.7,35.8,35.9,36.0,36.100002,36.2,36.3,36.4,36.5,36.600002,36.7,36.8,36.9,37.0,37.100002,37.2,37.3,37.4,37.5,37.600002,37.7,37.8,37.9,38.0,38.100002,38.2,38.3,38.4,38.5,38.600002,38.7,38.8,38.9,39.0,39.100002,39.2,39.3,39.4,39.5,39.600002,39.7,39.8,39.9,40.0,40.100002,40.2,40.3,40.4,40.5,40.600002,40.7,40.8,40.9,41.0,41.100002,41.2,41.3,41.4,41.5,41.600002,41.7,41.8,41.9,42.0,42.100002,42.2,42.3,42.4,42.5,42.600002,42.7,42.8,42.9,43.0,43.100002,43.2,43.3,43.4,43.5,43.600002,43.7,43.8,43.9,44.0,44.100002,44.2,44.3,44.4,44.5,44.600002,44.7,44.8,44.9,45.0,45.100002,45.2,45.3,45.4,45.5,45.600002,45.7,45.8,45.9,46.0,46.100002,46.2,46.3,46.4,46.5,46.600002,46.7,46.8,46.9,47.0,47.100002,47.2,47.3,47.4,47.5,47.600002,47.7,47.8,47.9,48.0,48.100002,48.2,48.3,48.4,48.5,48.600002,48.7,48.8,48.9,49.0,49.100002,49.2,49.3,49.4,49.5,49.600002,49.7,49.8,49.9,50.0,50.100002,50.2,50.3,50.4,50.5,50.600002,50.7,50.8,50.9,51.0,51.100002,51.2,51.3,51.4,51.5,51.600002,51.7,51.8,51.9,52.0,52.100002,52.2,52.3,52.4,52.5,52.600002,52.7,52.8,52.9,53.0,53.100002,53.2,53.3,53.4,53.5,53.600002,53.7,53.8,53.9,54.0,54.100002,54.2,54.3,54.4,54.5,54.600002,54.7,54.8,54.9,55.0,55.100002,55.2,55.3,55.4,55.5,55.600002,55.7,55.8,55.9,56.0,56.100002,56.2,56.3,56.4,56.5,56.600002,56.7,56.8,56.9,57.0,57.100002,57.2,57.3,57.4,57.5,57.600002,57.7,57.8,57.9,58.0,58.100002,58.2,58.3,58.4,58.5,58.600002,58.7,58.8,58.9,59.0,59.100002,59.2,59.3,59.4,59.5,59.600002,59.7,59.8,59.9,60.0;
lon = 70.0,70.1,70.2,70.3,70.4,70.5,70.6,70.7,70.8,70.9,71.0,71.1,71.2,71.3,71.4,71.5,71.6,71.7,71.8,71.9,72.0,72.1,72.2,72.3,72.4,72.5,72.6,72.7,72.8,72.9,73.0,73.1,73.2,73.3,73.4,73.5,73.6,73.7,73.8,73.9,74.0,74.1,74.2,74.3,74.4,74.5,74.6,74.7,74.8,74.9,75.0,75.1,75.2,75.3,75.4,75.5,75.6,75.7,75.8,75.9,76.0,76.1,76.2,76.3,76.4,76.5,76.6,76.7,76.8,76.9,77.0,77.1,77.2,77.3,77.4,77.5,77.6,77.7,77.8,77.9,78.0,78.1,78.2,78.3,78.4,78.5,78.6,78.7,78.8,78.9,79.0,79.1,79.2,79.3,79.4,79.5,79.6,79.7,79.8,79.9,80.0,80.1,80.2,80.3,80.4,80.5,80.6,80.7,80.8,80.9,81.0,81.1,81.2,81.3,81.4,81.5,81.6,81.7,81.8,81.9,82.0,82.1,82.2,82.3,82.4,82.5,82.6,82.7,82.8,82.9,83.0,83.1,83.2,83.3,83.4,83.5,83.6,83.7,83.8,83.9,84.0,84.1,84.2,84.3,84.4,84.5,84.6,84.7,84.8,84.9,85.0,85.1,85.2,85.3,85.4,85.5,85.6,85.7,85.8,85.9,86.0,86.1,86.2,86.3,86.4,86.5,86.6,86.7,86.8,86.9,87.0,87.1,87.2,87.3,87.4,87.5,87.6,87.7,87.8,87.9,88.0,88.1,88.2,88.3,88.4,88.5,88.6,88.7,88.8,88.9,89.0,89.1,89.2,89.3,89.4,89.5,89.6,89.7,89.8,89.9,90.0,90.1,90.2,90.3,90.4,90.5,90.6,90.7,90.8,90.9,91.0,91.1,91.2,91.3,91.4,91.5,91.6,91.7,91.8,91.9,92.0,92.1,92.2,92.3,92.4,92.5,92.6,92.7,92.8,92.9,93.0,93.1,93.2,93.3,93.4,93.5,93.6,93.7,93.8,93.9,94.0,94.1,94.2,94.3,94.4,94.5,94.6,94.7,94.8,94.9,95.0,95.1,95.2,95.3,95.4,95.5,95.6,95.7,95.8,95.9,96.0,96.1,96.2,96.3,96.4,96.5,96.6,96.7,96.8,96.9,97.0,97.1,97.2,97.3,97.4,97.5,97.6,97.7,97.8,97.9,98.0,98.1,98.2,98.3,98.4,98.5,98.6,98.7,98.8,98.9,99.0,99.1,99.2,99.3,99.4,99.5,99.6,99.7,99.8,99.9,100.0,100.1,100.2,100.3,100.4,100.5,100.6,100.7,100.8,100.9,101.0,101.1,101.2,101.3,101.4,101.5,101.6,101.7,101.8,101.9,102.0,102.100006,102.2,102.3,102.4,102.5,102.600006,102.7,102.8,102.9,103.0,103.100006,103.2,103.3,103.4,103.5,103.600006,103.7,103.8,103.9,104.0,104.100006,104.2,104.3,104.4,104.5,104.600006,104.7,104.8,104.9,105.0,105.100006,105.2,105.3,105.4,105.5,105.600006,105.7,105.8,105.9,106.0,106.100006,106.2,106.3,106.4,106.5,106.600006,106.7,106.8,106.9,107.0,107.100006,107.2,107.3,107.4,107.5,107.600006,107.7,107.8,107.9,108.0,108.100006,108.2,108.3,108.4,108.5,108.600006,108.7,108.8,108.9,109.0,109.100006,109.2,109.3,109.4,109.5,109.600006,109.7,109.8,109.9,110.0,110.100006,110.2,110.3,110.4,110.5,110.600006,110.7,110.8,110.9,111.0,111.100006,111.2,111.3,111.4,111.5,111.600006,111.7,111.8,111.9,112.0,112.100006,112.2,112.3,112.4,112.5,112.600006,112.7,112.8,112.9,113.0,113.100006,113.2,113.3,113.4,113.5,113.600006,113.7,113.8,113.9,114.0,114.100006,114.2,114.3,114.4,114.5,114.600006,114.7,114.8,114.9,115.0,115.100006,115.2,115.3,115.4,115.5,115.600006,115.7,115.8,115.9,116.0,116.100006,116.2,116.3,116.4,116.5,116.600006,116.7,116.8,116.9,117.0,117.100006,117.2,117.3,117.4,117.5,117.600006,117.7,117.8,117.9,118.0,118.100006,118.2,118.3,118.4,118.5,118.600006,118.7,118.8,118.9,119.0,119.100006,119.2,119.3,119.4,119.5,119.600006,119.7,119.8,119.9,120.0,120.100006,120.2,120.3,120.4,120.5,120.600006,120.7,120.8,120.9,121.0,121.100006,121.2,121.3,121.4,121.5,121.600006,121.7,121.8,121.9,122.0,122.100006,122.2,122.3,122.4,122.5,122.600006,122.7,122.8,122.9,123.0,123.100006,123.2,123.3,123.4,123.5,123.600006,123.7,123.8,123.9,124.0,124.100006,124.2,124.3,124.4,124.5,124.600006,124.7,124.8,124.9,125.0,125.100006,125.2,125.3,125.4,125.5,125.600006,125.7,125.8,125.9,126.0,126.100006,126.2,126.3,126.4,126.5,126.600006,126.7,126.8,126.9,127.0,127.100006,127.2,127.3,127.4,127.5,127.600006,127.7,127.8,127.9,128.0,128.1,128.2,128.3,128.4,128.5,128.6,128.7,128.8,128.9,129.0,129.1,129.2,129.3,129.4,129.5,129.6,129.7,129.8,129.9,130.0,130.1,130.2,130.3,130.4,130.5,130.6,130.7,130.8,130.9,131.0,131.1,131.2,131.3,131.4,131.5,131.6,131.7,131.8,131.9,132.0,132.1,132.2,132.3,132.4,132.5,132.6,132.7,132.8,132.9,133.0,133.1,133.2,133.3,133.4,133.5,133.6,133.7,133.8,133.9,134.0,134.1,134.20001,134.3,134.4,134.5,134.6,134.70001,134.8,134.9,135.0,135.1,135.20001,135.3,135.4,135.5,135.6,135.70001,135.8,135.9,136.0,136.1,136.20001,136.3,136.4,136.5,136.6,136.70001,136.8,136.9,137.0,137.1,137.20001,137.3,137.4,137.5,137.6,137.70001,137.8,137.9,138.0,138.1,138.20001,138.3,138.4,138.5,138.6,138.70001,138.8,138.9,139.0,139.1,139.20001,139.3,139.4,139.5,139.6,139.70001,139.8,139.9,140.0;
APCP_24 = 0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,0.74964523,1.3235924,1.901444,2.475391,3.049338,3.6232853,4.911738,6.2001905,7.4886436,8.773191,10.061645,9.4018,8.738052,8.074304,7.4105554,6.7507114,7.0513506,7.348085,7.648724,7.9493628,8.250002,10.0382185,11.826434,13.610746,15.398962,17.18718,17.03881,16.88654,16.738173,16.585901,16.437534,17.651802,18.862167,20.076437,21.2868,22.50107,20.349745,18.19842,16.050997,13.899672,11.748346,10.674636,9.600925,8.52331,7.4495993,6.375889,7.2856145,8.1992445,9.112875,10.0265045,10.936231,10.951848,10.963562,10.975275,10.986988,10.998701,9.874233,8.749765,7.6252975,6.5008297,5.376362,5.8370814,6.3017054,6.7624245,7.223144,7.687768,8.437413,9.187058,9.936704,10.686349,11.435994,12.173926,12.911859,13.64979,14.387722,15.125654,15.410676,15.699601,15.988527,16.273548,16.562475,14.575133,12.587793,10.600452,8.6131115,6.6257706,6.676528,6.7233806,6.774138,6.824895,6.8756523,6.5984397,6.3251314,6.0518236,5.774611,5.5013027,6.9264097,8.351517,9.776623,11.20173,12.626837,12.825961,13.025085,13.224211,13.423335,13.626364,15.012426,16.398489,17.788456,19.174519,20.560583,23.137487,25.71049,28.287394,30.8643,33.4373,32.226936,31.012667,29.798397,28.588034,27.373764,27.026272,26.674877,26.32348,25.975988,25.624592,23.699722,21.77485,19.849981,17.92511,16.00024,15.223265,14.450192,13.673217,12.900145,12.123169,10.213917,8.300759,6.387602,4.474445,2.5612879,2.2489357,1.9365835,1.6242313,1.3118792,0.999527,1.3235924,1.6515622,1.9756275,2.2996929,2.6237583,3.474918,4.3260775,5.173333,6.0244927,6.8756523,7.5003567,8.125061,8.749765,9.37447,9.999174,11.998228,14.001186,16.00024,17.999294,19.998348,21.048632,22.098917,23.1492,24.199486,25.24977,22.563541,19.873407,17.18718,14.50095,11.810817,10.975275,10.135828,9.300286,8.460839,7.6252975,7.800996,7.9766936,8.148487,8.324185,8.499884,7.9259367,7.348085,6.774138,6.2001905,5.6262436,4.985922,4.349504,3.7130866,3.076669,2.436347,1.9873407,1.5383345,1.0893283,0.63641757,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.1639849,0.3240654,0.48805028,0.6481308,0.81211567,0.698888,0.58566034,0.47633708,0.3631094,0.24988174,0.3513962,0.44900626,0.5505207,0.6481308,0.74964523,0.60127795,0.44900626,0.30063897,0.14836729,0.0,0.3631094,0.7262188,1.0893283,1.4485333,1.8116426,2.2489357,2.6862288,3.1235218,3.5608149,3.998108,6.375889,8.749765,11.123642,13.501423,15.875299,13.025085,10.174872,7.3246584,4.474445,1.6242313,1.8389735,2.0498111,2.260649,2.475391,2.6862288,2.7018464,2.7135596,2.7252727,2.736986,2.7486992,2.612045,2.475391,2.338737,2.1981785,2.0615244,2.0107672,1.9639144,1.9131571,1.8623998,1.8116426,1.9756275,2.135708,2.2996929,2.463678,2.6237583,2.3231194,2.0263848,1.7257458,1.4251068,1.1244678,2.9868677,4.8492675,6.7116675,8.574067,10.436467,8.437413,6.4383593,4.4393053,2.436347,0.43729305,1.3235924,2.2137961,3.1000953,3.9863946,4.8765984,4.900025,4.9234514,4.950782,4.9742084,5.001539,5.4115014,5.825368,6.239235,6.649197,7.0630636,6.2860875,5.5130157,4.73604,3.9629683,3.1859922,2.5495746,1.9131571,1.2767396,0.63641757,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.22645533,0.3240654,0.42557985,0.5231899,0.62470436,0.58566034,0.5505207,0.5114767,0.47633708,0.43729305,0.43729305,0.43729305,0.43729305,0.43729305,0.43729305,1.5500476,2.6628022,3.775557,4.8883114,6.001066,4.900025,3.7989833,2.7018464,1.6008049,0.4997635,2.8267872,5.1499066,7.47693,9.80005,12.123169,10.760532,9.4018,8.039165,6.676528,5.3138914,5.5013027,5.688714,5.8761253,6.0635366,6.250948,6.688241,7.125534,7.562827,8.00012,8.437413,15.500477,22.563541,29.626604,36.685764,43.74883,38.099155,32.449486,26.799816,21.150146,15.500477,14.59856,13.700547,12.798631,11.900618,10.998701,14.848442,18.698183,22.551826,26.401567,30.251308,27.764204,25.273195,22.78609,20.298986,17.811884,23.914463,30.01314,36.111816,42.214397,48.313072,40.148968,31.988768,23.824663,15.660558,7.5003567,8.238289,8.976221,9.714153,10.44818,11.186112,9.788337,8.386656,6.98888,5.5871997,4.1894236,5.298274,6.4110284,7.523783,8.636538,9.749292,9.749292,9.749292,9.749292,9.749292,9.749292,10.350571,10.951848,11.549222,12.150499,12.751778,10.237343,7.726812,5.212377,2.7018464,0.18741131,0.38653582,0.58566034,0.78868926,0.9878138,1.1869383,1.4485333,1.7140326,1.9756275,2.2372224,2.4988174,2.8111696,3.1235218,3.435874,3.7482262,4.0605783,9.300286,14.53609,19.775797,25.0116,30.251308,26.823244,23.399082,19.974922,16.55076,13.1266,12.911859,12.70102,12.486279,12.27544,12.0606985,13.376482,14.688361,16.00024,17.31212,18.623999,14.899199,11.174399,7.4495993,3.7247996,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,1.9131571,3.3265507,4.73604,6.1494336,7.562827,8.36323,9.163632,9.964035,10.764437,11.560935,10.487225,9.413514,8.335898,7.262188,6.1884775,5.2748475,4.3612175,3.4514916,2.5378613,1.6242313,2.338737,3.049338,3.7638438,4.474445,5.1889505,5.9268827,6.66091,7.3988423,8.136774,8.874706,9.089449,9.300286,9.511124,9.725866,9.936704,9.187058,8.437413,7.687768,6.9381227,6.1884775,5.001539,3.8106966,2.6237583,1.43682,0.24988174,1.901444,3.5491016,5.2006636,6.8483214,8.499884,7.137247,5.774611,4.4119744,3.049338,1.6867018,1.9131571,2.135708,2.3621633,2.5886188,2.8111696,3.1235218,3.435874,3.7482262,4.0605783,4.376835,4.9624953,5.548156,6.13772,6.7233806,7.3129454,6.3251314,5.337318,4.349504,3.3616903,2.3738766,2.3114061,2.2489357,2.1864653,2.1239948,2.0615244,1.6632754,1.261122,0.8628729,0.46071947,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.47633708,0.57394713,0.6754616,0.77307165,0.8745861,0.737932,0.60127795,0.46071947,0.3240654,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.31235218,0.4997635,0.6871748,0.8745861,1.0619974,1.3509232,1.6359446,1.9248703,2.2137961,2.4988174,2.9634414,3.4241607,3.8887846,4.349504,4.814128,5.376362,5.938596,6.5008297,7.0630636,7.6252975,7.125534,6.6257706,6.126007,5.6262436,5.12648,4.8883114,4.650143,4.4119744,4.173806,3.9356375,0.10151446,0.12103647,0.14055848,0.16008049,0.1796025,0.19912452,0.19522011,0.19131571,0.1835069,0.1796025,0.1756981,0.1717937,0.1717937,0.1678893,0.1639849,0.1639849,0.1717937,0.1756981,0.1835069,0.19131571,0.19912452,0.1796025,0.16008049,0.14055848,0.12103647,0.10151446,0.08589685,0.07027924,0.05466163,0.039044023,0.023426414,0.023426414,0.019522011,0.015617609,0.015617609,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.1756981,0.28111696,0.38263142,0.48414588,0.58566034,0.76135844,0.93315214,1.1049459,1.2767396,1.4485333,1.8741131,2.2957885,2.717464,3.1391394,3.5608149,4.8180323,6.0791545,7.336372,8.59359,9.850807,9.284669,8.718531,8.156297,7.590158,7.0240197,7.687768,8.351517,9.01136,9.675109,10.338858,11.603884,12.872814,14.141745,15.406772,16.675701,16.261835,15.844065,15.430198,15.016331,14.59856,16.004145,17.405825,18.807507,20.209187,21.610867,20.19357,18.772366,17.351164,15.933866,14.512663,13.497519,12.482374,11.46723,10.452085,9.43694,9.753197,10.065549,10.381805,10.698062,11.014318,10.971371,10.932326,10.893282,10.8542385,10.81129,9.885946,8.960603,8.039165,7.113821,6.1884775,6.617962,7.0474463,7.47693,7.9064145,8.335898,8.933272,9.526741,10.124115,10.717585,11.311053,11.931853,12.548749,13.165645,13.78254,14.399435,14.95386,15.5082855,16.066616,16.62104,17.175465,15.141272,13.110983,11.076789,9.0465,7.012306,7.1489606,7.28171,7.4183645,7.551114,7.687768,7.621393,7.558923,7.492548,7.426173,7.363703,8.6131115,9.866425,11.119738,12.373051,13.626364,13.606842,13.583415,13.563893,13.544372,13.524849,14.645412,15.765976,16.88654,18.003199,19.123762,21.025206,22.926651,24.82419,26.725634,28.623173,28.306917,27.986755,27.666594,27.346434,27.026272,26.850574,26.674877,26.499178,26.32348,26.151686,24.36347,22.579159,20.794846,19.010534,17.226223,16.69132,16.156416,15.621513,15.086611,14.551707,12.654168,10.760532,8.866898,6.969358,5.0757227,4.2284675,3.3851168,2.541766,1.6945106,0.8511597,1.1439898,1.43682,1.7257458,2.018576,2.3114061,2.979059,3.6467118,4.3143644,4.9820175,5.64967,6.126007,6.5984397,7.0747766,7.551114,8.023546,9.784432,11.545318,13.306203,15.063184,16.82407,18.003199,19.178425,20.357553,21.536682,22.711908,21.142338,19.57277,18.003199,16.43363,14.864059,14.590752,14.317443,14.044135,13.770826,13.501423,13.360865,13.220306,13.079747,12.939189,12.798631,11.72492,10.651209,9.573594,8.499884,7.426173,6.3836975,5.3412223,4.298747,3.2562714,2.2137961,1.893635,1.5773785,1.261122,0.94096094,0.62470436,0.5309987,0.44119745,0.3474918,0.25378615,0.1639849,0.26159495,0.3631094,0.46071947,0.5622339,0.6637484,0.5700427,0.47633708,0.38653582,0.29283017,0.19912452,0.32016098,0.44119745,0.5583295,0.679366,0.80040246,0.6442264,0.48414588,0.3279698,0.1717937,0.011713207,0.3435874,0.679366,1.0112402,1.3431144,1.6749885,2.05762,2.4402514,2.822883,3.2055142,3.5881457,5.883934,8.175818,10.471607,12.767395,15.063184,12.326198,9.593117,6.8561306,4.123049,1.3860629,1.7413634,2.096664,2.4519646,2.8072653,3.1625657,2.97125,2.77603,2.5847144,2.3933985,2.1981785,2.1005683,1.999054,1.901444,1.7999294,1.698415,1.7023194,1.7062237,1.7062237,1.7101282,1.7140326,1.7999294,1.8858263,1.9756275,2.0615244,2.1513257,2.0068626,1.8663043,1.7218413,1.5812829,1.43682,3.0883822,4.743849,6.395411,8.046973,9.698535,7.9454584,6.196286,4.4432096,2.690133,0.93705654,1.639849,2.3426414,3.0454338,3.7482262,4.4510183,4.5681505,4.6852827,4.802415,4.919547,5.036679,5.364649,5.6926184,6.0205884,6.348558,6.676528,5.969831,5.263134,4.560342,3.853645,3.1508527,2.5183394,1.8897307,1.261122,0.62860876,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.26159495,0.39434463,0.5309987,0.6637484,0.80040246,0.74574083,0.6910792,0.63641757,0.58175594,0.5231899,0.5388075,0.5505207,0.5622339,0.57394713,0.58566034,1.7335546,2.8814487,4.029343,5.1772375,6.3251314,5.309987,4.2948427,3.279698,2.2645533,1.2494087,3.1977055,5.1460023,7.094299,9.0386915,10.986988,10.120211,9.253433,8.386656,7.5159745,6.649197,6.5359693,6.426646,6.3134184,6.2001905,6.086963,6.4500723,6.813182,7.1762915,7.5394006,7.898606,13.884054,19.865599,25.847143,31.828688,37.814137,34.155712,30.497286,26.838861,23.184341,19.525915,18.74894,17.971964,17.191084,16.414106,15.637131,17.44487,19.252607,21.060347,22.868084,24.675823,25.296621,25.913517,26.534317,27.155117,27.775917,30.200552,32.625187,35.04982,37.474453,39.899086,33.163994,26.4289,19.693806,12.958711,6.223617,7.08649,7.9454584,8.804427,9.663396,10.526268,9.897659,9.269051,8.644346,8.015738,7.387129,7.9064145,8.421796,8.941081,9.456462,9.975748,9.788337,9.60483,9.421323,9.2339115,9.050405,9.561881,10.069453,10.58093,11.088503,11.599979,9.319808,7.039637,4.759466,2.4792955,0.19912452,0.44900626,0.698888,0.94876975,1.1986516,1.4485333,1.5969005,1.7452679,1.893635,2.0380979,2.1864653,2.5730011,2.9556324,3.3421683,3.7287042,4.1113358,8.128965,12.146595,16.164225,20.181856,24.199486,21.493734,18.791887,16.086138,13.380386,10.674636,10.471607,10.264673,10.061645,9.854712,9.651682,10.760532,11.869383,12.978233,14.090988,15.199838,12.158309,9.120684,6.0791545,3.0415294,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,1.8584955,3.3187418,4.7789884,6.239235,7.699481,8.011833,8.320281,8.628729,8.941081,9.249529,8.39056,7.531592,6.6687193,5.8097506,4.950782,4.513489,4.0801005,3.6467118,3.2094188,2.77603,3.1664703,3.5569105,3.9434462,4.3338866,4.7243266,5.270943,5.8214636,6.36808,6.914696,7.461313,7.578445,7.6916723,7.8088045,7.9220324,8.039165,7.7892823,7.5394006,7.2856145,7.0357327,6.785851,5.4700675,4.154284,2.8345962,1.5188124,0.19912452,1.8311646,3.4593005,5.0913405,6.719476,8.351517,7.551114,6.754616,5.958118,5.1616197,4.3612175,4.041056,3.7208953,3.4007344,3.0805733,2.7643168,2.9751544,3.1859922,3.4007344,3.611572,3.8263142,4.4119744,4.9937305,5.579391,6.165051,6.7507114,5.8566036,4.958591,4.0644827,3.1703746,2.2762666,2.1981785,2.1200905,2.0420024,1.9639144,1.8858263,1.5188124,1.1517987,0.78478485,0.41777104,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.19131571,0.3240654,0.45291066,0.58175594,0.7106012,0.57394713,0.43338865,0.29283017,0.15227169,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.093705654,0.113227665,0.13665408,0.15617609,0.1756981,0.23426414,0.28892577,0.3474918,0.40605783,0.46071947,0.5192855,0.57394713,0.62860876,0.6832704,0.737932,0.62079996,0.5075723,0.39434463,0.27721256,0.1639849,0.14836729,0.13665408,0.12494087,0.113227665,0.10151446,0.37482262,0.6481308,0.92534333,1.1986516,1.475864,1.698415,1.9248703,2.1513257,2.3738766,2.6003318,3.0610514,3.5256753,3.9863946,4.4510183,4.911738,5.3841705,5.8566036,6.329036,6.801469,7.2739015,6.914696,6.5554914,6.196286,5.833177,5.473972,5.5169206,5.5559645,5.5950084,5.6340523,5.6730967,0.07418364,0.113227665,0.15617609,0.19522011,0.23426414,0.27330816,0.27721256,0.28111696,0.28111696,0.28502136,0.28892577,0.28111696,0.27721256,0.27330816,0.26940376,0.26159495,0.26549935,0.26940376,0.26940376,0.27330816,0.27330816,0.24597734,0.21864653,0.19131571,0.1639849,0.13665408,0.12103647,0.10151446,0.08589685,0.06637484,0.05075723,0.046852827,0.039044023,0.03513962,0.031235218,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.3318742,0.5114767,0.6910792,0.8706817,1.0502841,1.2689307,1.4914817,1.7101282,1.9287747,2.1513257,2.4207294,2.690133,2.959537,3.2289407,3.4983444,4.728231,5.9542136,7.1841,8.410083,9.636065,9.171441,8.702912,8.234385,7.7658563,7.3012323,8.324185,9.351044,10.373997,11.400854,12.423808,13.173453,13.919194,14.668839,15.41458,16.164225,15.480955,14.801589,14.122223,13.442857,12.763491,14.356487,15.945579,17.538574,19.13157,20.724567,20.033487,19.346313,18.655233,17.964155,17.273075,16.320402,15.363823,14.411149,13.45457,12.501896,12.216875,11.935758,11.650736,11.369619,11.088503,10.994797,10.901091,10.81129,10.717585,10.6238785,9.901564,9.175345,8.449126,7.726812,7.000593,7.3988423,7.793187,8.191436,8.589685,8.987934,9.4291315,9.866425,10.307622,10.748819,11.186112,11.685876,12.181735,12.681499,13.177358,13.673217,14.4970455,15.320874,16.140799,16.964628,17.788456,15.711315,13.634172,11.553126,9.475985,7.3988423,7.621393,7.8400397,8.058686,8.281238,8.499884,8.644346,8.78881,8.933272,9.081639,9.226103,10.303718,11.385237,12.466757,13.544372,14.625891,14.383818,14.145649,13.903577,13.665408,13.423335,14.278399,15.129559,15.980719,16.835783,17.686943,18.912924,20.138906,21.360985,22.586967,23.81295,24.386896,24.95694,25.530886,26.10093,26.674877,26.674877,26.674877,26.674877,26.674877,26.674877,25.031122,23.383465,21.739712,20.095959,18.448301,18.15547,17.858736,17.565907,17.26917,16.976341,15.098324,13.220306,11.342289,9.464272,7.5862536,6.211904,4.83365,3.455396,2.077142,0.698888,0.96048295,1.2181735,1.4797685,1.7413634,1.999054,2.4831998,2.97125,3.455396,3.9395418,4.423688,4.7516575,5.0757227,5.3997884,5.7238536,6.0518236,7.570636,9.089449,10.608261,12.130978,13.64979,14.95386,16.261835,17.565907,18.869976,20.174046,19.721136,19.268225,18.81922,18.366308,17.913397,18.206228,18.499058,18.791887,19.080814,19.373644,18.920732,18.463919,18.011007,17.554192,17.101282,15.523903,13.950429,12.373051,10.799577,9.226103,7.7775693,6.329036,4.884407,3.435874,1.9873407,1.8038338,1.6164225,1.4329157,1.2494087,1.0619974,0.9136301,0.76916724,0.62079996,0.47243267,0.3240654,0.3631094,0.39824903,0.43729305,0.47633708,0.5114767,0.44119745,0.3670138,0.29673457,0.22255093,0.14836729,0.28892577,0.42948425,0.5700427,0.7106012,0.8511597,0.6832704,0.5192855,0.3553006,0.19131571,0.023426414,0.3279698,0.62860876,0.93315214,1.2337911,1.5383345,1.8663043,2.194274,2.5183394,2.8463092,3.174279,5.388075,7.605776,9.8195715,12.033368,14.251068,11.631214,9.01136,6.3915067,3.7716527,1.1517987,1.6476578,2.1435168,2.6432803,3.1391394,3.638903,3.240654,2.8424048,2.4441557,2.0459068,1.6515622,1.5890918,1.5266213,1.4641509,1.4016805,1.33921,1.3938715,1.4485333,1.5031948,1.5578566,1.6125181,1.6242313,1.6359446,1.6515622,1.6632754,1.6749885,1.6906061,1.7062237,1.7218413,1.7335546,1.7491722,3.193801,4.6345253,6.0791545,7.519879,8.960603,7.4574084,5.9542136,4.447114,2.9439192,1.43682,1.9561055,2.4714866,2.9907722,3.506153,4.025439,4.2362766,4.4432096,4.6540475,4.8648853,5.0757227,5.3177958,5.559869,5.801942,6.044015,6.2860875,5.6535745,5.017157,4.380739,3.7482262,3.1118085,2.4910088,1.8663043,1.2455044,0.62079996,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.29673457,0.46462387,0.63641757,0.80430686,0.97610056,0.9019169,0.8316377,0.75745404,0.6832704,0.61299115,0.63641757,0.6637484,0.6871748,0.7106012,0.737932,1.9209659,3.1039999,4.283129,5.466163,6.649197,5.7199492,4.7907014,3.8614538,2.9283018,1.999054,3.5686235,5.138193,6.7116675,8.281238,9.850807,9.475985,9.105066,8.734148,8.359325,7.988407,7.57454,7.1606736,6.7507114,6.336845,5.9268827,6.211904,6.5008297,6.785851,7.0747766,7.363703,12.263727,17.167656,22.071587,26.971611,31.87554,30.20836,28.545084,26.88181,25.21463,23.551353,22.895414,22.239475,21.583536,20.931501,20.27556,20.041296,19.803127,19.568865,19.3346,19.100336,22.82904,26.55384,30.282543,34.01125,37.73605,36.48664,35.237232,33.987823,32.738415,31.489004,26.179018,20.872934,15.562947,10.256865,4.950782,5.930787,6.914696,7.898606,8.878611,9.86252,10.006983,10.151445,10.295909,10.444276,10.588739,10.510651,10.432563,10.354475,10.276386,10.198298,9.8312845,9.460366,9.089449,8.718531,8.351517,8.769287,9.190963,9.608734,10.03041,10.44818,8.402273,6.356367,4.3065557,2.260649,0.21083772,0.5114767,0.81211567,1.1127546,1.4133936,1.7140326,1.7452679,1.7765031,1.8116426,1.8428779,1.8741131,2.330928,2.7916477,3.2484627,3.7052777,4.1620927,6.9615493,9.757101,12.556558,15.35211,18.151566,16.164225,14.180789,12.193448,10.2100115,8.226576,8.027451,7.8283267,7.633106,7.433982,7.238762,8.144583,9.054309,9.96013,10.865952,11.775677,9.421323,7.066968,4.7087092,2.3543546,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,1.8077383,3.3148375,4.8219366,6.329036,7.8361354,7.656533,7.47693,7.297328,7.1177254,6.9381227,6.2938967,5.645766,5.001539,4.357313,3.7130866,3.7560349,3.7989833,3.8419318,3.8809757,3.9239242,3.9942036,4.0605783,4.126953,4.193328,4.263607,4.618908,4.9781127,5.3334136,5.6926184,6.0518236,6.067441,6.083059,6.1025805,6.1181984,6.13772,6.387602,6.6374836,6.8873653,7.137247,7.387129,5.938596,4.493967,3.0454338,1.5969005,0.14836729,1.7608855,3.3694992,4.9781127,6.590631,8.1992445,7.968885,7.734621,7.504261,7.269997,7.0357327,6.17286,5.3060827,4.4432096,3.5764325,2.7135596,2.8267872,2.9361105,3.049338,3.1625657,3.2757936,3.8575494,4.4393053,5.0210614,5.606722,6.1884775,5.3841705,4.5837684,3.7794614,2.979059,2.174752,2.0810463,1.9912452,1.8975395,1.8038338,1.7140326,1.3782539,1.0424755,0.7066968,0.3709182,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.359205,0.59346914,0.8316377,1.0659018,1.3001659,1.0463798,0.78868926,0.5349031,0.28111696,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.19131571,0.23035973,0.26940376,0.30844778,0.3513962,0.39044023,0.42948425,0.46852827,0.5114767,0.5505207,0.5583295,0.5700427,0.58175594,0.58956474,0.60127795,0.5075723,0.41386664,0.3240654,0.23035973,0.13665408,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.43729305,0.80040246,1.1635119,1.5266213,1.8858263,2.0498111,2.2137961,2.3738766,2.5378613,2.7018464,3.1625657,3.6232853,4.087909,4.548629,5.0132523,5.395884,5.7785153,6.1611466,6.5437784,6.9264097,6.703859,6.4852123,6.266566,6.044015,5.825368,6.141625,6.461786,6.7780423,7.094299,7.4105554,0.05075723,0.10932326,0.1717937,0.23035973,0.28892577,0.3513962,0.359205,0.3709182,0.37872702,0.39044023,0.39824903,0.39434463,0.38653582,0.37872702,0.3709182,0.3631094,0.359205,0.359205,0.3553006,0.3513962,0.3513962,0.31625658,0.28111696,0.24597734,0.21083772,0.1756981,0.15617609,0.13665408,0.113227665,0.093705654,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.22645533,0.48414588,0.7418364,0.9956226,1.2533131,1.5110037,1.7804074,2.0459068,2.3153105,2.5808098,2.8502135,2.9673457,3.084478,3.2016098,3.3187418,3.435874,4.6345253,5.833177,7.0318284,8.226576,9.425227,9.054309,8.683391,8.316377,7.9454584,7.57454,8.960603,10.350571,11.736633,13.1266,14.512663,14.739119,14.965574,15.195933,15.422389,15.648844,14.703979,13.759113,12.814248,11.869383,10.924518,12.708829,14.489237,16.273548,18.053955,19.838268,19.877312,19.916355,19.959305,19.998348,20.037392,19.143284,18.249176,17.351164,16.457056,15.562947,14.684457,13.802062,12.923572,12.041177,11.162686,11.018223,10.87376,10.729298,10.58093,10.436467,9.913278,9.386183,8.862993,8.335898,7.812709,8.175818,8.542832,8.905942,9.272955,9.636065,9.921086,10.206107,10.491129,10.77615,11.061172,11.4398985,11.818625,12.193448,12.572175,12.950902,14.040231,15.129559,16.218887,17.308216,18.401447,16.277452,14.153459,12.033368,9.909373,7.7892823,8.093826,8.398369,8.702912,9.007456,9.311999,9.6673,10.0226,10.377901,10.733202,11.088503,11.994324,12.90405,13.809871,14.7156925,15.625418,15.164699,14.703979,14.243259,13.786445,13.325725,13.911386,14.493141,15.078801,15.664462,16.250122,16.800642,17.351164,17.901684,18.448301,18.998821,20.466877,21.931028,23.395178,24.85933,26.32348,26.499178,26.674877,26.850574,27.026272,27.198067,25.694872,24.191677,22.684578,21.181383,19.674282,19.619621,19.56496,19.510298,19.455637,19.400974,17.538574,15.680079,13.821584,11.959184,10.100689,8.191436,6.278279,4.369026,2.4597735,0.5505207,0.77697605,1.0034313,1.2337911,1.4602464,1.6867018,1.9912452,2.2918842,2.5964274,2.8970666,3.2016098,3.3734035,3.5491016,3.7247996,3.900498,4.0761957,5.35684,6.6335793,7.914223,9.194867,10.475512,11.908427,13.341343,14.774258,16.20327,17.636185,18.303837,18.967587,19.631334,20.298986,20.962736,21.821705,22.67677,23.535736,24.3908,25.24977,24.480602,23.711435,22.938364,22.169195,21.400028,19.326792,17.24965,15.176412,13.09927,11.0260315,9.171441,7.320754,5.466163,3.6154766,1.7608855,1.7101282,1.6593709,1.6047094,1.5539521,1.4992905,1.2962615,1.0932326,0.8941081,0.6910792,0.48805028,0.46071947,0.43729305,0.41386664,0.38653582,0.3631094,0.30844778,0.25769055,0.20693332,0.15227169,0.10151446,0.26159495,0.42167544,0.58175594,0.7418364,0.9019169,0.7262188,0.5544251,0.38263142,0.21083772,0.039044023,0.30844778,0.58175594,0.8550641,1.1283722,1.4016805,1.6710842,1.9443923,2.2177005,2.4910088,2.7643168,4.8961205,7.0318284,9.167537,11.303245,13.438952,10.932326,8.4257,5.9229784,3.416352,0.9136301,1.5539521,2.194274,2.8306916,3.4710135,4.1113358,3.5100577,2.9087796,2.3035975,1.7023194,1.1010414,1.0737107,1.0502841,1.0268579,0.999527,0.97610056,1.0815194,1.1908426,1.2962615,1.4055848,1.5110037,1.4485333,1.3860629,1.3235924,1.261122,1.1986516,1.3743496,1.5461433,1.717937,1.8897307,2.0615244,3.2953155,4.5291066,5.758993,6.9927845,8.226576,6.969358,5.708236,4.4510183,3.193801,1.9365835,2.2684577,2.6042364,2.9361105,3.2679846,3.5998588,3.9044023,4.2050414,4.50568,4.8102236,5.1108627,5.270943,5.4271193,5.5832953,5.743376,5.899552,5.3334136,4.7711797,4.2050414,3.638903,3.076669,2.4597735,1.8467822,1.2298868,0.61689556,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.3318742,0.5349031,0.7418364,0.94486535,1.1517987,1.0580931,0.96829176,0.8784905,0.78868926,0.698888,0.737932,0.77307165,0.81211567,0.8511597,0.8862993,2.1044729,3.3226464,4.5408196,5.758993,6.9732623,6.1299114,5.2865605,4.4393053,3.5959544,2.7486992,3.9434462,5.134289,6.329036,7.519879,8.710721,8.835662,8.956698,9.081639,9.202676,9.323712,8.6131115,7.898606,7.1880045,6.473499,5.7628975,5.9737353,6.1884775,6.3993154,6.6140575,6.824895,10.647305,14.469715,18.292124,22.114534,25.936945,26.264914,26.592884,26.920853,27.248823,27.576794,27.04189,26.510891,25.975988,25.44499,24.91399,22.63382,20.357553,18.081287,15.801116,13.524849,20.361458,27.194162,34.03077,40.863476,47.70008,42.77663,37.849274,32.925823,27.998468,23.075018,19.194042,15.31697,11.435994,7.5550184,3.6740425,4.7789884,5.883934,6.98888,8.093826,9.198771,10.116306,11.033841,11.951375,12.86891,13.786445,13.114887,12.44333,11.771772,11.096312,10.424754,9.870329,9.315904,8.761478,8.203149,7.648724,7.9805984,8.308568,8.640442,8.968412,9.300286,7.4847393,5.6691923,3.853645,2.0380979,0.22645533,0.57394713,0.92534333,1.2767396,1.6242313,1.9756275,1.893635,1.8116426,1.7257458,1.6437533,1.5617609,2.0927596,2.6237583,3.1508527,3.6818514,4.21285,5.7902284,7.367607,8.944985,10.522364,12.099743,10.834716,9.56969,8.304664,7.039637,5.774611,5.5832953,5.395884,5.2045684,5.0132523,4.825841,5.5286336,6.2353306,6.9381227,7.6448197,8.351517,6.6804323,5.009348,3.338264,1.6710842,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,1.756981,3.310933,4.8648853,6.4188375,7.9766936,7.3051367,6.6335793,5.9659266,5.2943697,4.6267166,4.193328,3.7638438,3.3343596,2.9048753,2.475391,2.9946766,3.513962,4.0332475,4.5564375,5.0757227,4.8219366,4.564246,4.31046,4.056674,3.7989833,3.9668727,4.134762,4.3026514,4.4705405,4.6384296,4.5564375,4.478349,4.396357,4.318269,4.2362766,4.985922,5.735567,6.4891167,7.238762,7.988407,6.4110284,4.83365,3.2562714,1.678893,0.10151446,1.6906061,3.279698,4.8687897,6.461786,8.050878,8.382751,8.714626,9.0465,9.378374,9.714153,8.300759,6.89127,5.481781,4.0722914,2.6628022,2.6745155,2.6862288,2.7018464,2.7135596,2.7252727,3.3031244,3.8848803,4.466636,5.044488,5.6262436,4.9156423,4.2050414,3.49444,2.7838387,2.0732377,1.9678187,1.8584955,1.7530766,1.6437533,1.5383345,1.2337911,0.93315214,0.62860876,0.3279698,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.5270943,0.8667773,1.2064602,1.5461433,1.8858263,1.5188124,1.1478943,0.77697605,0.40605783,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.22645533,0.28502136,0.3435874,0.40605783,0.46462387,0.5231899,0.5466163,0.5700427,0.59346914,0.61689556,0.63641757,0.60127795,0.5661383,0.5309987,0.4958591,0.46071947,0.39434463,0.3240654,0.25378615,0.1835069,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.4997635,0.94876975,1.4016805,1.8506867,2.2996929,2.4012074,2.4988174,2.6003318,2.7018464,2.7994564,3.2640803,3.7247996,4.1894236,4.650143,5.1108627,5.4036927,5.6965227,5.989353,6.282183,6.575013,6.4969254,6.4149327,6.336845,6.2548523,6.1767645,6.7702336,7.363703,7.9610763,8.554545,9.151918,0.023426414,0.10541886,0.1835069,0.26549935,0.3435874,0.42557985,0.44119745,0.46071947,0.47633708,0.4958591,0.5114767,0.5036679,0.49195468,0.48414588,0.47243267,0.46071947,0.45681506,0.44900626,0.44119745,0.43338865,0.42557985,0.38263142,0.339683,0.29673457,0.25378615,0.21083772,0.19131571,0.1678893,0.14446288,0.12103647,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.30063897,0.63641757,0.96829176,1.3040704,1.639849,1.9756275,2.2918842,2.6042364,2.920493,3.2367494,3.5491016,3.513962,3.4788225,3.4436827,3.408543,3.3734035,4.5408196,5.708236,6.8756523,8.043069,9.21439,8.941081,8.667773,8.3944645,8.121157,7.8517528,9.600925,11.350098,13.09927,14.848442,16.601519,16.30869,16.015858,15.723028,15.430198,15.137367,13.927003,12.716639,11.506273,10.295909,9.089449,11.061172,13.032895,15.004618,16.976341,18.948065,19.721136,20.490303,21.25947,22.028637,22.801708,21.966167,21.130625,20.295082,19.459541,18.623999,17.148134,15.668366,14.192502,12.716639,11.23687,11.04165,10.8425255,10.6434,10.44818,10.249056,9.924991,9.600925,9.276859,8.94889,8.624825,8.956698,9.288573,9.6243515,9.956225,10.2881,10.416945,10.545791,10.67854,10.807385,10.936231,11.193921,11.4516115,11.709302,11.966993,12.224684,13.583415,14.938243,16.296974,17.655706,19.014439,16.843592,14.676648,12.509705,10.342762,8.175818,8.566258,8.956698,9.343235,9.733675,10.124115,10.690253,11.256392,11.818625,12.384764,12.950902,13.68493,14.418958,15.15689,15.890917,16.624945,15.945579,15.266212,14.586847,13.903577,13.224211,13.544372,13.860628,14.176885,14.493141,14.813302,14.688361,14.56342,14.438479,14.313539,14.188598,16.546856,18.90121,21.25947,23.61773,25.975988,26.32348,26.674877,27.026272,27.373764,27.72516,26.35862,24.995983,23.629442,22.266806,20.900265,21.083773,21.271183,21.45469,21.638197,21.82561,19.98273,18.139853,16.296974,14.454097,12.611219,10.170968,7.726812,5.2865605,2.8424048,0.39824903,0.59346914,0.78868926,0.98390937,1.1791295,1.3743496,1.4953861,1.6164225,1.7335546,1.8545911,1.9756275,1.999054,2.0263848,2.0498111,2.0732377,2.1005683,3.1391394,4.181615,5.2201858,6.2587566,7.3012323,8.859089,10.42085,11.978706,13.540467,15.098324,16.882635,18.663042,20.447355,22.231667,24.012074,25.433277,26.858383,28.279585,29.700788,31.125895,30.04047,28.955048,27.869623,26.784199,25.698776,23.125774,20.548868,17.975868,15.398962,12.825961,10.569217,8.308568,6.0518236,3.795079,1.5383345,1.6164225,1.698415,1.7765031,1.8584955,1.9365835,1.678893,1.4212024,1.1635119,0.9058213,0.6481308,0.5622339,0.47633708,0.38653582,0.30063897,0.21083772,0.1796025,0.14836729,0.113227665,0.08199245,0.05075723,0.23035973,0.40996224,0.58956474,0.76916724,0.94876975,0.76916724,0.58956474,0.40996224,0.23035973,0.05075723,0.29283017,0.5349031,0.77697605,1.0190489,1.261122,1.4797685,1.698415,1.9131571,2.1318035,2.35045,4.4041657,6.461786,8.515501,10.569217,12.626837,10.2334385,7.843944,5.45445,3.0649557,0.6754616,1.456342,2.241127,3.0220075,3.8067923,4.5876727,3.7794614,2.97125,2.1630387,1.358732,0.5505207,0.5622339,0.57394713,0.58566034,0.60127795,0.61299115,0.77307165,0.93315214,1.0932326,1.2533131,1.4133936,1.2767396,1.1361811,0.999527,0.8628729,0.7262188,1.0541886,1.3860629,1.7140326,2.0459068,2.3738766,3.39683,4.4197836,5.4427366,6.46569,7.4886436,6.477403,5.466163,4.4588275,3.4475873,2.436347,2.5847144,2.7330816,2.8814487,3.0259118,3.174279,3.5686235,3.9668727,4.3612175,4.755562,5.1499066,5.22409,5.2943697,5.368553,5.4388323,5.5130157,5.017157,4.521298,4.029343,3.533484,3.0376248,2.4285383,1.8233559,1.2142692,0.60908675,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.3631094,0.60518235,0.8433509,1.0854238,1.3235924,1.2181735,1.1088502,1.0034313,0.8941081,0.78868926,0.8394465,0.8862993,0.93705654,0.9878138,1.038571,2.2918842,3.541293,4.794606,6.0479193,7.3012323,6.5398736,5.7785153,5.0210614,4.2597027,3.4983444,4.3143644,5.1303844,5.9464045,6.75852,7.57454,8.191436,8.8083315,9.4291315,10.046027,10.662923,9.651682,8.636538,7.6252975,6.6140575,5.5989127,5.735567,5.8761253,6.012779,6.1494336,6.2860875,9.030883,11.771772,14.516567,17.257458,19.998348,22.321468,24.640682,26.959898,29.279112,31.598328,31.188366,30.778402,30.36844,29.958479,29.548515,25.230247,20.911978,16.589806,12.271536,7.9493628,17.893875,27.834484,37.778996,47.719604,57.664116,49.062717,40.46132,31.863827,23.262428,14.661031,12.209065,9.757101,7.3051367,4.853172,2.4012074,3.6271896,4.853172,6.083059,7.309041,8.538928,10.229534,11.916236,13.606842,15.297448,16.988054,15.719124,14.454097,13.185166,11.916236,10.651209,9.909373,9.171441,8.429605,7.6916723,6.949836,7.191909,7.4300776,7.6682463,7.910319,8.148487,6.5672045,4.985922,3.4007344,1.8194515,0.23816854,0.63641757,1.038571,1.43682,1.8389735,2.2372224,2.0380979,1.8428779,1.6437533,1.4485333,1.2494087,1.8506867,2.455869,3.057147,3.6584249,4.263607,4.618908,4.9781127,5.3334136,5.6926184,6.0518236,5.505207,4.958591,4.415879,3.8692627,3.3265507,3.1430438,2.959537,2.77603,2.5964274,2.4129205,2.9165885,3.416352,3.9200199,4.423688,4.9234514,3.9395418,2.9556324,1.9717231,0.98390937,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,1.7023194,3.3031244,4.9078336,6.5086384,8.113348,6.9537406,5.794133,4.630621,3.4710135,2.3114061,2.096664,1.8819219,1.6671798,1.4524376,1.2376955,2.233318,3.232845,4.2284675,5.2279944,6.223617,5.645766,5.0718184,4.493967,3.9161155,3.338264,3.3148375,3.2914112,3.2718892,3.2484627,3.2250361,3.049338,2.8697357,2.6940374,2.514435,2.338737,3.5881457,4.8375545,6.086963,7.336372,8.58578,6.8795567,5.173333,3.4632049,1.756981,0.05075723,1.620327,3.1898966,4.759466,6.329036,7.898606,8.796618,9.694631,10.592644,11.490656,12.388668,10.432563,8.476458,6.524256,4.5681505,2.612045,2.5261483,2.436347,2.35045,2.260649,2.174752,2.7526035,3.330455,3.9083066,4.4861584,5.0640097,4.4432096,3.8263142,3.2094188,2.592523,1.9756275,1.8506867,1.7296503,1.6086137,1.4836729,1.3626363,1.0932326,0.8238289,0.5544251,0.28111696,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.6949836,1.1400855,1.5851873,2.0302892,2.475391,1.9912452,1.5031948,1.0190489,0.5349031,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.30063897,0.37872702,0.46071947,0.5388075,0.62079996,0.698888,0.7066968,0.7106012,0.7145056,0.71841,0.7262188,0.6442264,0.5661383,0.48414588,0.40605783,0.3240654,0.27721256,0.23035973,0.1835069,0.13665408,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.5622339,1.1010414,1.6359446,2.174752,2.7135596,2.7486992,2.787743,2.8267872,2.8619268,2.900971,3.3616903,3.8263142,4.2870336,4.7516575,5.212377,5.4154058,5.618435,5.8214636,6.0205884,6.223617,6.2860875,6.3446536,6.4032197,6.46569,6.524256,7.3988423,8.269524,9.14411,10.0147915,10.889378,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.5231899,0.5505207,0.57394713,0.60127795,0.62470436,0.61299115,0.60127795,0.58566034,0.57394713,0.5622339,0.5505207,0.5388075,0.5231899,0.5114767,0.4997635,0.44900626,0.39824903,0.3513962,0.30063897,0.24988174,0.22645533,0.19912452,0.1756981,0.14836729,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.37482262,0.78868926,1.1986516,1.6125181,2.0263848,2.436347,2.7994564,3.1625657,3.5256753,3.8887846,4.251894,4.0605783,3.873167,3.6857557,3.4983444,3.310933,4.4510183,5.5871997,6.7233806,7.8634663,8.999647,8.823949,8.648251,8.476458,8.300759,8.125061,10.237343,12.349625,14.461906,16.574188,18.68647,17.874353,17.062239,16.250122,15.438006,14.625891,13.150026,11.674163,10.198298,8.726339,7.250475,9.413514,11.576552,13.735687,15.8987255,18.061766,19.561056,21.06425,22.563541,24.062832,25.562122,24.78905,24.012074,23.239002,22.462027,21.688955,19.611813,17.538574,15.461433,13.388195,11.311053,11.061172,10.81129,10.561408,10.311526,10.061645,9.936704,9.811763,9.686822,9.561881,9.43694,9.737579,10.0382185,10.338858,10.6355915,10.936231,10.912805,10.889378,10.862047,10.838621,10.81129,10.951848,11.088503,11.225157,11.361811,11.498465,13.1266,14.750832,16.375063,17.999294,19.623526,17.413633,15.199838,12.986042,10.77615,8.562354,9.0386915,9.511124,9.987461,10.4637985,10.936231,11.713207,12.486279,13.263254,14.036326,14.813302,15.375536,15.93777,16.500004,17.062239,17.624472,16.72646,15.824542,14.92653,14.024612,13.1266,13.173453,13.224211,13.274967,13.325725,13.376482,12.576079,11.775677,10.975275,10.174872,9.37447,12.626837,15.875299,19.123762,22.37613,25.624592,26.151686,26.674877,27.198067,27.72516,28.24835,27.026272,25.80029,24.574308,23.348326,22.126247,22.551826,22.973503,23.399082,23.824663,24.250242,22.426888,20.599627,18.77627,16.94901,15.125654,12.150499,9.175345,6.2001905,3.2250361,0.24988174,0.41386664,0.57394713,0.737932,0.9019169,1.0619974,0.999527,0.93705654,0.8745861,0.81211567,0.74964523,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.92534333,1.7257458,2.5261483,3.3265507,4.123049,5.813655,7.5003567,9.187058,10.87376,12.564366,15.461433,18.362404,21.263374,24.164345,27.061413,29.048752,31.036093,33.023434,35.010777,36.998116,35.600338,34.198658,32.800884,31.399202,30.001427,26.924759,23.851994,20.775324,17.698656,14.625891,11.963089,9.300286,6.6374836,3.9746814,1.3118792,1.5266213,1.737459,1.9482968,2.1630387,2.3738766,2.0615244,1.7491722,1.43682,1.1244678,0.81211567,0.6637484,0.5114767,0.3631094,0.21083772,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.19912452,0.39824903,0.60127795,0.80040246,0.999527,0.81211567,0.62470436,0.43729305,0.24988174,0.062470436,0.27330816,0.48805028,0.698888,0.9136301,1.1244678,1.2884527,1.4485333,1.6125181,1.7765031,1.9365835,3.912211,5.8878384,7.8634663,9.839094,11.810817,9.538455,7.262188,4.985922,2.7135596,0.43729305,1.3626363,2.2879796,3.213323,4.138666,5.0640097,4.0488653,3.0376248,2.0263848,1.0112402,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.46071947,0.6754616,0.8862993,1.1010414,1.3118792,1.1010414,0.8862993,0.6754616,0.46071947,0.24988174,0.737932,1.2259823,1.7140326,2.1981785,2.6862288,3.4983444,4.3143644,5.12648,5.938596,6.7507114,5.989353,5.22409,4.462732,3.7013733,2.9361105,2.900971,2.8619268,2.8267872,2.787743,2.7486992,3.2367494,3.7247996,4.21285,4.7009,5.1889505,5.173333,5.1616197,5.1499066,5.138193,5.12648,4.7009,4.2753205,3.8497405,3.4241607,2.998581,2.4012074,1.7999294,1.1986516,0.60127795,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.39824903,0.6754616,0.94876975,1.2259823,1.4992905,1.3743496,1.2494087,1.1244678,0.999527,0.8745861,0.93705654,0.999527,1.0619974,1.1244678,1.1869383,2.475391,3.7638438,5.0483923,6.336845,7.6252975,6.949836,6.2743745,5.5989127,4.9234514,4.251894,4.689187,5.12648,5.563773,6.001066,6.4383593,7.551114,8.663869,9.776623,10.889378,11.998228,10.686349,9.37447,8.062591,6.7507114,5.4388323,5.5013027,5.563773,5.6262436,5.688714,5.7511845,7.4144597,9.073831,10.737106,12.400381,14.063657,18.374117,22.688482,26.998941,31.313307,35.623768,35.338745,35.04982,34.760895,34.475872,34.186947,27.822771,21.4625,15.098324,8.738052,2.3738766,15.426293,28.474806,41.52722,54.575733,67.624245,55.34881,43.07727,30.797924,18.526388,6.250948,5.22409,4.2011366,3.174279,2.1513257,1.1244678,2.475391,3.8263142,5.173333,6.524256,7.8751793,10.338858,12.798631,15.262308,17.725986,20.18576,18.32336,16.46096,14.59856,12.73616,10.87376,9.948417,9.026978,8.101635,7.1762915,6.250948,6.3993154,6.551587,6.699954,6.8483214,7.000593,5.64967,4.298747,2.951728,1.6008049,0.24988174,0.698888,1.1517987,1.6008049,2.0498111,2.4988174,2.1864653,1.8741131,1.5617609,1.2494087,0.93705654,1.6125181,2.2879796,2.9634414,3.638903,4.3143644,3.4514916,2.5886188,1.7257458,0.8628729,0.0,0.1756981,0.3513962,0.5231899,0.698888,0.8745861,0.698888,0.5231899,0.3513962,0.1756981,0.0,0.30063897,0.60127795,0.9019169,1.1986516,1.4992905,1.1986516,0.9019169,0.60127795,0.30063897,0.0,0.0,0.0,0.0,0.0,0.0,1.6515622,3.2992198,4.950782,6.5984397,8.250002,6.5984397,4.950782,3.2992198,1.6515622,0.0,0.0,0.0,0.0,0.0,0.0,1.475864,2.951728,4.423688,5.899552,7.375416,6.473499,5.575486,4.6735697,3.775557,2.87364,2.6628022,2.4480603,2.2372224,2.0263848,1.8116426,1.5383345,1.261122,0.9878138,0.7106012,0.43729305,2.1864653,3.9356375,5.688714,7.437886,9.187058,7.348085,5.5130157,3.6740425,1.8389735,0.0,1.5500476,3.1000953,4.650143,6.2001905,7.7502384,9.21439,10.674636,12.138786,13.599033,15.063184,12.560462,10.061645,7.562827,5.0640097,2.5612879,2.3738766,2.1864653,1.999054,1.8116426,1.6242313,2.1981785,2.77603,3.349977,3.9239242,4.5017757,3.9746814,3.4514916,2.9243972,2.4012074,1.8741131,1.737459,1.6008049,1.4641509,1.3235924,1.1869383,0.94876975,0.7106012,0.47633708,0.23816854,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.8628729,1.4133936,1.9639144,2.5105307,3.0610514,2.463678,1.8623998,1.261122,0.6637484,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.37482262,0.47633708,0.57394713,0.6754616,0.77307165,0.8745861,0.8628729,0.8511597,0.8394465,0.8238289,0.81211567,0.6871748,0.5622339,0.43729305,0.31235218,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.62470436,1.2494087,1.8741131,2.4988174,3.1235218,3.1000953,3.076669,3.049338,3.0259118,2.998581,3.4632049,3.9239242,4.388548,4.8492675,5.3138914,5.423215,5.5364423,5.64967,5.7628975,5.8761253,6.0752497,6.2743745,6.473499,6.676528,6.8756523,8.023546,9.175345,10.323239,11.475039,12.626837,0.5505207,0.62079996,0.6949836,0.76916724,0.8394465,0.9136301,0.93315214,0.95267415,0.97219616,0.9917182,1.0112402,0.97610056,0.94096094,0.9058213,0.8706817,0.8394465,0.80040246,0.76135844,0.7262188,0.6871748,0.6481308,0.61689556,0.58566034,0.5544251,0.5192855,0.48805028,0.48805028,0.48805028,0.48805028,0.48805028,0.48805028,0.5153811,0.5427119,0.5700427,0.59737355,0.62470436,0.698888,0.77307165,0.8511597,0.92534333,0.999527,1.3860629,1.7765031,2.1630387,2.5495746,2.9361105,3.1625657,3.3890212,3.611572,3.8380275,4.0605783,3.9317331,3.802888,3.6740425,3.541293,3.4124475,4.224563,5.036679,5.8487945,6.66091,7.47693,7.348085,7.2192397,7.094299,6.9654536,6.8366084,8.675582,10.510651,12.349625,14.188598,16.023666,15.5082855,14.989,14.473619,13.954333,13.438952,12.423808,11.408664,10.393518,9.378374,8.36323,10.100689,11.838148,13.575606,15.313066,17.050524,18.655233,20.259943,21.864653,23.469362,25.074072,24.539167,24.00036,23.461554,22.926651,22.387842,20.103767,17.815788,15.531713,13.247637,10.963562,10.971371,10.983084,10.990892,11.002605,11.014318,10.569217,10.124115,9.679013,9.2339115,8.78881,9.066022,9.343235,9.620447,9.897659,10.174872,10.471607,10.764437,11.061172,11.354002,11.650736,11.803008,11.955279,12.107552,12.259823,12.412095,13.501423,14.586847,15.676175,16.761599,17.850927,16.074425,14.294017,12.517513,10.741011,8.960603,9.280765,9.600925,9.921086,10.241247,10.561408,11.424281,12.28325,13.142218,14.001186,14.864059,15.231073,15.601992,15.97291,16.343828,16.710842,16.062712,15.410676,14.762545,14.114414,13.462379,13.513136,13.563893,13.610746,13.661504,13.712261,13.021181,12.334006,11.642927,10.951848,10.260769,12.946998,15.633226,18.319456,21.00178,23.68801,24.047213,24.406418,24.765623,25.128733,25.487938,24.796858,24.101875,23.410795,22.715813,22.024733,22.161386,22.294136,22.430792,22.563541,22.700195,21.048632,19.393166,17.741604,16.090042,14.438479,11.994324,9.554072,7.1099167,4.6657605,2.2255092,2.0615244,1.901444,1.737459,1.5734742,1.4133936,1.3314011,1.2533131,1.1713207,1.0932326,1.0112402,0.8433509,0.679366,0.5114767,0.3435874,0.1756981,0.80821127,1.4407244,2.0732377,2.7057507,3.338264,4.841459,6.348558,7.8517528,9.358852,10.862047,13.55218,16.242313,18.932447,21.62258,24.312714,27.108265,29.90772,32.703274,35.50273,38.298283,36.74433,35.186474,33.628616,32.07076,30.512903,27.748587,24.98427,22.21605,19.451733,16.687416,14.063657,11.443803,8.8200445,6.196286,3.5764325,3.3460727,3.1157131,2.8853533,2.6549935,2.4246337,2.2255092,2.0263848,1.8233559,1.6242313,1.4251068,1.3235924,1.2259823,1.1244678,1.0268579,0.92534333,0.8472553,0.76916724,0.6910792,0.61689556,0.5388075,0.6949836,0.8511597,1.0112402,1.1674163,1.3235924,1.175225,1.0268579,0.8745861,0.7262188,0.57394713,0.6637484,0.74964523,0.8394465,0.92534333,1.0112402,1.475864,1.9365835,2.4012074,2.8619268,3.3265507,4.552533,5.7785153,7.008402,8.234385,9.464272,7.6409154,5.8175592,3.9942036,2.1708477,0.3513962,1.0893283,1.8311646,2.5690966,3.310933,4.0488653,3.240654,2.4285383,1.620327,0.80821127,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.39044023,0.58175594,0.76916724,0.96048295,1.1517987,1.0151446,0.8784905,0.74574083,0.60908675,0.47633708,0.8238289,1.175225,1.5266213,1.8741131,2.2255092,2.8658314,3.5100577,4.154284,4.794606,5.4388323,4.9663997,4.493967,4.0215344,3.5491016,3.076669,3.018103,2.9634414,2.9087796,2.854118,2.7994564,3.193801,3.5842414,3.978586,4.369026,4.7633705,4.845363,4.927356,5.009348,5.0913405,5.173333,4.958591,4.743849,4.5291066,4.3143644,4.0996222,3.5373883,2.9751544,2.4129205,1.8506867,1.2884527,1.2689307,1.2494087,1.2259823,1.2064602,1.1869383,1.1517987,1.1127546,1.0737107,1.038571,0.999527,0.93315214,0.8667773,0.79649806,0.7301232,0.6637484,0.8316377,0.9956226,1.1635119,1.3314011,1.4992905,1.3821584,1.2650263,1.1478943,1.0307622,0.9136301,0.92143893,0.92924774,0.93315214,0.94096094,0.94876975,2.1786566,3.408543,4.6384296,5.8683167,7.098203,7.816613,8.535024,9.253433,9.971844,10.686349,9.772718,8.859089,7.941554,7.027924,6.114294,7.2543793,8.39056,9.530646,10.670732,11.810817,11.806912,11.803008,11.799104,11.791295,11.787391,10.475512,9.163632,7.8517528,6.5359693,5.22409,6.8639393,8.503788,10.143637,11.783486,13.423335,16.976341,20.529346,24.082354,27.635359,31.188366,30.649557,30.11075,29.575848,29.037039,28.498232,23.926178,19.354122,14.782067,10.2100115,5.6379566,15.363823,25.085785,34.81165,44.537518,54.263382,44.447716,34.635952,24.82419,15.012426,5.2006636,4.478349,3.7560349,3.0337205,2.3114061,1.5890918,5.0483923,8.511597,11.974802,15.438006,18.90121,19.07691,19.248703,19.4244,19.6001,19.775797,18.32336,16.874826,15.426293,13.973856,12.525322,12.415999,12.306676,12.193448,12.084125,11.974802,11.057267,10.139732,9.2221985,8.304664,7.387129,6.141625,4.892216,3.6467118,2.397303,1.1517987,1.4133936,1.678893,1.9443923,2.2098918,2.475391,2.2762666,2.0732377,1.8741131,1.6749885,1.475864,2.077142,2.67842,3.2836022,3.8848803,4.4861584,3.5881457,2.6940374,1.796025,0.8980125,0.0,1.5110037,3.0259118,4.5369153,6.0518236,7.562827,6.0518236,4.5369153,3.0259118,1.5110037,0.0,2.4714866,4.9468775,7.4183645,9.889851,12.361338,9.889851,7.4183645,4.9468775,2.4714866,0.0,0.0,0.0,0.0,0.0,0.0,1.475864,2.951728,4.423688,5.899552,7.375416,5.899552,4.423688,2.951728,1.475864,0.0,0.39824903,0.79649806,1.1908426,1.5890918,1.9873407,2.7682211,3.5530062,4.3338866,5.1186714,5.899552,5.2006636,4.5017757,3.7989833,3.1000953,2.4012074,2.241127,2.084951,1.9287747,1.7686942,1.6125181,1.3665408,1.116659,0.8706817,0.62079996,0.37482262,2.1474214,3.9200199,5.6926184,7.465217,9.237816,7.433982,5.6262436,3.8224099,2.018576,0.21083772,1.698415,3.182088,4.6657605,6.153338,7.6370106,8.55845,9.483793,10.405232,11.326671,12.24811,10.2334385,8.218767,6.2040954,4.1894236,2.174752,2.0927596,2.0107672,1.9287747,1.8467822,1.7608855,2.2137961,2.6628022,3.1118085,3.5608149,4.0137253,3.5256753,3.0376248,2.5495746,2.0615244,1.5734742,1.4485333,1.3235924,1.1986516,1.0737107,0.94876975,0.76135844,0.5700427,0.37872702,0.19131571,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.093705654,0.1756981,0.26159495,0.3435874,0.42557985,0.92924774,1.43682,1.9404879,2.4441557,2.951728,2.377781,1.8038338,1.2337911,0.659844,0.08589685,0.14836729,0.21083772,0.27330816,0.3357786,0.39824903,0.47633708,0.5505207,0.62470436,0.698888,0.77307165,0.75745404,0.7418364,0.7223144,0.7066968,0.6871748,0.58566034,0.48414588,0.37872702,0.27721256,0.1756981,0.15227169,0.12884527,0.10932326,0.08589685,0.062470436,0.058566034,0.05075723,0.046852827,0.042948425,0.039044023,0.5388075,1.038571,1.5383345,2.0380979,2.5378613,2.592523,2.6471848,2.7018464,2.7565079,2.8111696,3.2289407,3.6467118,4.0644827,4.482254,4.900025,4.9234514,4.950782,4.9742084,5.001539,5.024966,5.2006636,5.380266,5.5559645,5.735567,5.911265,6.9615493,8.011833,9.062118,10.112402,11.162686,1.1010414,1.1439898,1.1908426,1.2337911,1.2806439,1.3235924,1.33921,1.3548276,1.3704453,1.3860629,1.4016805,1.3431144,1.2845483,1.2259823,1.1713207,1.1127546,1.0502841,0.9878138,0.92534333,0.8628729,0.80040246,0.78478485,0.76916724,0.75354964,0.7418364,0.7262188,0.74964523,0.77307165,0.80040246,0.8238289,0.8511597,0.91753453,0.98390937,1.0541886,1.1205635,1.1869383,1.2767396,1.3626363,1.4485333,1.5383345,1.6242313,1.9873407,2.35045,2.7135596,3.076669,3.435874,3.5256753,3.611572,3.7013733,3.78727,3.873167,3.802888,3.7287042,3.6584249,3.5842414,3.513962,3.998108,4.4861584,4.9742084,5.462259,5.950309,5.8683167,5.7902284,5.708236,5.630148,5.548156,7.113821,8.675582,10.237343,11.799104,13.360865,13.138313,12.915763,12.693212,12.470661,12.24811,11.693685,11.139259,10.584834,10.03041,9.475985,10.787864,12.099743,13.411622,14.723501,16.039284,17.749413,19.455637,21.165764,22.875893,24.586021,24.289286,23.988647,23.68801,23.38737,23.086731,20.591818,18.096905,15.601992,13.107079,10.612165,10.881569,11.150972,11.424281,11.693685,11.963089,11.197825,10.432563,9.6673,8.902037,8.136774,8.39056,8.648251,8.902037,9.155824,9.413514,10.0265045,10.6434,11.256392,11.873287,12.486279,12.654168,12.822057,12.989946,13.157836,13.325725,13.8762455,14.426766,14.973383,15.523903,16.074425,14.73131,13.388195,12.0489855,10.705871,9.362757,9.526741,9.690726,9.858616,10.0226,10.186585,11.131451,12.076316,13.021181,13.966047,14.9109125,15.090515,15.266212,15.445815,15.621513,15.801116,15.398962,15.000713,14.59856,14.200311,13.798158,13.848915,13.899672,13.950429,14.001186,14.051944,13.470188,12.888432,12.31058,11.728825,11.150972,13.271063,15.391153,17.511244,19.631334,21.751425,21.946646,22.141865,22.333181,22.5284,22.723621,22.563541,22.40346,22.24338,22.0833,21.923218,21.770947,21.61477,21.458595,21.306324,21.150146,19.670378,18.19061,16.710842,15.231073,13.751305,11.838148,9.928895,8.019642,6.1103897,4.2011366,3.7130866,3.2250361,2.736986,2.2489357,1.7608855,1.6632754,1.5656652,1.4680552,1.3743496,1.2767396,1.0659018,0.8550641,0.6442264,0.43338865,0.22645533,0.6910792,1.1557031,1.620327,2.084951,2.5495746,3.873167,5.196759,6.5164475,7.8400397,9.163632,11.642927,14.122223,16.601519,19.080814,21.564014,25.17168,28.775444,32.387016,35.99078,39.598446,37.884415,36.170383,34.45635,32.738415,31.02438,28.568512,26.116547,23.660677,21.20481,18.74894,16.168129,13.583415,11.002605,8.421796,5.8370814,5.165524,4.493967,3.8185053,3.1469483,2.475391,2.3855898,2.2996929,2.2137961,2.1239948,2.0380979,1.9873407,1.9365835,1.8858263,1.8389735,1.7882162,1.6437533,1.5031948,1.358732,1.2181735,1.0737107,1.1908426,1.3040704,1.4212024,1.53443,1.6515622,1.5383345,1.4251068,1.3118792,1.1986516,1.0893283,1.0502841,1.0112402,0.97610056,0.93705654,0.9019169,1.6632754,2.4246337,3.1859922,3.951255,4.7126136,5.192855,5.6730967,6.153338,6.6335793,7.113821,5.743376,4.3729305,3.0024853,1.6320401,0.26159495,0.8160201,1.3743496,1.9287747,2.4831998,3.0376248,2.4285383,1.8233559,1.2142692,0.60908675,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.31625658,0.48414588,0.6520352,0.8199245,0.9878138,0.92924774,0.8706817,0.8160201,0.75745404,0.698888,0.9136301,1.1244678,1.33921,1.5500476,1.7608855,2.233318,2.7057507,3.1781836,3.6506162,4.126953,3.9434462,3.7599394,3.5764325,3.39683,3.213323,3.1391394,3.06886,2.9946766,2.9243972,2.8502135,3.1469483,3.4436827,3.7443218,4.041056,4.337791,4.513489,4.6930914,4.8687897,5.0483923,5.22409,5.2201858,5.2162814,5.2084727,5.2045684,5.2006636,4.6735697,4.1503797,3.6232853,3.1000953,2.5769055,2.522244,2.4714866,2.416825,2.366068,2.3114061,2.2137961,2.1122816,2.0107672,1.9131571,1.8116426,1.6906061,1.5656652,1.4446288,1.3235924,1.1986516,1.261122,1.319688,1.3782539,1.4407244,1.4992905,1.3899672,1.2806439,1.1713207,1.0580931,0.94876975,0.9019169,0.8550641,0.80821127,0.76135844,0.7106012,1.8858263,3.057147,4.2284675,5.4036927,6.575013,8.683391,10.795672,12.90405,15.016331,17.124708,14.856251,12.591698,10.323239,8.054782,5.786324,6.9537406,8.121157,9.288573,10.455989,11.623405,12.927476,14.231546,15.531713,16.835783,18.135948,15.449719,12.763491,10.073358,7.387129,4.7009,6.3173227,7.9337454,9.554072,11.170495,12.786918,15.578565,18.374117,21.165764,23.957413,26.74906,25.964275,25.175587,24.386896,23.598207,22.813423,20.029583,17.245745,14.465811,11.681972,8.898132,15.3013525,21.700668,28.099983,34.4993,40.898613,33.55053,26.19854,18.850454,11.498465,4.1503797,3.7287042,3.310933,2.8892577,2.4714866,2.0498111,7.6252975,13.200784,18.77627,24.351757,29.92334,27.811058,25.698776,23.586494,21.474213,19.36193,18.32336,17.288692,16.250122,15.211552,14.176885,14.879677,15.586374,16.289165,16.995863,17.698656,15.7152195,13.731783,11.744442,9.761005,7.773665,6.629675,5.4856853,4.3416953,3.193801,2.0498111,2.1318035,2.2098918,2.2918842,2.3699722,2.4480603,2.3621633,2.2762666,2.1864653,2.1005683,2.0107672,2.541766,3.0727646,3.6037633,4.1308575,4.661856,3.7287042,2.7994564,1.8663043,0.93315214,0.0,2.8502135,5.700427,8.550641,11.400854,14.251068,11.400854,8.550641,5.700427,2.8502135,0.0,4.646239,9.288573,13.934812,18.58105,23.223385,18.58105,13.934812,9.288573,4.646239,0.0,0.0,0.0,0.0,0.0,0.0,1.3001659,2.6003318,3.900498,5.2006636,6.5008297,5.2006636,3.900498,2.6003318,1.3001659,0.0,0.79649806,1.5890918,2.3855898,3.1781836,3.9746814,4.0644827,4.154284,4.2440853,4.3338866,4.423688,3.9239242,3.4241607,2.9243972,2.4246337,1.9248703,1.8233559,1.7218413,1.6164225,1.5149081,1.4133936,1.1908426,0.97219616,0.75354964,0.5309987,0.31235218,2.1083772,3.900498,5.6965227,7.492548,9.288573,7.5159745,5.743376,3.970777,2.1981785,0.42557985,1.8467822,3.2640803,4.6852827,6.1064854,7.523783,7.9064145,8.289046,8.671678,9.054309,9.43694,7.9064145,6.375889,4.8492675,3.3187418,1.7882162,1.8116426,1.8311646,1.8545911,1.8780174,1.901444,2.2255092,2.5495746,2.87364,3.2016098,3.5256753,3.076669,2.6237583,2.174752,1.7257458,1.2767396,1.1635119,1.0502841,0.93705654,0.8238289,0.7106012,0.5700427,0.42557985,0.28502136,0.14055848,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.12884527,0.23035973,0.3318742,0.43338865,0.5388075,0.9956226,1.456342,1.9170616,2.377781,2.8385005,2.2918842,1.7491722,1.2025559,0.6559396,0.113227665,0.1756981,0.23816854,0.30063897,0.3631094,0.42557985,0.47633708,0.5231899,0.57394713,0.62470436,0.6754616,0.6520352,0.62860876,0.60908675,0.58566034,0.5622339,0.48414588,0.40215343,0.3240654,0.24207294,0.1639849,0.14055848,0.12103647,0.10151446,0.08199245,0.062470436,0.06637484,0.06637484,0.07027924,0.07418364,0.07418364,0.44900626,0.8238289,1.1986516,1.5734742,1.9482968,2.084951,2.2216048,2.3543546,2.4910088,2.6237583,2.998581,3.3694992,3.7443218,4.11524,4.4861584,4.423688,4.3612175,4.298747,4.2362766,4.173806,4.3299823,4.4861584,4.6384296,4.794606,4.950782,5.899552,6.8483214,7.800996,8.749765,9.698535,1.6515622,1.6671798,1.6867018,1.7023194,1.7218413,1.737459,1.7491722,1.756981,1.7686942,1.7765031,1.7882162,1.7062237,1.6281357,1.5461433,1.4680552,1.3860629,1.3001659,1.2142692,1.1244678,1.038571,0.94876975,0.95267415,0.95657855,0.95657855,0.96048295,0.96438736,1.0112402,1.0619974,1.1127546,1.1635119,1.2142692,1.319688,1.4290112,1.53443,1.6437533,1.7491722,1.8506867,1.9482968,2.0498111,2.1513257,2.2489357,2.5886188,2.9243972,3.2640803,3.5998588,3.9356375,3.8887846,3.8380275,3.78727,3.736513,3.6857557,3.6740425,3.6584249,3.6428072,3.6271896,3.611572,3.775557,3.9356375,4.0996222,4.263607,4.423688,4.3924527,4.3612175,4.3260775,4.2948427,4.263607,5.548156,6.8366084,8.125061,9.413514,10.698062,10.772245,10.84643,10.916709,10.990892,11.061172,10.967466,10.87376,10.77615,10.682445,10.588739,11.475039,12.361338,13.251541,14.13784,15.024139,16.839687,18.655233,20.470781,22.286327,24.101875,24.039404,23.976934,23.910559,23.84809,23.785618,21.083773,18.378021,15.672271,12.96652,10.260769,10.791768,11.322766,11.8537655,12.380859,12.911859,11.826434,10.741011,9.655587,8.574067,7.4886436,7.719003,7.9532676,8.183627,8.4178915,8.648251,9.585307,10.518459,11.455516,12.388668,13.325725,13.509232,13.688834,13.872341,14.055848,14.239355,14.251068,14.262781,14.274494,14.286208,14.301826,13.392099,12.486279,11.576552,10.670732,9.761005,9.772718,9.784432,9.792241,9.803954,9.811763,10.8425255,11.873287,12.90405,13.930907,14.96167,14.946052,14.934339,14.918721,14.903104,14.8874855,14.739119,14.586847,14.438479,14.286208,14.13784,14.188598,14.239355,14.286208,14.336966,14.387722,13.919194,13.446761,12.978233,12.5058,12.037272,13.591225,15.14908,16.703033,18.256985,19.810938,19.842173,19.873407,19.900738,19.931974,19.96321,20.334127,20.70895,21.079868,21.450787,21.82561,21.380507,20.935406,20.490303,20.0452,19.6001,18.292124,16.98415,15.676175,14.3682,13.06413,11.685876,10.307622,8.929368,7.551114,6.1767645,5.3607445,4.548629,3.736513,2.9243972,2.1122816,1.999054,1.8819219,1.7686942,1.6515622,1.5383345,1.2845483,1.0307622,0.78088045,0.5270943,0.27330816,0.57394713,0.8706817,1.1674163,1.4641509,1.7608855,2.900971,4.041056,5.181142,6.321227,7.461313,9.733675,12.002132,14.274494,16.542952,18.81141,23.231194,27.647072,32.066856,36.482735,40.898613,39.028404,37.154293,35.284084,33.40997,31.535856,29.39234,27.248823,25.101402,22.957886,20.81437,18.268698,15.726933,13.185166,10.6434,8.101635,6.984976,5.8683167,4.755562,3.638903,2.5261483,2.5495746,2.5769055,2.6003318,2.6237583,2.6510892,2.6510892,2.6510892,2.6510892,2.6510892,2.6510892,2.4441557,2.233318,2.0263848,1.8194515,1.6125181,1.6867018,1.756981,1.8311646,1.901444,1.9756275,1.901444,1.8233559,1.7491722,1.6749885,1.6008049,1.43682,1.2767396,1.1127546,0.94876975,0.78868926,1.8506867,2.912684,3.9746814,5.036679,6.098676,5.833177,5.563773,5.298274,5.02887,4.7633705,3.8458362,2.9283018,2.0107672,1.0932326,0.1756981,0.5466163,0.9136301,1.2845483,1.6554666,2.0263848,1.620327,1.2142692,0.80821127,0.40605783,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.24597734,0.39044023,0.5349031,0.679366,0.8238289,0.8433509,0.8667773,0.8862993,0.9058213,0.92534333,0.999527,1.0737107,1.1517987,1.2259823,1.3001659,1.6008049,1.9053483,2.2059872,2.5105307,2.8111696,2.920493,3.0259118,3.135235,3.240654,3.349977,3.260176,3.1703746,3.0805733,2.9907722,2.900971,3.1039999,3.3031244,3.506153,3.7091823,3.912211,4.185519,4.4588275,4.728231,5.001539,5.2748475,5.481781,5.6848097,5.891743,6.094772,6.3017054,5.813655,5.3256044,4.8375545,4.349504,3.8614538,3.775557,3.6935644,3.6076677,3.521771,3.435874,3.2757936,3.1118085,2.951728,2.787743,2.6237583,2.4480603,2.2684577,2.0927596,1.9131571,1.737459,1.6906061,1.6437533,1.5969005,1.5461433,1.4992905,1.397776,1.2962615,1.1908426,1.0893283,0.9878138,0.8862993,0.78088045,0.679366,0.57785153,0.47633708,1.5890918,2.7057507,3.8185053,4.9351645,6.0518236,9.554072,13.056321,16.55857,20.06082,23.563068,19.943687,16.324306,12.70102,9.081639,5.462259,6.657006,7.8517528,9.0465,10.241247,11.435994,14.048039,16.65618,19.268225,21.876366,24.48841,20.423927,16.36335,12.298867,8.238289,4.173806,5.7707067,7.363703,8.960603,10.553599,12.150499,14.180789,16.214983,18.249176,20.279465,22.31366,21.275087,20.236517,19.20185,18.163279,17.124708,16.13299,15.141272,14.145649,13.153932,12.162213,15.238882,18.311647,21.388315,24.46108,27.537748,22.649437,17.761126,12.8767185,7.988407,3.1000953,2.9829633,2.8658314,2.7486992,2.631567,2.514435,10.202203,17.886066,25.573835,33.261604,40.94937,36.54911,32.14885,27.748587,23.348326,18.948065,18.32336,17.698656,17.073952,16.449247,15.824542,17.343355,18.866072,20.384884,21.903696,23.426414,20.37317,17.31993,14.2666855,11.213444,8.164105,7.1216297,6.0791545,5.036679,3.9942036,2.951728,2.8463092,2.7408905,2.6354716,2.5300527,2.4246337,2.4480603,2.475391,2.4988174,2.5261483,2.5495746,3.0063896,3.4632049,3.9239242,4.380739,4.8375545,3.8692627,2.900971,1.9365835,0.96829176,0.0,4.1894236,8.374943,12.564366,16.749886,20.93931,16.749886,12.564366,8.374943,4.185519,0.0,6.817086,13.634172,20.45126,27.268345,34.089336,27.268345,20.45126,13.634172,6.817086,0.0,0.0,0.0,0.0,0.0,0.0,1.1244678,2.2489357,3.3734035,4.5017757,5.6262436,4.5017757,3.3734035,2.2489357,1.1244678,0.0,1.1908426,2.3855898,3.5764325,4.7711797,5.9620223,5.3607445,4.759466,4.154284,3.5530062,2.951728,2.6510892,2.35045,2.0498111,1.7491722,1.4485333,1.4016805,1.3548276,1.3079748,1.261122,1.2142692,1.0190489,0.8277333,0.63641757,0.44119745,0.24988174,2.069333,3.8848803,5.704332,7.519879,9.339331,7.5979667,5.8566036,4.1191444,2.377781,0.63641757,1.9912452,3.3460727,4.7009,6.055728,7.4105554,7.2543793,7.098203,6.9381227,6.7819467,6.6257706,5.579391,4.5369153,3.4905357,2.4441557,1.4016805,1.5266213,1.6554666,1.7843118,1.9092526,2.0380979,2.2372224,2.436347,2.639376,2.8385005,3.0376248,2.6237583,2.2137961,1.7999294,1.3860629,0.97610056,0.8745861,0.77307165,0.6754616,0.57394713,0.47633708,0.37872702,0.28502136,0.19131571,0.093705654,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.16008049,0.28111696,0.40605783,0.5270943,0.6481308,1.0659018,1.4797685,1.893635,2.3114061,2.7252727,2.2059872,1.6906061,1.1713207,0.6559396,0.13665408,0.19912452,0.26159495,0.3240654,0.38653582,0.44900626,0.47633708,0.4997635,0.5231899,0.5505207,0.57394713,0.5466163,0.5192855,0.49195468,0.46462387,0.43729305,0.37872702,0.3240654,0.26549935,0.20693332,0.14836729,0.13274968,0.113227665,0.09761006,0.078088045,0.062470436,0.07418364,0.08199245,0.093705654,0.10151446,0.113227665,0.3631094,0.61299115,0.8628729,1.1127546,1.3626363,1.5773785,1.7921207,2.0068626,2.2216048,2.436347,2.7643168,3.0922866,3.4202564,3.7482262,4.0761957,3.9239242,3.775557,3.6232853,3.474918,3.3265507,3.4593005,3.5881457,3.7208953,3.853645,3.9863946,4.8375545,5.688714,6.5359693,7.387129,8.238289,2.1981785,2.1903696,2.1786566,2.1708477,2.1591344,2.1513257,2.15523,2.1591344,2.1669433,2.1708477,2.174752,2.0732377,1.9717231,1.8663043,1.7647898,1.6632754,1.5500476,1.43682,1.3235924,1.2142692,1.1010414,1.1205635,1.1400855,1.1596074,1.1791295,1.1986516,1.2767396,1.3509232,1.4251068,1.4992905,1.5734742,1.7218413,1.8702087,2.018576,2.1669433,2.3114061,2.4246337,2.5378613,2.6510892,2.7643168,2.87364,3.1859922,3.4983444,3.8106966,4.126953,4.4393053,4.251894,4.0605783,3.873167,3.6857557,3.4983444,3.541293,3.5842414,3.6271896,3.6701381,3.7130866,3.5491016,3.3890212,3.2250361,3.0610514,2.900971,2.9165885,2.9283018,2.9439192,2.959537,2.9751544,3.9863946,5.001539,6.012779,7.0240197,8.039165,8.406178,8.773191,9.140205,9.507219,9.874233,10.241247,10.604357,10.971371,11.334479,11.701493,12.162213,12.626837,13.087557,13.548276,14.012899,15.933866,17.850927,19.771893,21.69286,23.613825,23.785618,23.961317,24.137014,24.312714,24.48841,21.571823,18.659138,15.74255,12.825961,9.913278,10.701966,11.490656,12.28325,13.0719385,13.860628,12.458947,11.053363,9.647778,8.242193,6.8366084,7.0474463,7.2582836,7.4691215,7.676055,7.8868923,9.14411,10.397423,11.650736,12.907954,14.161267,14.360392,14.555612,14.754736,14.95386,15.14908,14.625891,14.098797,13.575606,13.048512,12.525322,12.05289,11.580457,11.108025,10.6355915,10.163159,10.018696,9.874233,9.725866,9.581403,9.43694,10.553599,11.666354,12.783013,13.895767,15.012426,14.805493,14.59856,14.391626,14.180789,13.973856,14.07537,14.176885,14.274494,14.376009,14.473619,14.524376,14.575133,14.625891,14.676648,14.723501,14.364296,14.005091,13.645885,13.286681,12.923572,13.91529,14.903104,15.894821,16.88654,17.874353,17.741604,17.60495,17.468296,17.335546,17.198893,18.104713,19.010534,19.916355,20.818274,21.724094,20.990067,20.256039,19.518106,18.784079,18.05005,16.91387,15.781594,14.645412,13.509232,12.376955,11.5297,10.686349,9.839094,8.995743,8.148487,7.012306,5.8761253,4.73604,3.5998588,2.463678,2.330928,2.1981785,2.0654287,1.9326792,1.7999294,1.5031948,1.2103647,0.9136301,0.62079996,0.3240654,0.45681506,0.58566034,0.7145056,0.8433509,0.97610056,1.9326792,2.8892577,3.8458362,4.806319,5.7628975,7.824422,9.882042,11.943566,14.001186,16.062712,21.290705,26.5187,31.746695,36.970783,42.19878,40.16849,38.138203,36.111816,34.081528,32.05124,30.21617,28.3811,26.54603,24.710962,22.875893,20.37317,17.87045,15.367727,12.8650055,10.362284,8.804427,7.2465706,5.688714,4.1308575,2.5769055,2.7135596,2.8502135,2.9868677,3.1235218,3.2640803,3.310933,3.3616903,3.4124475,3.4632049,3.513962,3.240654,2.9673457,2.6940374,2.4207294,2.1513257,2.1786566,2.2098918,2.241127,2.2684577,2.2996929,2.260649,2.2255092,2.1864653,2.1513257,2.1122816,1.8233559,1.5383345,1.2494087,0.96438736,0.6754616,2.0380979,3.4007344,4.7633705,6.126007,7.4886436,6.473499,5.4583545,4.4432096,3.4280653,2.4129205,1.9482968,1.4836729,1.0190489,0.5544251,0.08589685,0.27330816,0.45681506,0.6442264,0.8277333,1.0112402,0.80821127,0.60908675,0.40605783,0.20302892,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.1717937,0.29673457,0.41777104,0.5388075,0.6637484,0.76135844,0.8589685,0.95657855,1.0541886,1.1517987,1.0893283,1.0268579,0.96438736,0.9019169,0.8394465,0.96829176,1.1010414,1.2337911,1.3665408,1.4992905,1.8975395,2.2957885,2.6940374,3.0883822,3.4866312,3.3812122,3.2718892,3.1664703,3.057147,2.951728,3.057147,3.1664703,3.2718892,3.3812122,3.4866312,3.853645,4.220659,4.591577,4.958591,5.3256044,5.7394714,6.153338,6.571109,6.984976,7.3988423,6.949836,6.5008297,6.0518236,5.5989127,5.1499066,5.0327744,4.9156423,4.7985106,4.6813784,4.564246,4.337791,4.1113358,3.8887846,3.6623292,3.435874,3.2055142,2.97125,2.7408905,2.5066261,2.2762666,2.1200905,1.9639144,1.8116426,1.6554666,1.4992905,1.4055848,1.3118792,1.2142692,1.1205635,1.0268579,0.8667773,0.7106012,0.5544251,0.39434463,0.23816854,1.2962615,2.3543546,3.408543,4.466636,5.5247293,10.42085,15.313066,20.209187,25.105307,30.001427,25.027218,20.056915,15.0827055,10.108498,5.138193,6.3602715,7.5823493,8.804427,10.0265045,11.248583,15.168603,19.084719,23.000834,26.920853,30.83697,25.398136,19.96321,14.524376,9.085544,3.6506162,5.22409,6.79366,8.367134,9.940608,11.514082,12.786918,14.055848,15.328683,16.601519,17.874353,16.585901,15.3013525,14.012899,12.724447,11.435994,12.236397,13.032895,13.829392,14.625891,15.426293,15.176412,14.92653,14.676648,14.426766,14.176885,11.748346,9.323712,6.899079,4.474445,2.0498111,2.233318,2.4207294,2.6042364,2.7916477,2.9751544,12.775204,22.575254,32.375305,42.175354,51.975403,45.287163,38.59892,31.910679,25.226343,18.538101,18.32336,18.112522,17.901684,17.686943,17.476105,19.810938,22.14577,24.480602,26.815435,29.150267,25.031122,20.911978,16.788929,12.6697855,8.550641,7.60968,6.6687193,5.7316628,4.7907014,3.8497405,3.5608149,3.2718892,2.979059,2.690133,2.4012074,2.5378613,2.6745155,2.8111696,2.951728,3.0883822,3.4710135,3.8575494,4.2440853,4.6267166,5.0132523,4.009821,3.0063896,2.0068626,1.0034313,0.0,5.5247293,11.0494585,16.574188,22.098917,27.623646,22.098917,16.574188,11.0494585,5.5247293,0.0,8.991838,17.979773,26.971611,35.959545,44.95138,35.959545,26.971611,17.979773,8.987934,0.0,0.0,0.0,0.0,0.0,0.0,0.94876975,1.901444,2.8502135,3.7989833,4.7516575,3.7989833,2.8502135,1.901444,0.94876975,0.0,1.5890918,3.1781836,4.7711797,6.3602715,7.9493628,6.6531014,5.3607445,4.0644827,2.7682211,1.475864,1.3743496,1.2767396,1.175225,1.0737107,0.97610056,0.98390937,0.9917182,0.9956226,1.0034313,1.0112402,0.8472553,0.6832704,0.5192855,0.3513962,0.18741131,2.0263848,3.8692627,5.708236,7.5472097,9.386183,7.6799593,5.9737353,4.263607,2.5573835,0.8511597,2.1396124,3.4280653,4.7204223,6.008875,7.3012323,6.602344,5.903456,5.2084727,4.5095844,3.8106966,3.252367,2.6940374,2.1318035,1.5734742,1.0112402,1.2455044,1.475864,1.7101282,1.9443923,2.174752,2.2489357,2.3231194,2.4012074,2.475391,2.5495746,2.174752,1.7999294,1.4251068,1.0502841,0.6754616,0.58566034,0.4997635,0.41386664,0.3240654,0.23816854,0.19131571,0.14055848,0.093705654,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.19131571,0.3357786,0.47633708,0.62079996,0.76135844,1.1322767,1.5031948,1.8741131,2.241127,2.612045,2.1239948,1.6320401,1.1439898,0.6520352,0.1639849,0.22645533,0.28892577,0.3513962,0.41386664,0.47633708,0.47633708,0.47633708,0.47633708,0.47633708,0.47633708,0.44119745,0.40996224,0.37872702,0.3435874,0.31235218,0.27721256,0.24207294,0.20693332,0.1717937,0.13665408,0.12103647,0.10932326,0.093705654,0.078088045,0.062470436,0.078088045,0.09761006,0.113227665,0.13274968,0.14836729,0.27330816,0.39824903,0.5231899,0.6481308,0.77307165,1.0698062,1.3665408,1.6593709,1.9561055,2.2489357,2.533957,2.815074,3.096191,3.3812122,3.6623292,3.4241607,3.1859922,2.951728,2.7135596,2.475391,2.5847144,2.6940374,2.803361,2.9165885,3.0259118,3.775557,4.5252023,5.2748475,6.0244927,6.774138,2.7486992,2.7135596,2.6745155,2.639376,2.6003318,2.5612879,2.5612879,2.5612879,2.5612879,2.5612879,2.5612879,2.436347,2.3114061,2.1864653,2.0615244,1.9365835,1.7999294,1.6632754,1.5266213,1.3860629,1.2494087,1.2884527,1.3235924,1.3626363,1.4016805,1.43682,1.5383345,1.6359446,1.737459,1.8389735,1.9365835,2.1239948,2.3114061,2.4988174,2.6862288,2.87364,2.998581,3.1235218,3.2484627,3.3734035,3.4983444,3.78727,4.0761957,4.3612175,4.650143,4.939069,4.6110992,4.2870336,3.9629683,3.638903,3.310933,3.4124475,3.513962,3.611572,3.7130866,3.8106966,3.3265507,2.8385005,2.35045,1.8623998,1.3743496,1.43682,1.4992905,1.5617609,1.6242313,1.6867018,2.4246337,3.1625657,3.900498,4.6384296,5.376362,6.036206,6.699954,7.363703,8.023546,8.687295,9.511124,10.338858,11.162686,11.986515,12.814248,12.849388,12.888432,12.923572,12.962616,13.001659,15.024139,17.050524,19.07691,21.09939,23.125774,23.535736,23.949604,24.36347,24.773432,25.1873,22.063778,18.936352,15.812829,12.689307,9.561881,10.612165,11.66245,12.712734,13.763018,14.813302,13.087557,11.361811,9.636065,7.914223,6.1884775,6.375889,6.5633,6.7507114,6.9381227,7.125534,8.699008,10.276386,11.849861,13.423335,15.000713,15.211552,15.426293,15.637131,15.851873,16.062712,15.000713,13.938716,12.8767185,11.810817,10.748819,10.71368,10.674636,10.6355915,10.600452,10.561408,10.260769,9.964035,9.663396,9.362757,9.062118,10.260769,11.4633255,12.661977,13.860628,15.063184,14.661031,14.262781,13.860628,13.462379,13.06413,13.411622,13.763018,14.114414,14.461906,14.813302,14.864059,14.9109125,14.96167,15.012426,15.063184,14.813302,14.56342,14.313539,14.063657,13.813775,14.239355,14.661031,15.086611,15.51219,15.93777,15.637131,15.336493,15.035853,14.739119,14.438479,15.875299,17.31212,18.74894,20.18576,21.626484,20.599627,19.576674,18.549814,17.526861,16.500004,15.535617,14.575133,13.610746,12.650263,11.685876,11.373524,11.061172,10.748819,10.436467,10.124115,8.663869,7.1997175,5.735567,4.2753205,2.8111696,2.6628022,2.514435,2.3621633,2.2137961,2.0615244,1.7257458,1.3860629,1.0502841,0.7106012,0.37482262,0.3357786,0.30063897,0.26159495,0.22645533,0.18741131,0.96438736,1.737459,2.514435,3.2875066,4.0605783,5.911265,7.7619514,9.612638,11.4633255,13.314012,19.350218,25.386423,31.426535,37.462738,43.498947,41.31248,39.126015,36.935646,34.74918,32.562714,31.036093,29.513376,27.986755,26.464039,24.937418,22.47374,20.013966,17.550287,15.086611,12.626837,10.6238785,8.624825,6.6257706,4.6267166,2.6237583,2.87364,3.1235218,3.3734035,3.6232853,3.873167,3.9746814,4.0761957,4.173806,4.2753205,4.376835,4.037152,3.7013733,3.3616903,3.0259118,2.6862288,2.6745155,2.6628022,2.6510892,2.639376,2.6237583,2.6237583,2.6237583,2.6237583,2.6237583,2.6237583,2.2137961,1.7999294,1.3860629,0.97610056,0.5622339,2.2255092,3.8887846,5.548156,7.211431,8.874706,7.113821,5.349031,3.5881457,1.8233559,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.6754616,0.8511597,1.0268579,1.1986516,1.3743496,1.175225,0.97610056,0.77307165,0.57394713,0.37482262,0.3357786,0.30063897,0.26159495,0.22645533,0.18741131,0.8745861,1.5617609,2.2489357,2.9361105,3.6232853,3.4983444,3.3734035,3.2484627,3.1235218,2.998581,3.0141985,3.0259118,3.0376248,3.049338,3.0610514,3.5256753,3.9863946,4.4510183,4.911738,5.376362,6.001066,6.6257706,7.250475,7.8751793,8.499884,8.086017,7.676055,7.262188,6.8483214,6.4383593,6.2860875,6.13772,5.989353,5.8370814,5.688714,5.3997884,5.1108627,4.825841,4.5369153,4.251894,3.9629683,3.6740425,3.3890212,3.1000953,2.8111696,2.5495746,2.2879796,2.0263848,1.7608855,1.4992905,1.4133936,1.3235924,1.2376955,1.1517987,1.0619974,0.8511597,0.63641757,0.42557985,0.21083772,0.0,0.999527,1.999054,2.998581,3.998108,5.001539,11.287627,17.573715,23.863707,30.149794,36.435883,30.11075,23.789522,17.460487,11.139259,4.814128,6.0635366,7.3129454,8.562354,9.811763,11.061172,16.289165,21.513256,26.737347,31.961437,37.18943,30.37625,23.563068,16.749886,9.936704,3.1235218,4.6735697,6.223617,7.773665,9.323712,10.87376,11.389141,11.900618,12.412095,12.923572,13.438952,11.900618,10.362284,8.823949,7.2856145,5.7511845,8.335898,10.924518,13.513136,16.101755,18.68647,15.113941,11.537509,7.9610763,4.388548,0.81211567,0.8511597,0.8862993,0.92534333,0.96438736,0.999527,1.4875772,1.9756275,2.463678,2.951728,3.435874,15.35211,27.260536,39.176773,51.089104,63.001434,54.025215,45.048992,36.076675,27.100456,18.124235,18.32336,18.526388,18.725513,18.924637,19.123762,22.274614,25.425468,28.57632,31.723269,34.874123,29.689075,24.500124,19.311174,14.126127,8.937177,8.101635,7.262188,6.426646,5.5871997,4.7516575,4.2753205,3.7989833,3.3265507,2.8502135,2.3738766,2.6237583,2.87364,3.1235218,3.3734035,3.6232853,3.9356375,4.251894,4.564246,4.8765984,5.1889505,4.1503797,3.1118085,2.0732377,1.038571,0.0,6.8639393,13.723974,20.587914,27.451853,34.311886,27.447948,20.587914,13.723974,6.8639393,0.0,11.162686,22.325373,33.48806,44.650745,55.81343,44.650745,33.48806,22.325373,11.162686,0.0,0.0,0.0,0.0,0.0,0.0,0.77697605,1.5500476,2.3231194,3.1000953,3.873167,3.1000953,2.3231194,1.5500476,0.77307165,0.0,1.9873407,3.9746814,5.9620223,7.9493628,9.936704,7.9493628,5.9620223,3.9746814,1.9873407,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.5622339,0.62470436,0.6871748,0.74964523,0.81211567,0.6754616,0.5388075,0.39824903,0.26159495,0.12494087,1.9873407,3.8497405,5.7121406,7.57454,9.43694,7.7619514,6.086963,4.4119744,2.736986,1.0619974,2.2879796,3.513962,4.73604,5.9620223,7.1880045,5.950309,4.7126136,3.474918,2.2372224,0.999527,0.92534333,0.8511597,0.77307165,0.698888,0.62470436,0.96438736,1.3001659,1.6359446,1.9756275,2.3114061,2.260649,2.2137961,2.1630387,2.1122816,2.0615244,1.7257458,1.3860629,1.0502841,0.7106012,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.22645533,0.38653582,0.5505207,0.7106012,0.8745861,1.1986516,1.5266213,1.8506867,2.174752,2.4988174,2.0380979,1.5734742,1.1127546,0.6481308,0.18741131,0.24988174,0.31235218,0.37482262,0.43729305,0.4997635,0.47633708,0.44900626,0.42557985,0.39824903,0.37482262,0.3357786,0.30063897,0.26159495,0.22645533,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.5622339,0.93705654,1.3118792,1.6867018,2.0615244,2.2996929,2.5378613,2.77603,3.0141985,3.2484627,2.9243972,2.6003318,2.2762666,1.9482968,1.6242313,1.7140326,1.7999294,1.8858263,1.9756275,2.0615244,2.7135596,3.3616903,4.0137253,4.661856,5.3138914,2.3231194,2.338737,2.3543546,2.3699722,2.3855898,2.4012074,2.3933985,2.3894942,2.3855898,2.3816853,2.3738766,2.2840753,2.1903696,2.096664,2.0068626,1.9131571,1.8233559,1.7335546,1.6437533,1.5539521,1.4641509,1.4914817,1.5188124,1.5461433,1.5734742,1.6008049,1.7882162,1.9756275,2.1630387,2.35045,2.5378613,2.639376,2.7408905,2.8463092,2.9478238,3.049338,3.0610514,3.076669,3.0883822,3.1000953,3.1118085,3.3148375,3.5178664,3.7208953,3.9239242,4.123049,3.8614538,3.5959544,3.330455,3.0649557,2.7994564,2.8853533,2.97125,3.0532427,3.1391394,3.2250361,2.8892577,2.5495746,2.2137961,1.8741131,1.5383345,1.796025,2.0537157,2.3114061,2.5690966,2.8267872,3.349977,3.873167,4.4002614,4.9234514,5.4505453,5.9268827,6.3993154,6.8756523,7.348085,7.824422,8.624825,9.425227,10.22563,11.0260315,11.826434,11.814721,11.806912,11.795199,11.783486,11.775677,13.673217,15.57466,17.476105,19.373644,21.275087,22.024733,22.774378,23.524023,24.273668,25.023314,22.508879,19.99054,17.4722,14.95386,12.439425,12.712734,12.986042,13.263254,13.536563,13.813775,12.501896,11.186112,9.874233,8.562354,7.250475,7.180196,7.1099167,7.039637,6.969358,6.899079,8.347612,9.796145,11.240774,12.689307,14.13784,14.336966,14.53609,14.739119,14.938243,15.137367,14.438479,13.735687,13.036799,12.337912,11.639023,11.435994,11.23687,11.037745,10.838621,10.6355915,10.186585,9.733675,9.280765,8.827853,8.374943,9.565785,10.756628,11.943566,13.134409,14.325252,13.868437,13.411622,12.950902,12.494087,12.037272,12.404286,12.767395,13.134409,13.497519,13.860628,13.899672,13.938716,13.973856,14.012899,14.051944,13.923099,13.798158,13.673217,13.548276,13.423335,13.614651,13.805966,13.993378,14.184693,14.376009,14.188598,14.005091,13.821584,13.634172,13.450665,14.383818,15.320874,16.254026,17.191084,18.124235,17.40192,16.679607,15.957292,15.234978,14.512663,13.692739,12.872814,12.05289,11.232965,10.413041,10.295909,10.178777,10.061645,9.940608,9.823476,8.550641,7.28171,6.008875,4.73604,3.4632049,3.2445583,3.0259118,2.8111696,2.592523,2.3738766,1.9834363,1.5969005,1.2064602,0.8160201,0.42557985,0.45681506,0.48805028,0.5231899,0.5544251,0.58566034,1.4407244,2.2957885,3.1508527,4.0059166,4.860981,6.2353306,7.605776,8.980125,10.350571,11.72492,17.683039,23.641155,29.599274,35.553486,41.511604,38.840992,36.174286,33.503677,30.833065,28.162453,26.862288,25.562122,24.261955,22.96179,21.661623,19.73285,17.804073,15.871395,13.94262,12.013845,10.303718,8.59359,6.883461,5.173333,3.4632049,3.4983444,3.533484,3.5686235,3.6037633,3.638903,3.736513,3.8380275,3.9356375,4.037152,4.138666,3.9356375,3.736513,3.5373883,3.338264,3.1391394,3.2367494,3.3343596,3.4280653,3.5256753,3.6232853,3.4710135,3.3187418,3.1664703,3.0141985,2.8619268,2.592523,2.3231194,2.0537157,1.7843118,1.5110037,2.7447948,3.978586,5.2084727,6.4422636,7.676055,6.1494336,4.6267166,3.1000953,1.5734742,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.30844778,0.61689556,0.92143893,1.2298868,1.5383345,1.8038338,2.0732377,2.338737,2.6081407,2.87364,2.6510892,2.4285383,2.2059872,1.9834363,1.7608855,1.5500476,1.33921,1.1244678,0.9136301,0.698888,1.1400855,1.5812829,2.018576,2.4597735,2.900971,2.8111696,2.7213683,2.631567,2.541766,2.4480603,2.5261483,2.6042364,2.6823244,2.7604125,2.8385005,3.154757,3.4710135,3.7911747,4.1074314,4.423688,5.0757227,5.7238536,6.375889,7.0240197,7.676055,7.3129454,6.949836,6.5867267,6.223617,5.8644123,5.911265,5.9620223,6.012779,6.0635366,6.114294,5.989353,5.8644123,5.735567,5.610626,5.4856853,5.056201,4.6228123,4.1894236,3.7560349,3.3265507,3.1430438,2.959537,2.77603,2.5964274,2.4129205,2.1669433,1.9209659,1.678893,1.4329157,1.1869383,1.0502841,0.9136301,0.77307165,0.63641757,0.4997635,1.4992905,2.4988174,3.4983444,4.5017757,5.5013027,10.401327,15.3013525,20.201378,25.101402,30.001427,24.785145,19.568865,14.356487,9.140205,3.9239242,4.927356,5.930787,6.9342184,7.9337454,8.937177,13.228115,17.519053,21.806087,26.097025,30.387962,25.554314,20.724567,15.890917,11.057267,6.223617,7.5667315,8.909846,10.25296,11.596075,12.939189,13.563893,14.192502,14.821111,15.445815,16.074425,14.625891,13.181262,11.732729,10.284196,8.835662,10.944039,13.052417,15.160794,17.26917,19.373644,16.535143,13.696643,10.8542385,8.015738,5.173333,4.3026514,3.4319696,2.5573835,1.6867018,0.81211567,1.7335546,2.6510892,3.5725281,4.493967,5.4115014,16.632753,27.854006,39.071354,50.292606,61.51386,54.454697,47.399445,40.340282,33.281124,26.22587,24.906181,23.590399,22.27071,20.954927,19.639143,22.122343,24.605543,27.092648,29.575848,32.06295,27.373764,22.684578,17.991486,13.302299,8.6131115,7.6526284,6.6921453,5.7316628,4.7711797,3.8106966,3.4280653,3.049338,2.6667068,2.2840753,1.901444,2.4597735,3.018103,3.5803368,4.138666,4.7009,4.970304,5.239708,5.5091114,5.7785153,6.0518236,4.841459,3.631094,2.4207294,1.2103647,0.0,5.4895897,10.979179,16.46877,21.958359,27.451853,21.958359,16.46877,10.979179,5.4895897,0.0,8.929368,17.858736,26.792007,35.721375,44.650745,35.83851,27.026272,18.214037,9.4018,0.58566034,0.5583295,0.5309987,0.5036679,0.47633708,0.44900626,1.0424755,1.6359446,2.2294137,2.8189783,3.4124475,2.7330816,2.05762,1.3782539,0.7027924,0.023426414,1.6086137,3.193801,4.7789884,6.364176,7.9493628,6.4110284,4.8687897,3.330455,1.7882162,0.24988174,0.28111696,0.30844778,0.339683,0.3709182,0.39824903,0.46852827,0.5388075,0.60908675,0.679366,0.74964523,0.62079996,0.49195468,0.359205,0.23035973,0.10151446,1.8428779,3.5842414,5.3256044,7.0708723,8.812236,7.6682463,6.5281606,5.3841705,4.2440853,3.1000953,3.631094,4.165997,4.6969957,5.2318993,5.7628975,5.251421,4.743849,4.2323723,3.7208953,3.213323,3.1391394,3.06886,2.9946766,2.9243972,2.8502135,3.0415294,3.2367494,3.4280653,3.619381,3.8106966,3.6076677,3.4007344,3.1977055,2.9907722,2.787743,2.2918842,1.7921207,1.2962615,0.79649806,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.25378615,0.44119745,0.63251317,0.8238289,1.0112402,1.3665408,1.7218413,2.077142,2.4324427,2.787743,2.2684577,1.7530766,1.2337911,0.71841,0.19912452,0.25378615,0.30454338,0.359205,0.40996224,0.46071947,0.42948425,0.39824903,0.3631094,0.3318742,0.30063897,0.27330816,0.24597734,0.21864653,0.19131571,0.1639849,0.1639849,0.1678893,0.1717937,0.1717937,0.1756981,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.22645533,0.21864653,0.20693332,0.19912452,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.4958591,0.80821127,1.116659,1.4290112,1.737459,1.9482968,2.1630387,2.3738766,2.5886188,2.7994564,2.5183394,2.241127,1.9600099,1.678893,1.4016805,1.5617609,1.7257458,1.8858263,2.0498111,2.2137961,2.7916477,3.3694992,3.9434462,4.521298,5.099149,1.901444,1.9678187,2.0341935,2.1005683,2.1708477,2.2372224,2.2294137,2.2177005,2.2059872,2.1981785,2.1864653,2.1278992,2.069333,2.0068626,1.9482968,1.8858263,1.8467822,1.8038338,1.7608855,1.717937,1.6749885,1.6906061,1.7101282,1.7257458,1.7452679,1.7608855,2.0380979,2.3114061,2.5886188,2.8619268,3.1391394,3.154757,3.174279,3.1898966,3.2094188,3.2250361,3.1235218,3.0259118,2.9243972,2.8267872,2.7252727,2.8424048,2.959537,3.076669,3.193801,3.310933,3.1079042,2.900971,2.697942,2.4910088,2.2879796,2.358259,2.4285383,2.4988174,2.5690966,2.639376,2.4480603,2.260649,2.0732377,1.8858263,1.698415,2.1513257,2.6042364,3.057147,3.5100577,3.9629683,4.2753205,4.5876727,4.900025,5.212377,5.5247293,5.813655,6.098676,6.387602,6.676528,6.9615493,7.7385254,8.511597,9.288573,10.061645,10.838621,10.780055,10.721489,10.666827,10.608261,10.549695,12.326198,14.098797,15.875299,17.651802,19.4244,20.51373,21.599154,22.688482,23.773905,24.863234,22.953981,21.040823,19.13157,17.222319,15.313066,14.813302,14.313539,13.813775,13.314012,12.814248,11.912332,11.014318,10.112402,9.21439,8.312472,7.984503,7.656533,7.328563,7.000593,6.676528,7.996216,9.315904,10.6355915,11.955279,13.274967,13.462379,13.64979,13.837202,14.024612,14.212025,13.8762455,13.536563,13.200784,12.861101,12.525322,12.162213,11.799104,11.435994,11.076789,10.71368,10.108498,9.503315,8.898132,8.292951,7.687768,8.866898,10.046027,11.229061,12.408191,13.58732,13.0719385,12.556558,12.041177,11.525795,11.014318,11.393045,11.771772,12.154405,12.533132,12.911859,12.939189,12.962616,12.986042,13.013372,13.036799,13.036799,13.036799,13.036799,13.036799,13.036799,12.993851,12.946998,12.90405,12.857197,12.814248,12.743969,12.67369,12.603411,12.533132,12.4628525,12.89624,13.325725,13.759113,14.192502,14.625891,14.204215,13.786445,13.364769,12.943093,12.525322,11.845957,11.170495,10.491129,9.815667,9.136301,9.21439,9.292478,9.370565,9.448653,9.526741,8.441318,7.3597984,6.278279,5.196759,4.1113358,3.8263142,3.541293,3.2562714,2.97125,2.6862288,2.2450314,1.8038338,1.358732,0.91753453,0.47633708,0.57785153,0.679366,0.78088045,0.8862993,0.9878138,1.9209659,2.8580225,3.7911747,4.728231,5.661383,6.559396,7.453504,8.347612,9.24172,10.135828,16.015858,21.891983,27.772013,33.64814,39.524265,36.373413,33.218655,30.067802,26.913044,23.762192,22.688482,21.610867,20.537155,19.463446,18.38583,16.991959,15.594183,14.196406,12.798631,11.400854,9.979652,8.55845,7.141152,5.7199492,4.298747,4.1191444,3.9395418,3.7599394,3.5803368,3.4007344,3.4983444,3.5998588,3.7013733,3.7989833,3.900498,3.8380275,3.775557,3.7130866,3.6506162,3.5881457,3.795079,4.0020123,4.2089458,4.415879,4.6267166,4.318269,4.0137253,3.7091823,3.4046388,3.1000953,2.97125,2.8463092,2.717464,2.5886188,2.463678,3.2640803,4.068387,4.8687897,5.6730967,6.473499,5.1889505,3.900498,2.612045,1.3235924,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5153811,1.0307622,1.5461433,2.0615244,2.5769055,2.9361105,3.2953155,3.6545205,4.0137253,4.376835,4.1308575,3.8848803,3.638903,3.39683,3.1508527,2.7643168,2.3738766,1.9873407,1.6008049,1.2142692,1.4055848,1.5969005,1.7882162,1.9834363,2.174752,2.1200905,2.0654287,2.0107672,1.9561055,1.901444,2.0420024,2.1864653,2.3270237,2.4714866,2.612045,2.7838387,2.9556324,3.1313305,3.3031244,3.474918,4.1503797,4.825841,5.5013027,6.1767645,6.8483214,6.5359693,6.223617,5.911265,5.5989127,5.2865605,5.5364423,5.786324,6.036206,6.2860875,6.5359693,6.575013,6.6140575,6.649197,6.688241,6.7233806,6.1455293,5.571582,4.9937305,4.415879,3.8380275,3.736513,3.631094,3.5295796,3.4280653,3.3265507,2.9243972,2.5183394,2.1161861,1.7140326,1.3118792,1.2494087,1.1869383,1.1244678,1.0619974,0.999527,1.999054,2.998581,3.998108,5.001539,6.001066,9.511124,13.025085,16.539047,20.049105,23.563068,19.455637,15.35211,11.248583,7.141152,3.0376248,3.7911747,4.548629,5.3021784,6.055728,6.813182,10.167064,13.520945,16.87873,20.232613,23.586494,20.73628,17.882162,15.028045,12.177831,9.323712,10.459893,11.596075,12.728352,13.864532,15.000713,15.74255,16.484386,17.226223,17.96806,18.7138,17.355068,15.996336,14.641508,13.282777,11.924045,13.55218,15.180316,16.808453,18.436588,20.06082,17.956347,15.851873,13.7474,11.642927,9.538455,7.7541428,5.9737353,4.1894236,2.4090161,0.62470436,1.979532,3.330455,4.6813784,6.036206,7.387129,17.917301,28.443571,38.969837,49.49611,60.02628,54.884182,49.74599,44.60389,39.4657,34.3236,31.489004,28.654408,25.819813,22.985216,20.15062,21.970072,23.789522,25.608974,27.428427,29.251781,25.058455,20.865126,16.671797,12.47847,8.289046,7.2036223,6.1221027,5.040583,3.959064,2.87364,2.5847144,2.2957885,2.0068626,1.7140326,1.4251068,2.2957885,3.1664703,4.0332475,4.903929,5.774611,6.001066,6.2314262,6.4578815,6.6843367,6.910792,5.5286336,4.1464753,2.7643168,1.3821584,0.0,4.1191444,8.234385,12.353529,16.46877,20.587914,16.46877,12.353529,8.234385,4.1191444,0.0,6.6960497,13.396004,20.092054,26.792007,33.48806,27.026272,20.564487,14.098797,7.6370106,1.175225,1.1205635,1.0659018,1.0112402,0.95657855,0.9019169,1.3118792,1.7218413,2.1318035,2.541766,2.951728,2.3699722,1.7882162,1.2103647,0.62860876,0.05075723,1.2337911,2.416825,3.5959544,4.7789884,5.9620223,4.8687897,3.7794614,2.6862288,1.5929961,0.4997635,0.46071947,0.42167544,0.37872702,0.339683,0.30063897,0.37872702,0.45681506,0.5309987,0.60908675,0.6871748,0.5661383,0.44119745,0.32016098,0.19912452,0.07418364,1.698415,3.3187418,4.942973,6.5633,8.187531,7.578445,6.969358,6.356367,5.74728,5.138193,4.9781127,4.8180323,4.657952,4.4978714,4.337791,4.5564375,4.7711797,4.989826,5.2084727,5.423215,5.35684,5.2865605,5.2162814,5.1460023,5.0757227,5.1225758,5.169429,5.2162814,5.263134,5.3138914,4.950782,4.591577,4.2323723,3.873167,3.513962,2.854118,2.1981785,1.5383345,0.8823949,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.28111696,0.4958591,0.7145056,0.93315214,1.1517987,1.53443,1.9209659,2.3035975,2.690133,3.076669,2.5027218,1.9287747,1.358732,0.78478485,0.21083772,0.25378615,0.29673457,0.339683,0.38263142,0.42557985,0.38653582,0.3435874,0.30454338,0.26549935,0.22645533,0.20693332,0.19131571,0.1717937,0.15617609,0.13665408,0.15617609,0.1717937,0.19131571,0.20693332,0.22645533,0.26159495,0.30063897,0.3357786,0.37482262,0.41386664,0.3670138,0.3240654,0.27721256,0.23426414,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.43338865,0.679366,0.92143893,1.1674163,1.4133936,1.6008049,1.7882162,1.9756275,2.1630387,2.35045,2.1161861,1.8819219,1.6437533,1.4094892,1.175225,1.4133936,1.6515622,1.8858263,2.1239948,2.3621633,2.8658314,3.3734035,3.8770714,4.380739,4.8883114,1.475864,1.5969005,1.7140326,1.8350691,1.9561055,2.0732377,2.0615244,2.0459068,2.0302892,2.0146716,1.999054,1.9717231,1.9443923,1.9170616,1.8897307,1.8623998,1.8663043,1.8741131,1.8780174,1.8819219,1.8858263,1.893635,1.901444,1.9092526,1.9170616,1.9248703,2.2879796,2.6510892,3.0141985,3.3734035,3.736513,3.6701381,3.6037633,3.533484,3.4671092,3.4007344,3.1859922,2.9751544,2.7643168,2.5495746,2.338737,2.3699722,2.4012074,2.436347,2.4675822,2.4988174,2.3543546,2.2098918,2.0654287,1.9209659,1.7765031,1.8311646,1.8858263,1.9404879,1.9951496,2.0498111,2.0107672,1.9756275,1.9365835,1.901444,1.8623998,2.5105307,3.1586614,3.8067923,4.4510183,5.099149,5.2006636,5.298274,5.3997884,5.5013027,5.5989127,5.700427,5.801942,5.899552,6.001066,6.098676,6.8483214,7.601871,8.351517,9.101162,9.850807,9.745388,9.639969,9.534551,9.4291315,9.323712,10.975275,12.626837,14.274494,15.926057,17.573715,18.998821,20.423927,21.849035,23.274141,24.69925,23.399082,22.095013,20.790941,19.490776,18.186707,16.91387,15.637131,14.364296,13.087557,11.810817,11.326671,10.838621,10.350571,9.86252,9.37447,8.78881,8.203149,7.621393,7.0357327,6.4500723,7.6409154,8.835662,10.0265045,11.221252,12.412095,12.587793,12.763491,12.939189,13.110983,13.286681,13.314012,13.337439,13.360865,13.388195,13.411622,12.888432,12.361338,11.838148,11.311053,10.787864,10.03041,9.272955,8.515501,7.758047,7.000593,8.171914,9.339331,10.510651,11.678067,12.849388,12.2793455,11.705398,11.131451,10.561408,9.987461,10.381805,10.77615,11.174399,11.568744,11.963089,11.974802,11.986515,11.998228,12.013845,12.025558,12.150499,12.27544,12.400381,12.525322,12.650263,12.369146,12.091934,11.810817,11.5297,11.248583,11.295436,11.338385,11.385237,11.428185,11.475039,11.404759,11.334479,11.2642,11.193921,11.123642,11.00651,10.889378,10.772245,10.655114,10.537982,10.003078,9.468176,8.933272,8.398369,7.8634663,8.136774,8.406178,8.679486,8.952794,9.226103,8.331994,7.4417906,6.547683,5.6535745,4.7633705,4.40807,4.056674,3.7052777,3.3538816,2.998581,2.5066261,2.0107672,1.5149081,1.0190489,0.5231899,0.698888,0.8706817,1.0424755,1.2142692,1.3860629,2.4012074,3.416352,4.4314966,5.446641,6.461786,6.8795567,7.297328,7.715099,8.13287,8.550641,14.348679,20.146715,25.94085,31.738886,37.536922,33.901924,30.266926,26.631927,22.99693,19.36193,18.51077,17.663515,16.812357,15.961197,15.113941,14.247164,13.384291,12.517513,11.650736,10.787864,9.655587,8.527214,7.3988423,6.266566,5.138193,4.743849,4.3455997,3.951255,3.5569105,3.1625657,3.2640803,3.3616903,3.4632049,3.5608149,3.6623292,3.736513,3.8106966,3.8887846,3.9629683,4.037152,4.3534083,4.6735697,4.989826,5.3060827,5.6262436,5.169429,4.7087092,4.251894,3.795079,3.338264,3.3538816,3.3655949,3.3812122,3.39683,3.4124475,3.7833657,4.1581883,4.5291066,4.903929,5.2748475,4.224563,3.174279,2.1239948,1.0737107,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7223144,1.4446288,2.1669433,2.8892577,3.611572,4.0644827,4.5173936,4.970304,5.423215,5.8761253,5.606722,5.3412223,5.0718184,4.806319,4.5369153,3.9746814,3.4124475,2.8502135,2.2879796,1.7257458,1.6710842,1.6164225,1.5617609,1.5031948,1.4485333,1.4290112,1.4094892,1.3899672,1.3704453,1.3509232,1.5578566,1.7647898,1.9717231,2.1786566,2.3855898,2.416825,2.4441557,2.4714866,2.4988174,2.5261483,3.2250361,3.9239242,4.6267166,5.3256044,6.0244927,5.7628975,5.5013027,5.2358036,4.9742084,4.7126136,5.1616197,5.610626,6.0635366,6.5125427,6.9615493,7.1606736,7.363703,7.562827,7.7619514,7.9610763,7.238762,6.5164475,5.794133,5.0718184,4.349504,4.3260775,4.3065557,4.283129,4.2597027,4.2362766,3.677947,3.1157131,2.5573835,1.999054,1.43682,1.4485333,1.4641509,1.475864,1.4875772,1.4992905,2.4988174,3.4983444,4.5017757,5.5013027,6.5008297,8.624825,10.748819,12.8767185,15.000713,17.124708,14.130032,11.135355,8.140678,5.1460023,2.1513257,2.6588979,3.1664703,3.6740425,4.181615,4.689187,7.1060123,9.526741,11.947471,14.3682,16.788929,15.914344,15.043662,14.169076,13.298394,12.423808,13.353056,14.278399,15.207646,16.136894,17.062239,17.921206,18.77627,19.635239,20.494207,21.349272,20.084246,18.815315,17.546383,16.281357,15.012426,16.16032,17.308216,18.45611,19.604004,20.751898,19.381453,18.011007,16.640562,15.270117,13.899672,11.205634,8.515501,5.8214636,3.1313305,0.43729305,2.2216048,4.0059166,5.794133,7.578445,9.362757,19.197947,29.033134,38.868324,48.703514,58.538704,55.313667,52.092533,48.871403,45.646366,42.425236,38.071827,33.71842,29.368914,25.015505,20.662096,21.8178,22.973503,24.129206,25.281004,26.436708,22.743143,19.045673,15.35211,11.6585455,7.9610763,6.75852,5.55206,4.3455997,3.1430438,1.9365835,1.7413634,1.542239,1.3431144,1.1478943,0.94876975,2.1318035,3.310933,4.4900627,5.6691923,6.8483214,7.0357327,7.2192397,7.406651,7.590158,7.773665,6.2197127,4.6657605,3.1118085,1.5539521,0.0,2.7447948,5.4895897,8.234385,10.979179,13.723974,10.979179,8.234385,5.4895897,2.7447948,0.0,4.466636,8.929368,13.396004,17.858736,22.325373,18.214037,14.098797,9.987461,5.8761253,1.7608855,1.678893,1.5969005,1.5149081,1.4329157,1.3509232,1.5773785,1.8038338,2.0341935,2.260649,2.4871042,2.0068626,1.5227169,1.038571,0.5583295,0.07418364,0.8550641,1.6359446,2.416825,3.193801,3.9746814,3.330455,2.6862288,2.0380979,1.3938715,0.74964523,0.64032197,0.5309987,0.42167544,0.30844778,0.19912452,0.28502136,0.3709182,0.45681506,0.5388075,0.62470436,0.5114767,0.39434463,0.28111696,0.1639849,0.05075723,1.5539521,3.0532427,4.5564375,6.0596323,7.562827,7.4847393,7.406651,7.328563,7.2543793,7.1762915,6.321227,5.4700675,4.618908,3.7638438,2.912684,3.8575494,4.802415,5.74728,6.6921453,7.6370106,7.570636,7.504261,7.433982,7.367607,7.3012323,7.2036223,7.1060123,7.008402,6.910792,6.813182,6.297801,5.7824197,5.267039,4.7516575,4.2362766,3.4202564,2.6042364,1.7843118,0.96829176,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.30844778,0.5544251,0.79649806,1.0424755,1.2884527,1.7023194,2.1161861,2.533957,2.9478238,3.3616903,2.7330816,2.1083772,1.4797685,0.8511597,0.22645533,0.25769055,0.28892577,0.3240654,0.3553006,0.38653582,0.339683,0.29283017,0.24597734,0.19912452,0.14836729,0.14055848,0.13665408,0.12884527,0.12103647,0.113227665,0.14446288,0.1756981,0.21083772,0.24207294,0.27330816,0.3357786,0.39824903,0.46071947,0.5231899,0.58566034,0.5075723,0.42557985,0.3474918,0.26940376,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.3670138,0.5466163,0.7262188,0.9058213,1.0893283,1.2494087,1.4133936,1.5734742,1.737459,1.901444,1.7101282,1.5188124,1.3314011,1.1400855,0.94876975,1.261122,1.5734742,1.8858263,2.1981785,2.514435,2.9439192,3.377308,3.8106966,4.2440853,4.6735697,1.0502841,1.2220778,1.3938715,1.5656652,1.7413634,1.9131571,1.893635,1.8741131,1.8506867,1.8311646,1.8116426,1.8194515,1.8233559,1.8272603,1.8311646,1.8389735,1.8897307,1.9443923,1.9951496,2.0459068,2.1005683,2.096664,2.096664,2.0927596,2.0888553,2.0888553,2.5378613,2.9868677,3.435874,3.8887846,4.337791,4.185519,4.0332475,3.8809757,3.7287042,3.5764325,3.2484627,2.9243972,2.6003318,2.2762666,1.9482968,1.8975395,1.8467822,1.7921207,1.7413634,1.6867018,1.6008049,1.5188124,1.4329157,1.3470187,1.261122,1.3040704,1.3431144,1.3821584,1.4212024,1.4641509,1.5734742,1.6867018,1.7999294,1.9131571,2.0263848,2.8658314,3.7091823,4.552533,5.395884,6.239235,6.126007,6.012779,5.899552,5.786324,5.6730967,5.5871997,5.5013027,5.4115014,5.3256044,5.2358036,5.9620223,6.688241,7.4144597,8.136774,8.862993,8.710721,8.55845,8.406178,8.253906,8.101635,9.6243515,11.150972,12.67369,14.200311,15.726933,17.487818,19.248703,21.013493,22.774378,24.539167,23.844185,23.1492,22.454218,21.759233,21.06425,19.014439,16.960724,14.9109125,12.861101,10.81129,10.737106,10.662923,10.588739,10.510651,10.436467,9.593117,8.75367,7.910319,7.066968,6.223617,7.289519,8.355421,9.421323,10.48332,11.549222,11.713207,11.873287,12.037272,12.201257,12.361338,12.751778,13.138313,13.524849,13.911386,14.301826,13.610746,12.923572,12.236397,11.549222,10.862047,9.952321,9.042596,8.13287,7.223144,6.3134184,7.473026,8.632633,9.792241,10.951848,12.111456,11.482847,10.8542385,10.221725,9.593117,8.960603,9.370565,9.784432,10.194394,10.604357,11.014318,11.014318,11.014318,11.014318,11.014318,11.014318,11.2642,11.514082,11.763964,12.013845,12.263727,11.748346,11.232965,10.717585,10.202203,9.686822,9.846903,10.006983,10.167064,10.327144,10.487225,9.913278,9.343235,8.769287,8.1992445,7.6252975,7.8088045,7.996216,8.179723,8.36323,8.550641,8.156297,7.7658563,7.3715115,6.9810715,6.5867267,7.055255,7.523783,7.988407,8.456935,8.925464,8.2226715,7.519879,6.817086,6.114294,5.4115014,4.9937305,4.572055,4.154284,3.7326086,3.310933,2.7643168,2.2177005,1.6710842,1.1205635,0.57394713,0.8160201,1.0580931,1.3040704,1.5461433,1.7882162,2.8814487,3.978586,5.0718184,6.168956,7.262188,7.2036223,7.141152,7.082586,7.0240197,6.9615493,12.681499,18.397543,24.113588,29.833538,35.549583,31.434343,27.315199,23.196054,19.080814,14.96167,14.336966,13.712261,13.087557,12.4628525,11.838148,11.506273,11.174399,10.838621,10.506746,10.174872,9.335425,8.495979,7.656533,6.813182,5.9737353,5.364649,4.755562,4.1464753,3.533484,2.9243972,3.0259118,3.1235218,3.2250361,3.3265507,3.4241607,3.638903,3.8497405,4.0605783,4.2753205,4.4861584,4.9156423,5.3412223,5.7707067,6.196286,6.6257706,6.016684,5.4036927,4.794606,4.185519,3.5764325,3.7326086,3.8887846,4.0488653,4.2050414,4.3612175,4.3065557,4.2479897,4.1894236,4.1308575,4.0761957,3.2640803,2.4519646,1.6359446,0.8238289,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.92924774,1.8584955,2.7916477,3.7208953,4.650143,5.196759,5.7394714,6.2860875,6.8287997,7.375416,7.08649,6.79366,6.504734,6.2158084,5.9268827,5.1889505,4.4510183,3.7130866,2.9751544,2.2372224,1.9365835,1.6320401,1.3314011,1.0268579,0.7262188,0.7418364,0.75354964,0.76916724,0.78478485,0.80040246,1.0737107,1.3431144,1.6164225,1.8897307,2.1630387,2.0459068,1.9287747,1.8116426,1.6906061,1.5734742,2.2996929,3.0259118,3.7482262,4.474445,5.2006636,4.985922,4.775084,4.564246,4.349504,4.138666,4.786797,5.4388323,6.086963,6.7389984,7.387129,7.7502384,8.113348,8.476458,8.835662,9.198771,8.331994,7.465217,6.5984397,5.7316628,4.860981,4.919547,4.9781127,5.036679,5.0913405,5.1499066,4.4314966,3.7130866,2.998581,2.280171,1.5617609,1.6515622,1.737459,1.8233559,1.9131571,1.999054,2.998581,3.998108,5.001539,6.001066,7.000593,7.7385254,8.476458,9.21439,9.948417,10.686349,8.800523,6.918601,5.0327744,3.1469483,1.261122,1.5227169,1.7843118,2.0420024,2.3035975,2.5612879,4.0488653,5.532538,7.016211,8.503788,9.987461,11.096312,12.201257,13.310107,14.418958,15.523903,16.246218,16.964628,17.686943,18.405352,19.123762,20.095959,21.068155,22.044254,23.01645,23.988647,22.809519,21.634293,20.455164,19.276033,18.10081,18.768461,19.436115,20.103767,20.77142,21.439074,20.802654,20.166237,19.533724,18.897306,18.26089,14.661031,11.057267,7.453504,3.853645,0.24988174,2.4675822,4.6852827,6.902983,9.120684,11.338385,20.482494,29.6227,38.76681,47.907017,57.051125,55.743153,54.43908,53.13501,51.83094,50.52687,44.654648,38.78633,32.914112,27.045794,21.173573,21.665527,22.153578,22.645533,23.133583,23.625538,20.427834,17.230127,14.032422,10.834716,7.6370106,6.309514,4.9820175,3.6545205,2.3270237,0.999527,0.8941081,0.78868926,0.6832704,0.58175594,0.47633708,1.9639144,3.455396,4.9468775,6.434455,7.9259367,8.066495,8.210958,8.351517,8.495979,8.636538,6.910792,5.181142,3.455396,1.7257458,0.0,1.3743496,2.7447948,4.1191444,5.4895897,6.8639393,5.4895897,4.1191444,2.7447948,1.3743496,0.0,2.233318,4.466636,6.6960497,8.929368,11.162686,9.4018,7.6370106,5.8761253,4.1113358,2.35045,2.241127,2.1318035,2.018576,1.9092526,1.7999294,1.8467822,1.8897307,1.9365835,1.979532,2.0263848,1.639849,1.2533131,0.8706817,0.48414588,0.10151446,0.47633708,0.8550641,1.2337911,1.6086137,1.9873407,1.7882162,1.5929961,1.3938715,1.1986516,0.999527,0.8199245,0.64032197,0.46071947,0.28111696,0.10151446,0.19131571,0.28502136,0.37872702,0.46852827,0.5622339,0.45681506,0.3474918,0.23816854,0.13274968,0.023426414,1.4094892,2.7916477,4.173806,5.5559645,6.9381227,7.3910336,7.8478484,8.300759,8.757574,9.21439,7.6682463,6.1221027,4.575959,3.0337205,1.4875772,3.1586614,4.83365,6.504734,8.175818,9.850807,9.784432,9.718058,9.655587,9.589212,9.526741,9.280765,9.0386915,8.796618,8.554545,8.312472,7.6409154,6.9732623,6.3017054,5.6340523,4.9624953,3.9863946,3.0063896,2.0302892,1.0541886,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.3357786,0.60908675,0.8784905,1.1517987,1.4251068,1.8702087,2.3153105,2.7604125,3.2055142,3.6506162,2.9673457,2.2840753,1.6008049,0.92143893,0.23816854,0.26159495,0.28111696,0.30454338,0.3279698,0.3513962,0.29673457,0.23816854,0.1835069,0.12884527,0.07418364,0.078088045,0.078088045,0.08199245,0.08589685,0.08589685,0.13665408,0.1835069,0.23035973,0.27721256,0.3240654,0.41386664,0.4997635,0.58566034,0.6754616,0.76135844,0.6481308,0.5309987,0.41777104,0.30063897,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.30063897,0.41777104,0.5309987,0.6481308,0.76135844,0.9019169,1.038571,1.175225,1.3118792,1.4485333,1.3040704,1.1596074,1.0151446,0.8706817,0.7262188,1.1127546,1.4992905,1.8858263,2.2762666,2.6628022,3.0220075,3.3812122,3.7443218,4.1035266,4.462732,0.62470436,0.8511597,1.0737107,1.3001659,1.5266213,1.7491722,1.7257458,1.698415,1.6749885,1.6515622,1.6242313,1.6632754,1.698415,1.737459,1.7765031,1.8116426,1.9131571,2.0107672,2.1122816,2.2137961,2.3114061,2.2996929,2.2879796,2.2762666,2.260649,2.2489357,2.787743,3.3265507,3.8614538,4.4002614,4.939069,4.7009,4.462732,4.224563,3.9863946,3.7482262,3.310933,2.87364,2.436347,1.999054,1.5617609,1.4251068,1.2884527,1.1517987,1.0112402,0.8745861,0.8511597,0.8238289,0.80040246,0.77307165,0.74964523,0.77307165,0.80040246,0.8238289,0.8511597,0.8745861,1.1361811,1.4016805,1.6632754,1.9248703,2.1864653,3.2250361,4.263607,5.298274,6.336845,7.375416,7.0513506,6.7233806,6.3993154,6.0752497,5.7511845,5.473972,5.2006636,4.9234514,4.650143,4.376835,5.0757227,5.774611,6.473499,7.1762915,7.8751793,7.676055,7.47693,7.2739015,7.0747766,6.8756523,8.273428,9.675109,11.076789,12.4745655,13.8762455,15.976814,18.073479,20.174046,22.274614,24.375183,24.289286,24.199486,24.113588,24.023787,23.937891,21.111103,18.28822,15.461433,12.63855,9.811763,10.151445,10.487225,10.826907,11.162686,11.498465,10.401327,9.300286,8.1992445,7.098203,6.001066,6.9381227,7.8751793,8.812236,9.749292,10.686349,10.838621,10.986988,11.139259,11.287627,11.435994,12.185639,12.939189,13.688834,14.438479,15.188125,14.336966,13.4858055,12.63855,11.787391,10.936231,9.874233,8.812236,7.7502384,6.688241,5.6262436,6.774138,7.9259367,9.073831,10.22563,11.373524,10.686349,9.999174,9.311999,8.624825,7.9376497,8.36323,8.78881,9.21439,9.636065,10.061645,10.049932,10.0382185,10.0265045,10.010887,9.999174,10.373997,10.748819,11.123642,11.498465,11.873287,11.123642,10.373997,9.6243515,8.874706,8.125061,8.398369,8.675582,8.94889,9.226103,9.499411,8.4257,7.348085,6.2743745,5.2006636,4.123049,4.6110992,5.099149,5.5871997,6.0752497,6.5633,6.3134184,6.0635366,5.813655,5.563773,5.3138914,5.9737353,6.6374836,7.3012323,7.9610763,8.624825,8.113348,7.601871,7.08649,6.575013,6.0635366,5.575486,5.087436,4.5993857,4.1113358,3.6232853,3.0259118,2.4246337,1.8233559,1.2259823,0.62470436,0.93705654,1.2494087,1.5617609,1.8741131,2.1864653,3.3616903,4.5369153,5.7121406,6.8873653,8.062591,7.523783,6.98888,6.4500723,5.911265,5.376362,11.014318,16.64837,22.286327,27.924286,33.56224,28.962856,24.36347,19.764084,15.160794,10.561408,10.163159,9.761005,9.362757,8.960603,8.562354,8.761478,8.960603,9.163632,9.362757,9.561881,9.01136,8.460839,7.914223,7.363703,6.813182,5.989353,5.1616197,4.337791,3.513962,2.6862288,2.787743,2.8892577,2.9868677,3.0883822,3.1859922,3.5373883,3.8887846,4.2362766,4.5876727,4.939069,5.473972,6.012779,6.551587,7.08649,7.6252975,6.8639393,6.098676,5.337318,4.575959,3.8106966,4.1113358,4.4119744,4.7126136,5.0132523,5.3138914,4.825841,4.337791,3.8497405,3.3616903,2.87364,2.2996929,1.7257458,1.1517987,0.57394713,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1361811,2.2762666,3.4124475,4.548629,5.688714,6.3251314,6.9615493,7.601871,8.238289,8.874706,8.562354,8.250002,7.9376497,7.6252975,7.3129454,6.3993154,5.4856853,4.575959,3.6623292,2.7486992,2.1981785,1.6515622,1.1010414,0.5505207,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.58566034,0.92534333,1.261122,1.6008049,1.9365835,1.6749885,1.4133936,1.1517987,0.8862993,0.62470436,1.3743496,2.1239948,2.87364,3.6232853,4.376835,4.21285,4.0488653,3.8887846,3.7247996,3.5608149,4.4119744,5.263134,6.114294,6.9615493,7.812709,8.335898,8.862993,9.386183,9.913278,10.436467,9.425227,8.413987,7.3988423,6.387602,5.376362,5.5130157,5.64967,5.786324,5.9268827,6.0635366,5.1889505,4.3143644,3.435874,2.5612879,1.6867018,1.8506867,2.0107672,2.174752,2.338737,2.4988174,3.4983444,4.5017757,5.5013027,6.5008297,7.5003567,6.8483214,6.2001905,5.548156,4.900025,4.251894,3.474918,2.7018464,1.9248703,1.1517987,0.37482262,0.38653582,0.39824903,0.41386664,0.42557985,0.43729305,0.9878138,1.5383345,2.0888553,2.639376,3.1859922,6.2743745,9.362757,12.4511385,15.535617,18.623999,19.13938,19.650856,20.162333,20.67381,21.189192,22.274614,23.363943,24.449368,25.538694,26.624119,25.538694,24.449368,23.363943,22.274614,21.189192,21.376602,21.564014,21.751425,21.938837,22.126247,22.223858,22.325373,22.426888,22.524496,22.62601,18.112522,13.599033,9.085544,4.575959,0.062470436,2.7135596,5.3607445,8.011833,10.662923,13.314012,21.763138,30.212265,38.661392,47.11442,55.56355,56.17654,56.785625,57.398617,58.01161,58.6246,51.237473,43.85034,36.46321,29.076084,21.688955,21.513256,21.337559,21.16186,20.986162,20.81437,18.112522,15.410676,12.712734,10.010887,7.3129454,5.860508,4.4119744,2.9634414,1.5110037,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,1.7999294,3.5998588,5.3997884,7.1997175,8.999647,9.101162,9.198771,9.300286,9.4018,9.499411,7.5979667,5.700427,3.7989833,1.901444,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.58566034,1.175225,1.7608855,2.35045,2.9361105,2.7994564,2.6628022,2.5261483,2.3855898,2.2489357,2.1122816,1.9756275,1.8389735,1.698415,1.5617609,1.2767396,0.9878138,0.698888,0.41386664,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.24988174,0.4997635,0.74964523,0.999527,1.2494087,0.999527,0.74964523,0.4997635,0.24988174,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,1.261122,2.5261483,3.78727,5.0483923,6.3134184,7.3012323,8.289046,9.276859,10.260769,11.248583,9.01136,6.774138,4.5369153,2.2996929,0.062470436,2.463678,4.860981,7.262188,9.663396,12.0606985,11.998228,11.935758,11.873287,11.810817,11.748346,11.361811,10.975275,10.588739,10.198298,9.811763,8.987934,8.164105,7.336372,6.5125427,5.688714,4.548629,3.4124475,2.2762666,1.1361811,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.3631094,0.6637484,0.96438736,1.261122,1.5617609,2.0380979,2.514435,2.9868677,3.4632049,3.9356375,3.2016098,2.463678,1.7257458,0.9878138,0.24988174,0.26159495,0.27330816,0.28892577,0.30063897,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.37482262,0.48805028,0.60127795,0.7106012,0.8238289,0.93705654,0.78868926,0.63641757,0.48805028,0.3357786,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.23816854,0.28892577,0.3357786,0.38653582,0.43729305,0.5505207,0.6637484,0.77307165,0.8862993,0.999527,0.9019169,0.80040246,0.698888,0.60127795,0.4997635,0.96438736,1.4251068,1.8858263,2.35045,2.8111696,3.1000953,3.3890212,3.6740425,3.9629683,4.251894,0.92534333,1.0932326,1.261122,1.4290112,1.5969005,1.7608855,1.7335546,1.7023194,1.6710842,1.6437533,1.6125181,1.6125181,1.6125181,1.6125181,1.6125181,1.6125181,1.7140326,1.8116426,1.9131571,2.0107672,2.1122816,2.1005683,2.0888553,2.0732377,2.0615244,2.0498111,2.463678,2.8814487,3.2953155,3.7091823,4.123049,3.9083066,3.68966,3.4710135,3.2562714,3.0376248,2.6823244,2.3270237,1.9717231,1.6164225,1.261122,1.1557031,1.0541886,0.94876975,0.8433509,0.737932,0.78478485,0.8316377,0.8784905,0.92924774,0.97610056,0.9917182,1.0112402,1.0268579,1.0463798,1.0619974,1.358732,1.6515622,1.9482968,2.241127,2.5378613,3.4632049,4.388548,5.3138914,6.239235,7.1606736,6.8756523,6.5867267,6.3017054,6.012779,5.7238536,5.5091114,5.290465,5.0718184,4.853172,4.6384296,5.1889505,5.735567,6.2860875,6.8366084,7.387129,7.3246584,7.262188,7.1997175,7.137247,7.0747766,8.156297,9.24172,10.323239,11.404759,12.486279,14.067561,15.648844,17.226223,18.807507,20.388788,20.423927,20.459068,20.494207,20.529346,20.560583,18.22575,15.890917,13.556085,11.221252,8.886419,9.120684,9.351044,9.585307,9.815667,10.049932,9.24172,8.429605,7.621393,6.8092775,6.001066,7.2153354,8.429605,9.643873,10.858143,12.076316,11.783486,11.490656,11.197825,10.904996,10.612165,11.283723,11.951375,12.622932,13.2905855,13.962143,13.087557,12.212971,11.338385,10.4637985,9.589212,8.675582,7.7619514,6.8483214,5.938596,5.024966,6.168956,7.3168497,8.460839,9.60483,10.748819,10.034314,9.319808,8.605303,7.890797,7.1762915,7.5276875,7.8790836,8.234385,8.58578,8.937177,9.085544,9.2339115,9.378374,9.526741,9.675109,10.018696,10.366188,10.709775,11.053363,11.400854,10.71368,10.03041,9.343235,8.659965,7.9766936,8.113348,8.253906,8.3944645,8.535024,8.675582,7.6916723,6.7116675,5.727758,4.743849,3.7638438,4.181615,4.60329,5.0210614,5.4427366,5.8644123,5.8566036,5.8487945,5.840986,5.833177,5.825368,6.196286,6.571109,6.942027,7.3168497,7.687768,7.211431,6.7311897,6.2548523,5.7785153,5.298274,4.884407,4.466636,4.0488653,3.631094,3.213323,2.7643168,2.3192148,1.8702087,1.4212024,0.97610056,1.2767396,1.5734742,1.8741131,2.174752,2.475391,3.4983444,4.521298,5.5442514,6.5633,7.5862536,7.1216297,6.6531014,6.184573,5.716045,5.251421,9.866425,14.4853325,19.10424,23.719244,28.338152,24.613352,20.888552,17.163752,13.438952,9.714153,9.390087,9.066022,8.745861,8.421796,8.101635,8.331994,8.566258,8.796618,9.030883,9.261242,9.101162,8.937177,8.773191,8.6131115,8.449126,7.605776,6.75852,5.9151692,5.0718184,4.224563,4.056674,3.8887846,3.7208953,3.5569105,3.3890212,3.7911747,4.1972322,4.60329,5.009348,5.4115014,5.911265,6.4110284,6.910792,7.4144597,7.914223,7.4144597,6.910792,6.4110284,5.911265,5.4115014,5.251421,5.0913405,4.93126,4.7711797,4.6110992,4.1503797,3.6857557,3.2250361,2.7643168,2.2996929,1.8389735,1.3782539,0.92143893,0.46071947,0.0,0.046852827,0.08980125,0.13665408,0.1796025,0.22645533,0.19912452,0.1756981,0.14836729,0.12494087,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,1.0268579,2.0537157,3.084478,4.1113358,5.138193,5.8175592,6.4969254,7.1762915,7.8556576,8.538928,8.097731,7.656533,7.2192397,6.7780423,6.336845,5.520825,4.7009,3.8848803,3.06886,2.2489357,1.901444,1.5539521,1.2064602,0.8589685,0.5114767,0.47633708,0.43729305,0.39824903,0.3631094,0.3240654,0.58566034,0.8511597,1.1127546,1.3743496,1.6359446,1.4133936,1.1869383,0.96438736,0.737932,0.5114767,1.116659,1.717937,2.3192148,2.9243972,3.5256753,3.4632049,3.4046388,3.3460727,3.2836022,3.2250361,3.9356375,4.650143,5.3607445,6.0752497,6.785851,7.473026,8.156297,8.843472,9.526741,10.213917,9.468176,8.726339,7.984503,7.2426662,6.5008297,6.7233806,6.949836,7.1762915,7.3988423,7.6252975,6.606249,5.5832953,4.564246,3.5451972,2.5261483,2.9087796,3.2914112,3.6740425,4.056674,4.4393053,4.93126,5.423215,5.9151692,6.407124,6.899079,6.4422636,5.985449,5.5286336,5.0718184,4.6110992,4.0801005,3.5491016,3.0141985,2.4831998,1.9482968,1.8741131,1.7999294,1.7257458,1.6515622,1.5734742,1.8311646,2.0888553,2.3465457,2.6042364,2.8619268,5.270943,7.6838636,10.09288,12.501896,14.9109125,15.594183,16.273548,16.952915,17.63228,18.311647,19.373644,20.435642,21.501543,22.563541,23.625538,22.645533,21.665527,20.685524,19.705519,18.725513,19.162806,19.6001,20.037392,20.474686,20.911978,20.494207,20.076437,19.658665,19.240894,18.823124,15.070992,11.314958,7.558923,3.8067923,0.05075723,2.8345962,5.6145306,8.398369,11.178304,13.962143,20.119385,26.272722,32.42606,38.5833,44.73664,45.298874,45.86111,46.423344,46.985577,47.551716,41.6873,35.826794,29.962383,24.097971,18.237463,18.221846,18.206228,18.19061,18.178898,18.163279,15.824542,13.4858055,11.150972,8.812236,6.473499,5.559869,4.646239,3.7287042,2.815074,1.901444,1.7101282,1.5188124,1.3314011,1.1400855,0.94876975,2.4480603,3.9434462,5.4427366,6.9381227,8.437413,8.421796,8.406178,8.39056,8.378847,8.36323,6.688241,5.017157,3.3460727,1.6710842,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.47243267,0.94486535,1.4172981,1.8897307,2.3621633,2.4246337,2.4871042,2.5495746,2.612045,2.6745155,2.4207294,2.1669433,1.9092526,1.6554666,1.4016805,1.1400855,0.8784905,0.62079996,0.359205,0.10151446,0.26159495,0.42167544,0.58175594,0.7418364,0.9019169,0.92143893,0.94096094,0.96048295,0.98000497,0.999527,0.80040246,0.60127795,0.39824903,0.19912452,0.0,0.13665408,0.27330816,0.41386664,0.5505207,0.6871748,0.79649806,0.9019169,1.0112402,1.116659,1.2259823,2.3933985,3.5647192,4.73604,5.903456,7.0747766,7.461313,7.843944,8.23048,8.6131115,8.999647,7.2153354,5.4310236,3.6467118,1.8584955,0.07418364,1.9912452,3.9083066,5.8292727,7.746334,9.663396,9.721962,9.784432,9.8429985,9.901564,9.964035,9.651682,9.339331,9.023073,8.710721,8.398369,7.715099,7.0318284,6.3446536,5.661383,4.9742084,3.978586,2.9868677,1.9912452,0.9956226,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.58956474,1.0815194,1.5695697,2.0615244,2.5495746,3.1781836,3.8067923,4.4314966,5.0601053,5.688714,5.0718184,4.4588275,3.8419318,3.2289407,2.612045,2.2762666,1.9443923,1.6086137,1.2728351,0.93705654,0.8160201,0.6910792,0.5700427,0.44900626,0.3240654,0.3318742,0.339683,0.3474918,0.3553006,0.3631094,0.3631094,0.3670138,0.3709182,0.3709182,0.37482262,0.5036679,0.62860876,0.75745404,0.8862993,1.0112402,0.92924774,0.8472553,0.76526284,0.6832704,0.60127795,0.5583295,0.5192855,0.48024148,0.44119745,0.39824903,0.42948425,0.46071947,0.48805028,0.5192855,0.5505207,0.60127795,0.6559396,0.7066968,0.76135844,0.81211567,0.74964523,0.6871748,0.62470436,0.5622339,0.4997635,0.97610056,1.4485333,1.9248703,2.4012074,2.87364,3.1469483,3.4202564,3.6935644,3.9668727,4.2362766,1.2259823,1.3353056,1.4446288,1.5539521,1.6632754,1.7765031,1.7413634,1.7062237,1.6710842,1.6359446,1.6008049,1.5617609,1.5266213,1.4875772,1.4485333,1.4133936,1.5110037,1.6125181,1.7140326,1.8116426,1.9131571,1.901444,1.8858263,1.8741131,1.8623998,1.8506867,2.1435168,2.436347,2.7291772,3.018103,3.310933,3.1157131,2.9165885,2.7213683,2.522244,2.3231194,2.0537157,1.7804074,1.5070993,1.2337911,0.96438736,0.8902037,0.8160201,0.74574083,0.6715572,0.60127795,0.71841,0.8394465,0.96048295,1.0815194,1.1986516,1.2103647,1.2181735,1.2298868,1.2415999,1.2494087,1.5773785,1.9053483,2.233318,2.5612879,2.8892577,3.7013733,4.513489,5.3256044,6.13772,6.949836,6.699954,6.4500723,6.2001905,5.950309,5.700427,5.5403466,5.380266,5.2201858,5.0601053,4.900025,5.298274,5.700427,6.098676,6.5008297,6.899079,6.9732623,7.0513506,7.125534,7.1997175,7.2739015,8.039165,8.804427,9.56969,10.334952,11.100216,12.158309,13.220306,14.278399,15.340397,16.398489,16.55857,16.714746,16.870922,17.031002,17.18718,15.344301,13.497519,11.650736,9.807858,7.9610763,8.089922,8.218767,8.343708,8.472553,8.601398,8.078208,7.558923,7.039637,6.520352,6.001066,7.492548,8.98403,10.479416,11.970898,13.462379,12.728352,11.994324,11.256392,10.522364,9.788337,10.377901,10.967466,11.557031,12.146595,12.73616,11.838148,10.936231,10.0382185,9.136301,8.238289,7.47693,6.7116675,5.950309,5.1889505,4.423688,5.563773,6.703859,7.843944,8.98403,10.124115,9.382278,8.640442,7.898606,7.1567693,6.4110284,6.6921453,6.9732623,7.2543793,7.531592,7.812709,8.121157,8.4257,8.734148,9.042596,9.351044,9.663396,9.979652,10.295909,10.608261,10.924518,10.303718,9.686822,9.066022,8.445222,7.824422,7.8283267,7.8361354,7.8400397,7.843944,7.8517528,6.9615493,6.0713453,5.181142,4.290938,3.4007344,3.7521305,4.1035266,4.4588275,4.8102236,5.1616197,5.395884,5.6340523,5.8683167,6.1025805,6.336845,6.4188375,6.5008297,6.5867267,6.6687193,6.7507114,6.3056097,5.8644123,5.423215,4.9781127,4.5369153,4.1894236,3.8419318,3.49444,3.1469483,2.7994564,2.5066261,2.2098918,1.9131571,1.620327,1.3235924,1.6125181,1.901444,2.1864653,2.475391,2.7643168,3.631094,4.5017757,5.3724575,6.2431393,7.113821,6.715572,6.3173227,5.919074,5.520825,5.12648,8.722435,12.318389,15.918248,19.514202,23.114061,20.263847,17.413633,14.56342,11.713207,8.862993,8.617016,8.371038,8.128965,7.882988,7.6370106,7.90251,8.16801,8.433509,8.699008,8.960603,9.187058,9.413514,9.636065,9.86252,10.088976,9.2221985,8.359325,7.492548,6.6257706,5.7628975,5.3256044,4.892216,4.4588275,4.0215344,3.5881457,4.0488653,4.50568,4.9663997,5.4271193,5.8878384,6.348558,6.813182,7.2739015,7.7385254,8.1992445,7.9610763,7.726812,7.4886436,7.250475,7.012306,6.3915067,5.7707067,5.153811,4.533011,3.912211,3.474918,3.0376248,2.6003318,2.1630387,1.7257458,1.3782539,1.0346665,0.6910792,0.3435874,0.0,0.08980125,0.1796025,0.26940376,0.359205,0.44900626,0.39824903,0.3513962,0.30063897,0.24988174,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.91753453,1.8350691,2.7526035,3.6701381,4.5876727,5.309987,6.0323014,6.754616,7.47693,8.1992445,7.633106,7.066968,6.4969254,5.930787,5.3607445,4.6384296,3.9161155,3.193801,2.4714866,1.7491722,1.6047094,1.4602464,1.3157835,1.1713207,1.0268579,0.9019169,0.77307165,0.6481308,0.5231899,0.39824903,0.58566034,0.77307165,0.96438736,1.1517987,1.33921,1.1517987,0.96438736,0.77307165,0.58566034,0.39824903,0.8550641,1.3118792,1.7647898,2.2216048,2.6745155,2.717464,2.7604125,2.803361,2.8463092,2.8892577,3.4632049,4.037152,4.6110992,5.1889505,5.7628975,6.606249,7.453504,8.296855,9.14411,9.987461,9.515028,9.042596,8.570163,8.097731,7.6252975,7.9376497,8.250002,8.562354,8.874706,9.187058,8.023546,6.8561306,5.6926184,4.5291066,3.3616903,3.9668727,4.5681505,5.169429,5.7707067,6.375889,6.3602715,6.3446536,6.329036,6.3134184,6.3017054,6.036206,5.7707067,5.505207,5.239708,4.9742084,4.6852827,4.396357,4.1035266,3.814601,3.5256753,3.3616903,3.2016098,3.0376248,2.87364,2.7135596,2.67842,2.6432803,2.6081407,2.5730011,2.5378613,4.271416,6.001066,7.734621,9.468176,11.20173,12.0489855,12.89624,13.743496,14.590752,15.438006,16.476578,17.511244,18.549814,19.588387,20.626957,19.75237,18.88169,18.007103,17.136421,16.261835,16.94901,17.636185,18.32336,19.014439,19.701614,18.764557,17.831406,16.894348,15.961197,15.024139,12.025558,9.030883,6.0323014,3.0337205,0.039044023,2.951728,5.8683167,8.781001,11.697589,14.614178,18.471727,22.333181,26.190731,30.052185,33.91364,34.425114,34.936592,35.451973,35.963448,36.474926,32.137135,27.799343,23.461554,19.123762,14.785972,14.934339,15.078801,15.223265,15.367727,15.51219,13.536563,11.560935,9.589212,7.6135845,5.6379566,5.2592297,4.8765984,4.4978714,4.1191444,3.736513,3.3694992,3.0024853,2.6354716,2.2684577,1.901444,3.096191,4.290938,5.4856853,6.6804323,7.8751793,7.746334,7.6135845,7.4847393,7.355894,7.223144,5.7785153,4.3338866,2.8892577,1.4446288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.359205,0.7145056,1.0737107,1.4290112,1.7882162,2.0498111,2.3114061,2.5769055,2.8385005,3.1000953,2.7291772,2.3543546,1.9834363,1.6086137,1.2376955,1.0034313,0.77307165,0.5388075,0.30844778,0.07418364,0.42167544,0.76526284,1.1088502,1.456342,1.7999294,1.5890918,1.3782539,1.1713207,0.96048295,0.74964523,0.60127795,0.44900626,0.30063897,0.14836729,0.0,0.1756981,0.3513962,0.5231899,0.698888,0.8745861,1.1908426,1.5031948,1.8194515,2.135708,2.4480603,3.5256753,4.60329,5.6809053,6.75852,7.8361354,7.621393,7.4027467,7.1841,6.969358,6.7507114,5.4193106,4.084005,2.7526035,1.4212024,0.08589685,1.5227169,2.9556324,4.3924527,5.8292727,7.262188,7.445695,7.629202,7.8088045,7.9923115,8.175818,7.9376497,7.699481,7.461313,7.223144,6.98888,6.4422636,5.8956475,5.3529353,4.806319,4.263607,3.408543,2.5573835,1.7062237,0.8511597,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.13665408,0.8160201,1.4992905,2.1786566,2.8580225,3.5373883,4.318269,5.099149,5.8761253,6.657006,7.437886,6.9459314,6.453977,5.958118,5.466163,4.9742084,4.290938,3.611572,2.9283018,2.2450314,1.5617609,1.3782539,1.1986516,1.0151446,0.8316377,0.6481308,0.6520352,0.6559396,0.6559396,0.659844,0.6637484,0.60518235,0.5466163,0.48805028,0.43338865,0.37482262,0.5192855,0.659844,0.80430686,0.94486535,1.0893283,1.0737107,1.0580931,1.0424755,1.0268579,1.0112402,0.93315214,0.8511597,0.77307165,0.6910792,0.61299115,0.62079996,0.63251317,0.6442264,0.6520352,0.6637484,0.6559396,0.6481308,0.64032197,0.63251317,0.62470436,0.60127795,0.57394713,0.5505207,0.5231899,0.4997635,0.9878138,1.475864,1.9639144,2.4480603,2.9361105,3.193801,3.4514916,3.7091823,3.9668727,4.224563,1.5266213,1.5773785,1.6281357,1.6827974,1.7335546,1.7882162,1.7491722,1.7062237,1.6671798,1.6281357,1.5890918,1.5110037,1.43682,1.3626363,1.2884527,1.2142692,1.3118792,1.4133936,1.5110037,1.6125181,1.7140326,1.698415,1.6867018,1.6749885,1.6632754,1.6515622,1.8194515,1.9912452,2.1591344,2.330928,2.4988174,2.3231194,2.1435168,1.9678187,1.7882162,1.6125181,1.4212024,1.2337911,1.0424755,0.8511597,0.6637484,0.62079996,0.58175594,0.5427119,0.5036679,0.46071947,0.6559396,0.8472553,1.038571,1.2337911,1.4251068,1.4290112,1.4290112,1.4329157,1.43682,1.43682,1.796025,2.1591344,2.5183394,2.8775444,3.2367494,3.9356375,4.6384296,5.337318,6.036206,6.7389984,6.524256,6.3134184,6.098676,5.8878384,5.6730967,5.571582,5.4700675,5.368553,5.263134,5.1616197,5.4115014,5.661383,5.911265,6.1611466,6.4110284,6.6257706,6.8366084,7.0513506,7.262188,7.47693,7.9220324,8.371038,8.81614,9.265146,9.714153,10.25296,10.791768,11.330575,11.873287,12.412095,12.693212,12.974329,13.251541,13.532659,13.813775,12.458947,11.10412,9.749292,8.39056,7.0357327,7.0591593,7.082586,7.1060123,7.1294384,7.1489606,6.918601,6.688241,6.461786,6.2314262,6.001066,7.7697606,9.538455,11.311053,13.079747,14.848442,13.673217,12.494087,11.318862,10.139732,8.960603,9.47208,9.983557,10.491129,11.002605,11.514082,10.588739,9.663396,8.738052,7.812709,6.8873653,6.2743745,5.661383,5.0483923,4.4393053,3.8263142,4.958591,6.094772,7.230953,8.36323,9.499411,8.730244,7.9610763,7.191909,6.4188375,5.64967,5.8566036,6.0635366,6.2743745,6.481308,6.688241,7.1567693,7.621393,8.089922,8.55845,9.023073,9.308095,9.593117,9.878138,10.163159,10.44818,9.893755,9.339331,8.784905,8.23048,7.676055,7.5433054,7.4144597,7.2856145,7.1567693,7.0240197,6.2275214,5.4310236,4.630621,3.8341231,3.0376248,3.3226464,3.6076677,3.892689,4.1777105,4.462732,4.939069,5.4193106,5.8956475,6.3719845,6.8483214,6.6413884,6.434455,6.2275214,6.0205884,5.813655,5.4036927,4.997635,4.591577,4.181615,3.775557,3.4983444,3.2211318,2.9439192,2.6667068,2.3855898,2.2450314,2.1005683,1.9600099,1.815547,1.6749885,1.9482968,2.2255092,2.4988174,2.77603,3.049338,3.767748,4.4861584,5.2006636,5.919074,6.6374836,6.309514,5.9815445,5.6535745,5.3256044,5.001539,7.578445,10.155351,12.732256,15.309161,17.886066,15.914344,13.938716,11.963089,9.987461,8.011833,7.843944,7.676055,7.5081654,7.3441806,7.1762915,7.473026,7.7697606,8.066495,8.36323,8.663869,9.276859,9.885946,10.498938,11.111929,11.72492,10.838621,9.956225,9.069926,8.183627,7.3012323,6.5984397,5.8956475,5.192855,4.4900627,3.78727,4.3026514,4.8180323,5.3334136,5.8487945,6.364176,6.785851,7.211431,7.6370106,8.062591,8.488171,8.511597,8.538928,8.562354,8.58578,8.6131115,7.531592,6.453977,5.3724575,4.290938,3.213323,2.7994564,2.3855898,1.9756275,1.5617609,1.1517987,0.92143893,0.6910792,0.46071947,0.23035973,0.0,0.13665408,0.26940376,0.40605783,0.5388075,0.6754616,0.60127795,0.5231899,0.44900626,0.37482262,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.80821127,1.6164225,2.4207294,3.2289407,4.037152,4.802415,5.5676775,6.3329406,7.098203,7.8634663,7.168483,6.473499,5.7785153,5.083532,4.388548,3.7599394,3.1313305,2.5066261,1.8780174,1.2494087,1.3079748,1.3665408,1.4212024,1.4797685,1.5383345,1.3235924,1.1127546,0.9019169,0.6871748,0.47633708,0.58566034,0.698888,0.81211567,0.92534333,1.038571,0.8862993,0.737932,0.58566034,0.43729305,0.28892577,0.59346914,0.9019169,1.2103647,1.5188124,1.8233559,1.9717231,2.1161861,2.260649,2.4051118,2.5495746,2.9868677,3.4241607,3.8614538,4.298747,4.73604,5.743376,6.746807,7.7541428,8.757574,9.761005,9.561881,9.358852,9.155824,8.952794,8.749765,9.151918,9.550168,9.948417,10.350571,10.748819,9.440845,8.128965,6.8209906,5.5091114,4.2011366,5.0210614,5.84489,6.6687193,7.4886436,8.312472,7.7892823,7.266093,6.746807,6.223617,5.700427,5.6262436,5.5559645,5.481781,5.4115014,5.337318,5.290465,5.2436123,5.196759,5.1460023,5.099149,4.8492675,4.5993857,4.349504,4.0996222,3.8497405,3.521771,3.193801,2.8658314,2.541766,2.2137961,3.2679846,4.322173,5.376362,6.434455,7.4886436,8.503788,9.518932,10.534078,11.549222,12.564366,13.575606,14.586847,15.598087,16.613232,17.624472,16.85921,16.093946,15.328683,14.56342,13.798158,14.739119,15.676175,16.613232,17.550287,18.487345,17.034906,15.582469,14.130032,12.677594,11.225157,8.98403,6.746807,4.50568,2.2645533,0.023426414,3.0727646,6.1181984,9.167537,12.216875,15.262308,16.827974,18.393639,19.959305,21.521065,23.086731,23.551353,24.012074,24.476698,24.937418,25.398136,22.586967,19.775797,16.960724,14.149553,11.338385,11.642927,11.947471,12.252014,12.556558,12.861101,11.248583,9.636065,8.023546,6.4110284,4.7985106,4.9546866,5.1108627,5.263134,5.4193106,5.575486,5.02887,4.4861584,3.9395418,3.39683,2.8502135,3.7443218,4.6345253,5.5286336,6.4188375,7.3129454,7.066968,6.8209906,6.578918,6.3329406,6.086963,4.8687897,3.6506162,2.436347,1.2181735,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24207294,0.48414588,0.7262188,0.96829176,1.2142692,1.6749885,2.135708,2.6003318,3.0610514,3.5256753,3.0337205,2.5456703,2.0537157,1.5656652,1.0737107,0.8706817,0.6637484,0.46071947,0.25378615,0.05075723,0.58175594,1.1088502,1.639849,2.1708477,2.7018464,2.260649,1.8194515,1.3782539,0.94096094,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.21083772,0.42557985,0.63641757,0.8511597,1.0619974,1.5851873,2.1083772,2.631567,3.1508527,3.6740425,4.661856,5.645766,6.629675,7.6135845,8.601398,7.7814736,6.9615493,6.141625,5.3217,4.5017757,3.619381,2.7408905,1.8584955,0.98000497,0.10151446,1.0541886,2.0068626,2.9556324,3.9083066,4.860981,5.169429,5.473972,5.7785153,6.083059,6.387602,6.223617,6.0635366,5.899552,5.735567,5.575486,5.169429,4.7633705,4.3612175,3.9551594,3.5491016,2.8385005,2.1318035,1.4212024,0.7106012,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,1.0463798,1.9131571,2.7838387,3.6545205,4.5252023,5.4583545,6.3915067,7.320754,8.253906,9.187058,8.81614,8.449126,8.078208,7.70729,7.336372,6.3056097,5.278752,4.2479897,3.2172275,2.1864653,1.9443923,1.7023194,1.4602464,1.2181735,0.97610056,0.97219616,0.96829176,0.96829176,0.96438736,0.96438736,0.8433509,0.7262188,0.60908675,0.49195468,0.37482262,0.5309987,0.6910792,0.8472553,1.0034313,1.1635119,1.2142692,1.2689307,1.319688,1.3743496,1.4251068,1.3040704,1.183034,1.0659018,0.94486535,0.8238289,0.8160201,0.80430686,0.79649806,0.78478485,0.77307165,0.7066968,0.64032197,0.57394713,0.5036679,0.43729305,0.44900626,0.46071947,0.47633708,0.48805028,0.4997635,0.999527,1.4992905,1.999054,2.4988174,2.998581,3.240654,3.4866312,3.7287042,3.970777,4.21285,1.8233559,1.8194515,1.815547,1.8116426,1.8038338,1.7999294,1.7530766,1.7101282,1.6632754,1.620327,1.5734742,1.4641509,1.3509232,1.2376955,1.1244678,1.0112402,1.1127546,1.2142692,1.3118792,1.4133936,1.5110037,1.4992905,1.4875772,1.475864,1.4641509,1.4485333,1.4992905,1.5461433,1.5929961,1.639849,1.6867018,1.5305257,1.3743496,1.2142692,1.0580931,0.9019169,0.79259366,0.6832704,0.57785153,0.46852827,0.3631094,0.3553006,0.3474918,0.339683,0.3318742,0.3240654,0.58956474,0.8550641,1.1205635,1.3860629,1.6515622,1.6437533,1.639849,1.6359446,1.6281357,1.6242313,2.018576,2.4090161,2.803361,3.193801,3.5881457,4.173806,4.7633705,5.349031,5.938596,6.524256,6.348558,6.1767645,6.001066,5.825368,5.64967,5.606722,5.559869,5.5169206,5.4700675,5.423215,5.5247293,5.6262436,5.7238536,5.825368,5.9268827,6.2743745,6.6257706,6.9732623,7.3246584,7.676055,7.8049,7.9337454,8.066495,8.19534,8.324185,8.343708,8.36323,8.386656,8.406178,8.4257,8.827853,9.230007,9.63216,10.034314,10.436467,9.573594,8.706817,7.843944,6.9771667,6.114294,6.028397,5.9464045,5.8644123,5.7824197,5.700427,5.758993,5.8214636,5.8800297,5.938596,6.001066,8.046973,10.096785,12.142691,14.188598,16.238409,14.618082,12.997755,11.377428,9.757101,8.136774,8.566258,8.995743,9.4291315,9.858616,10.2881,9.339331,8.386656,7.437886,6.4891167,5.5364423,5.0757227,4.6110992,4.1503797,3.6857557,3.2250361,4.3534083,5.4856853,6.6140575,7.746334,8.874706,8.078208,7.28171,6.481308,5.6848097,4.8883114,5.0210614,5.1577153,5.2943697,5.4271193,5.563773,6.1884775,6.817086,7.445695,8.074304,8.699008,8.956698,9.2104845,9.464272,9.718058,9.975748,9.483793,8.995743,8.503788,8.015738,7.523783,7.2582836,6.996689,6.7311897,6.46569,6.2001905,5.493494,4.7907014,4.084005,3.3812122,2.6745155,2.893162,3.1118085,3.3265507,3.5451972,3.7638438,4.482254,5.2006636,5.9229784,6.6413884,7.363703,6.8639393,6.36808,5.8683167,5.3724575,4.8765984,4.5017757,4.1308575,3.7560349,3.3851168,3.0141985,2.803361,2.5964274,2.3894942,2.182561,1.9756275,1.9834363,1.9951496,2.0068626,2.0146716,2.0263848,2.2879796,2.5495746,2.8111696,3.076669,3.338264,3.9044023,4.466636,5.0327744,5.5989127,6.1611466,5.903456,5.645766,5.388075,5.134289,4.8765984,6.4305506,7.988407,9.546264,11.10412,12.661977,11.560935,10.4637985,9.362757,8.261715,7.1606736,7.0708723,6.9810715,6.89127,6.801469,6.7116675,7.043542,7.3715115,7.703386,8.031356,8.36323,9.362757,10.362284,11.361811,12.361338,13.360865,12.458947,11.553126,10.647305,9.741484,8.835662,7.8673706,6.899079,5.9268827,4.958591,3.9863946,4.5564375,5.12648,5.6965227,6.266566,6.8366084,7.223144,7.6135845,8.00012,8.386656,8.773191,9.062118,9.351044,9.636065,9.924991,10.213917,8.671678,7.1333427,5.591104,4.0527697,2.514435,2.1239948,1.737459,1.3509232,0.96438736,0.57394713,0.46071947,0.3435874,0.23035973,0.113227665,0.0,0.1796025,0.359205,0.5388075,0.71841,0.9019169,0.80040246,0.698888,0.60127795,0.4997635,0.39824903,0.32016098,0.23816854,0.16008049,0.078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.698888,1.3938715,2.0927596,2.7916477,3.4866312,4.2948427,5.1030536,5.911265,6.715572,7.523783,6.703859,5.8800297,5.056201,4.2362766,3.4124475,2.8814487,2.3465457,1.815547,1.2806439,0.74964523,1.0112402,1.2689307,1.5305257,1.7882162,2.0498111,1.7491722,1.4485333,1.1517987,0.8511597,0.5505207,0.58566034,0.62470436,0.6637484,0.698888,0.737932,0.62470436,0.5114767,0.39824903,0.28892577,0.1756981,0.3357786,0.4958591,0.6559396,0.8160201,0.97610056,1.2220778,1.4680552,1.717937,1.9639144,2.2137961,2.514435,2.8111696,3.1118085,3.4124475,3.7130866,4.8765984,6.044015,7.2075267,8.371038,9.538455,9.60483,9.671205,9.741484,9.807858,9.874233,10.362284,10.850334,11.338385,11.826434,12.31058,10.858143,9.4018,7.9493628,6.493021,5.036679,6.0791545,7.1216297,8.164105,9.20658,10.249056,9.218294,8.191436,7.1606736,6.1299114,5.099149,5.2201858,5.3412223,5.4583545,5.579391,5.700427,5.8956475,6.0908675,6.2860875,6.481308,6.676528,6.336845,6.001066,5.661383,5.3256044,4.985922,4.369026,3.7482262,3.1274261,2.5066261,1.8858263,2.2645533,2.6432803,3.018103,3.39683,3.775557,4.958591,6.141625,7.320754,8.503788,9.686822,10.674636,11.66245,12.650263,13.638077,14.625891,13.966047,13.310107,12.654168,11.994324,11.338385,12.525322,13.712261,14.899199,16.086138,17.273075,15.305257,13.333533,11.365715,9.393991,7.426173,5.9425,4.4588275,2.979059,1.4953861,0.011713207,3.193801,6.3719845,9.554072,12.732256,15.914344,15.18422,14.454097,13.723974,12.993851,12.263727,12.67369,13.087557,13.501423,13.911386,14.325252,13.036799,11.748346,10.4637985,9.175345,7.8868923,8.351517,8.81614,9.280765,9.749292,10.213917,8.960603,7.7111945,6.461786,5.212377,3.9629683,4.6540475,5.3412223,6.0323014,6.7233806,7.4105554,6.688241,5.9659266,5.2436123,4.521298,3.7989833,4.388548,4.9781127,5.571582,6.1611466,6.7507114,6.3915067,6.028397,5.6691923,5.309987,4.950782,3.959064,2.97125,1.979532,0.9917182,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12884527,0.25378615,0.38263142,0.5114767,0.63641757,1.3001659,1.9639144,2.6237583,3.2875066,3.951255,3.3421683,2.7330816,2.1278992,1.5188124,0.9136301,0.7340276,0.5583295,0.37872702,0.20302892,0.023426414,0.7418364,1.456342,2.1708477,2.8853533,3.5998588,2.9283018,2.260649,1.5890918,0.92143893,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.24988174,0.4997635,0.74964523,0.999527,1.2494087,1.979532,2.7096553,3.4397783,4.169902,4.900025,5.794133,6.6843367,7.578445,8.468649,9.362757,7.941554,6.5164475,5.095245,3.6740425,2.2489357,1.8233559,1.3938715,0.96829176,0.5388075,0.113227665,0.58175594,1.0541886,1.5227169,1.9912452,2.463678,2.8892577,3.3187418,3.7443218,4.173806,4.5993857,4.513489,4.423688,4.337791,4.251894,4.1620927,3.8965936,3.631094,3.3655949,3.1039999,2.8385005,2.2684577,1.7023194,1.1361811,0.5661383,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.1639849,0.1756981,0.18741131,0.19912452,0.21083772,1.2728351,2.330928,3.3929255,4.4510183,5.5130157,6.5984397,7.6838636,8.769287,9.850807,10.936231,10.690253,10.444276,10.194394,9.948417,9.698535,8.324185,6.9459314,5.5676775,4.1894236,2.8111696,2.5105307,2.2059872,1.9053483,1.6008049,1.3001659,1.2923572,1.2845483,1.2767396,1.2689307,1.261122,1.0854238,0.9058213,0.7301232,0.5544251,0.37482262,0.5466163,0.71841,0.8941081,1.0659018,1.2376955,1.358732,1.475864,1.5969005,1.717937,1.8389735,1.678893,1.5188124,1.358732,1.1986516,1.038571,1.0073358,0.97610056,0.94876975,0.91753453,0.8862993,0.76135844,0.63251317,0.5036679,0.37872702,0.24988174,0.30063897,0.3513962,0.39824903,0.44900626,0.4997635,1.0112402,1.5266213,2.0380979,2.5495746,3.0610514,3.2914112,3.5178664,3.7443218,3.970777,4.2011366,2.1239948,2.0615244,1.999054,1.9365835,1.8741131,1.8116426,1.7608855,1.7140326,1.6632754,1.6125181,1.5617609,1.4133936,1.261122,1.1127546,0.96438736,0.81211567,0.9136301,1.0112402,1.1127546,1.2142692,1.3118792,1.3001659,1.2884527,1.2767396,1.261122,1.2494087,1.175225,1.1010414,1.0268579,0.94876975,0.8745861,0.737932,0.60127795,0.46071947,0.3240654,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.5231899,0.8628729,1.1986516,1.5383345,1.8741131,1.8623998,1.8506867,1.8389735,1.8233559,1.8116426,2.2372224,2.6628022,3.0883822,3.513962,3.9356375,4.4119744,4.8883114,5.3607445,5.8370814,6.3134184,6.1767645,6.036206,5.899552,5.7628975,5.6262436,5.6379566,5.64967,5.661383,5.6730967,5.688714,5.6379566,5.5871997,5.5364423,5.4856853,5.4388323,5.9268827,6.4110284,6.899079,7.387129,7.8751793,7.687768,7.5003567,7.3129454,7.125534,6.9381227,6.4383593,5.938596,5.4388323,4.939069,4.4393053,4.9624953,5.4856853,6.012779,6.5359693,7.0630636,6.688241,6.3134184,5.938596,5.563773,5.1889505,5.001539,4.814128,4.6267166,4.4393053,4.251894,4.5993857,4.950782,5.298274,5.64967,6.001066,8.324185,10.651209,12.974329,15.3013525,17.624472,15.562947,13.501423,11.435994,9.37447,7.3129454,7.6643414,8.011833,8.36323,8.710721,9.062118,8.086017,7.113821,6.13772,5.1616197,4.1894236,3.873167,3.5608149,3.2484627,2.9361105,2.6237583,3.7482262,4.8765984,6.001066,7.125534,8.250002,7.426173,6.5984397,5.774611,4.950782,4.123049,4.1894236,4.251894,4.3143644,4.376835,4.4393053,5.22409,6.012779,6.801469,7.5862536,8.374943,8.601398,8.823949,9.050405,9.276859,9.499411,9.073831,8.648251,8.226576,7.800996,7.375416,6.9732623,6.575013,6.1767645,5.774611,5.376362,4.7633705,4.1503797,3.5373883,2.9243972,2.3114061,2.463678,2.612045,2.7643168,2.912684,3.0610514,4.025439,4.985922,5.950309,6.910792,7.8751793,7.08649,6.3017054,5.5130157,4.7243266,3.9356375,3.5998588,3.2640803,2.9243972,2.5886188,2.2489357,2.1122816,1.9756275,1.8389735,1.698415,1.5617609,1.7257458,1.8858263,2.0498111,2.2137961,2.3738766,2.6237583,2.87364,3.1235218,3.3734035,3.6232853,4.037152,4.4510183,4.860981,5.2748475,5.688714,5.5013027,5.3138914,5.12648,4.939069,4.7516575,5.2865605,5.825368,6.364176,6.899079,7.437886,7.211431,6.98888,6.7624245,6.5359693,6.3134184,6.3017054,6.2860875,6.2743745,6.262661,6.250948,6.6140575,6.9732623,7.336372,7.699481,8.062591,9.448653,10.838621,12.224684,13.610746,15.000713,14.07537,13.150026,12.224684,11.29934,10.373997,9.136301,7.898606,6.66091,5.423215,4.1894236,4.814128,5.4388323,6.0635366,6.688241,7.3129454,7.6643414,8.011833,8.36323,8.710721,9.062118,9.612638,10.163159,10.71368,11.2642,11.810817,9.811763,7.812709,5.813655,3.8106966,1.8116426,1.4485333,1.0893283,0.7262188,0.3631094,0.0,0.0,0.0,0.0,0.0,0.0,0.22645533,0.44900626,0.6754616,0.9019169,1.1244678,0.999527,0.8745861,0.74964523,0.62470436,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.0,0.0,0.0,0.0,0.0,0.58566034,1.175225,1.7608855,2.35045,2.9361105,3.78727,4.6384296,5.4856853,6.336845,7.1880045,6.239235,5.2865605,4.337791,3.3890212,2.436347,1.999054,1.5617609,1.1244678,0.6871748,0.24988174,0.7106012,1.175225,1.6359446,2.1005683,2.5612879,2.174752,1.7882162,1.4016805,1.0112402,0.62470436,0.58566034,0.5505207,0.5114767,0.47633708,0.43729305,0.3631094,0.28892577,0.21083772,0.13665408,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.47633708,0.8238289,1.175225,1.5266213,1.8741131,2.0380979,2.1981785,2.3621633,2.5261483,2.6862288,4.0137253,5.337318,6.66091,7.988407,9.311999,9.651682,9.987461,10.323239,10.662923,10.998701,11.576552,12.150499,12.724447,13.298394,13.8762455,12.27544,10.674636,9.073831,7.473026,5.8761253,7.137247,8.398369,9.663396,10.924518,12.185639,10.651209,9.112875,7.57454,6.036206,4.5017757,4.814128,5.12648,5.4388323,5.7511845,6.0635366,6.5008297,6.9381227,7.375416,7.812709,8.250002,7.824422,7.3988423,6.9732623,6.551587,6.126007,5.212377,4.298747,3.3890212,2.475391,1.5617609,1.261122,0.96438736,0.6637484,0.3631094,0.062470436,1.4133936,2.7643168,4.1113358,5.462259,6.813182,7.773665,8.738052,9.698535,10.662923,11.623405,11.076789,10.526268,9.975748,9.425227,8.874706,10.311526,11.748346,13.189071,14.625891,16.062712,13.575606,11.088503,8.601398,6.114294,3.6232853,2.900971,2.174752,1.4485333,0.7262188,0.0,3.310933,6.6257706,9.936704,13.251541,16.562475,13.536563,10.510651,7.4886436,4.462732,1.43682,1.7999294,2.1630387,2.5261483,2.8892577,3.2484627,3.4866312,3.7247996,3.9629683,4.2011366,4.4393053,5.0640097,5.688714,6.3134184,6.9381227,7.562827,6.676528,5.786324,4.900025,4.0137253,3.1235218,4.349504,5.575486,6.801469,8.023546,9.249529,8.351517,7.4495993,6.551587,5.64967,4.7516575,5.036679,5.3256044,5.610626,5.899552,6.1884775,5.7121406,5.2358036,4.7633705,4.2870336,3.8106966,3.049338,2.2879796,1.5266213,0.76135844,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.92534333,1.7882162,2.6510892,3.513962,4.376835,3.6506162,2.9243972,2.1981785,1.475864,0.74964523,0.60127795,0.44900626,0.30063897,0.14836729,0.0,0.9019169,1.7999294,2.7018464,3.5998588,4.5017757,3.5998588,2.7018464,1.7999294,0.9019169,0.0,0.0,0.0,0.0,0.0,0.0,0.28892577,0.57394713,0.8628729,1.1517987,1.43682,2.3738766,3.310933,4.251894,5.1889505,6.126007,6.9264097,7.726812,8.52331,9.323712,10.124115,8.101635,6.0752497,4.0488653,2.0263848,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.61299115,1.1635119,1.7140326,2.260649,2.8111696,2.7994564,2.787743,2.77603,2.7643168,2.7486992,2.6237583,2.4988174,2.3738766,2.2489357,2.1239948,1.698415,1.2767396,0.8511597,0.42557985,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,1.4992905,2.7486992,3.998108,5.251421,6.5008297,7.7385254,8.976221,10.213917,11.4516115,12.689307,12.564366,12.439425,12.31058,12.185639,12.0606985,10.338858,8.6131115,6.8873653,5.1616197,3.435874,3.076669,2.7135596,2.35045,1.9873407,1.6242313,1.6125181,1.6008049,1.5890918,1.5734742,1.5617609,1.3235924,1.0893283,0.8511597,0.61299115,0.37482262,0.5622339,0.74964523,0.93705654,1.1244678,1.3118792,1.4992905,1.6867018,1.8741131,2.0615244,2.2489357,2.0498111,1.8506867,1.6515622,1.4485333,1.2494087,1.1986516,1.1517987,1.1010414,1.0502841,0.999527,0.81211567,0.62470436,0.43729305,0.24988174,0.062470436,0.14836729,0.23816854,0.3240654,0.41386664,0.4997635,1.0268579,1.5500476,2.0732377,2.6003318,3.1235218,3.338264,3.5491016,3.7638438,3.9746814,4.1894236,1.737459,1.6867018,1.6320401,1.5812829,1.5266213,1.475864,1.43682,1.4016805,1.3626363,1.3235924,1.2884527,1.1908426,1.097137,1.0034313,0.9058213,0.81211567,0.9058213,1.0034313,1.097137,1.1908426,1.2884527,1.2689307,1.2494087,1.2259823,1.2064602,1.1869383,1.1010414,1.0190489,0.93315214,0.8472553,0.76135844,0.6481308,0.5309987,0.41777104,0.30063897,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.20693332,0.28502136,0.3631094,0.44510186,0.5231899,0.8394465,1.1517987,1.4641509,1.7765031,2.0888553,1.9951496,1.901444,1.8116426,1.717937,1.6242313,2.0263848,2.4285383,2.8306916,3.2367494,3.638903,4.056674,4.478349,4.8961205,5.3177958,5.735567,5.6418614,5.5442514,5.446641,5.349031,5.251421,5.196759,5.138193,5.083532,5.02887,4.9742084,4.903929,4.829746,4.755562,4.6852827,4.6110992,5.083532,5.55206,6.0205884,6.493021,6.9615493,6.8873653,6.813182,6.7389984,6.66091,6.5867267,6.1181984,5.6535745,5.185046,4.716518,4.251894,4.6735697,5.095245,5.5169206,5.938596,6.364176,6.1064854,5.8487945,5.591104,5.3334136,5.0757227,4.9156423,4.759466,4.60329,4.4432096,4.2870336,4.5837684,4.8765984,5.173333,5.466163,5.7628975,7.6643414,9.565785,11.471134,13.372578,15.274021,13.595129,11.916236,10.2334385,8.554545,6.8756523,7.141152,7.406651,7.6682463,7.9337454,8.1992445,7.3715115,6.5398736,5.708236,4.8805027,4.0488653,3.8575494,3.6662338,3.4710135,3.279698,3.0883822,3.9356375,4.786797,5.6379566,6.4891167,7.336372,6.7233806,6.114294,5.5013027,4.8883114,4.2753205,4.3534083,4.4314966,4.50568,4.5837684,4.661856,5.267039,5.872221,6.477403,7.082586,7.687768,7.7619514,7.8361354,7.914223,7.988407,8.062591,7.719003,7.3715115,7.027924,6.6843367,6.336845,6.036206,5.7316628,5.4310236,5.12648,4.825841,4.3143644,3.8067923,3.2953155,2.7838387,2.2762666,2.455869,2.6354716,2.815074,2.9946766,3.174279,3.951255,4.728231,5.5091114,6.2860875,7.0630636,6.4891167,5.919074,5.3451266,4.7711797,4.2011366,3.9161155,3.631094,3.3460727,3.0610514,2.77603,2.6432803,2.5105307,2.377781,2.2450314,2.1122816,2.233318,2.358259,2.4792955,2.6042364,2.7252727,2.9165885,3.1118085,3.3031244,3.49444,3.6857557,4.0488653,4.40807,4.7672753,5.12648,5.4856853,5.368553,5.251421,5.134289,5.017157,4.900025,5.3177958,5.735567,6.153338,6.571109,6.98888,6.824895,6.66091,6.5008297,6.336845,6.1767645,6.329036,6.481308,6.6335793,6.785851,6.9381227,7.1021075,7.266093,7.433982,7.5979667,7.7619514,9.097258,10.432563,11.767868,13.103174,14.438479,13.536563,12.630741,11.728825,10.826907,9.924991,9.054309,8.179723,7.309041,6.434455,5.563773,5.8566036,6.1494336,6.4383593,6.7311897,7.0240197,7.7970915,8.570163,9.343235,10.116306,10.889378,10.698062,10.506746,10.319335,10.128019,9.936704,8.238289,6.5437784,4.845363,3.1469483,1.4485333,1.1713207,0.8941081,0.61689556,0.339683,0.062470436,0.058566034,0.05075723,0.046852827,0.042948425,0.039044023,0.25378615,0.46852827,0.6832704,0.8980125,1.1127546,0.97219616,0.8316377,0.6910792,0.5544251,0.41386664,0.339683,0.26940376,0.19522011,0.12103647,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.76135844,1.4133936,2.0615244,2.7135596,3.3616903,3.9200199,4.478349,5.036679,5.591104,6.1494336,5.481781,4.8102236,4.138666,3.4710135,2.7994564,2.3738766,1.9443923,1.5188124,1.0893283,0.6637484,1.0541886,1.4407244,1.8311646,2.2216048,2.612045,2.4480603,2.2840753,2.1161861,1.9522011,1.7882162,1.6906061,1.5969005,1.5031948,1.4055848,1.3118792,1.0815194,0.8511597,0.62079996,0.39434463,0.1639849,0.14836729,0.13665408,0.12494087,0.113227665,0.10151446,0.40215343,0.7066968,1.0073358,1.3118792,1.6125181,1.815547,2.018576,2.2216048,2.4207294,2.6237583,3.6935644,4.759466,5.8292727,6.8951745,7.9610763,8.246098,8.531119,8.81614,9.101162,9.386183,9.96013,10.534078,11.10412,11.678067,12.24811,10.912805,9.573594,8.238289,6.899079,5.563773,6.551587,7.5433054,8.531119,9.522837,10.510651,9.483793,8.456935,7.4300776,6.4032197,5.376362,5.4271193,5.481781,5.532538,5.5832953,5.6379566,5.9151692,6.192382,6.4695945,6.746807,7.0240197,6.699954,6.375889,6.0518236,5.7238536,5.3997884,4.618908,3.8419318,3.0610514,2.280171,1.4992905,1.2767396,1.0541886,0.8316377,0.60908675,0.38653582,1.4290112,2.4714866,3.513962,4.5564375,5.5989127,7.0240197,8.449126,9.874233,11.29934,12.724447,11.62731,10.530173,9.433036,8.335898,7.238762,8.433509,9.63216,10.8308115,12.025558,13.224211,11.240774,9.253433,7.269997,5.2865605,3.2992198,4.193328,5.0913405,5.985449,6.8795567,7.773665,10.268578,12.763491,15.258404,17.753317,20.24823,16.816261,13.380386,9.944512,6.5086384,3.076669,5.5871997,8.101635,10.612165,13.1266,15.637131,13.540467,11.443803,9.343235,7.2465706,5.1499066,6.8366084,8.519405,10.206107,11.888905,13.575606,12.361338,11.143164,9.928895,8.714626,7.5003567,8.015738,8.531119,9.0465,9.561881,10.073358,9.17925,8.285142,7.3910336,6.4969254,5.5989127,5.7628975,5.9268827,6.086963,6.250948,6.4110284,5.7394714,5.067914,4.396357,3.7208953,3.049338,2.4402514,1.8311646,1.2181735,0.60908675,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.093705654,0.14055848,0.19131571,0.23816854,0.19912452,0.1639849,0.12494087,0.08589685,0.05075723,0.8160201,1.5851873,2.3543546,3.1196175,3.8887846,3.3265507,2.7682211,2.2059872,1.6476578,1.0893283,0.8902037,0.6910792,0.4958591,0.29673457,0.10151446,0.80040246,1.4992905,2.1981785,2.900971,3.5998588,2.8814487,2.1669433,1.4485333,0.7301232,0.011713207,0.14055848,0.26940376,0.39434463,0.5231899,0.6481308,0.96438736,1.2767396,1.5890918,1.901444,2.2137961,3.0532427,3.892689,4.732136,5.571582,6.4110284,6.9615493,7.5120697,8.062591,8.6131115,9.163632,7.5159745,5.8683167,4.220659,2.5730011,0.92534333,0.9136301,0.9058213,0.8941081,0.8862993,0.8745861,1.0932326,1.3157835,1.53443,1.7530766,1.9756275,2.3465457,2.7213683,3.0922866,3.4632049,3.8380275,3.6467118,3.4514916,3.260176,3.06886,2.87364,2.7057507,2.541766,2.3738766,2.2059872,2.0380979,1.6281357,1.2220778,0.8160201,0.40605783,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09761006,0.19522011,0.29283017,0.39044023,0.48805028,0.5622339,0.63641757,0.7106012,0.78868926,0.8628729,1.9287747,2.998581,4.0644827,5.134289,6.2001905,7.3012323,8.398369,9.499411,10.600452,11.701493,11.834243,11.970898,12.103647,12.240301,12.373051,10.901091,9.425227,7.9493628,6.473499,5.001539,4.5369153,4.068387,3.6037633,3.1391394,2.6745155,2.9946766,3.3148375,3.6349986,3.9551594,4.2753205,3.8458362,3.416352,2.9868677,2.5534792,2.1239948,2.2684577,2.416825,2.5612879,2.7057507,2.8502135,2.7682211,2.690133,2.6081407,2.5300527,2.4480603,2.4012074,2.35045,2.2996929,2.2489357,2.1981785,1.9756275,1.7530766,1.53443,1.3118792,1.0893283,0.95657855,0.8238289,0.6910792,0.5583295,0.42557985,0.5192855,0.61689556,0.7106012,0.80430686,0.9019169,1.3782539,1.8545911,2.330928,2.8111696,3.2875066,3.357786,3.4280653,3.4983444,3.5686235,3.638903,1.3509232,1.3079748,1.2650263,1.2220778,1.1791295,1.1361811,1.1127546,1.0893283,1.0619974,1.038571,1.0112402,0.97219616,0.93315214,0.8941081,0.8511597,0.81211567,0.9019169,0.9917182,1.0815194,1.1713207,1.261122,1.2337911,1.2064602,1.1791295,1.1517987,1.1244678,1.0307622,0.93315214,0.8394465,0.74574083,0.6481308,0.5583295,0.46462387,0.3709182,0.28111696,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.3240654,0.45681506,0.59346914,0.7262188,0.8628729,1.1517987,1.43682,1.7257458,2.0107672,2.2996929,2.1278992,1.9561055,1.7843118,1.6086137,1.43682,1.815547,2.1981785,2.5769055,2.9556324,3.338264,3.7013733,4.068387,4.4314966,4.7985106,5.1616197,5.1030536,5.0483923,4.989826,4.93126,4.8765984,4.7516575,4.630621,4.50568,4.3846436,4.263607,4.165997,4.0722914,3.978586,3.8809757,3.78727,4.240181,4.6930914,5.1460023,5.5989127,6.0518236,6.086963,6.126007,6.1611466,6.2001905,6.239235,5.801942,5.368553,4.93126,4.4978714,4.0605783,4.380739,4.7009,5.0210614,5.3412223,5.661383,5.520825,5.3841705,5.2436123,5.1030536,4.9624953,4.83365,4.7087092,4.579864,4.4510183,4.3260775,4.564246,4.806319,5.044488,5.2865605,5.5247293,7.0044975,8.484266,9.964035,11.443803,12.923572,11.62731,10.331048,9.030883,7.734621,6.4383593,6.617962,6.7975645,6.9771667,7.1567693,7.336372,6.6531014,5.9659266,5.282656,4.5993857,3.912211,3.8419318,3.767748,3.6935644,3.6232853,3.5491016,4.123049,4.7009,5.2748475,5.8487945,6.426646,6.0244927,5.6262436,5.22409,4.825841,4.423688,4.5173936,4.6110992,4.7009,4.794606,4.8883114,5.309987,5.7316628,6.153338,6.578918,7.000593,6.9264097,6.8483214,6.774138,6.699954,6.6257706,6.3602715,6.094772,5.8292727,5.563773,5.298274,5.095245,4.8883114,4.6852827,4.478349,4.2753205,3.8692627,3.4593005,3.0532427,2.6432803,2.2372224,2.4480603,2.6588979,2.8658314,3.076669,3.2875066,3.8809757,4.4705405,5.0640097,5.657479,6.250948,5.891743,5.5364423,5.1772375,4.8219366,4.462732,4.2284675,3.998108,3.7638438,3.533484,3.2992198,3.174279,3.0454338,2.9165885,2.7916477,2.6628022,2.7447948,2.8267872,2.9087796,2.9907722,3.076669,3.2094188,3.3460727,3.4788225,3.6154766,3.7482262,4.056674,4.365122,4.6735697,4.9781127,5.2865605,5.239708,5.192855,5.1460023,5.099149,5.0483923,5.349031,5.645766,5.9425,6.239235,6.5359693,6.4383593,6.336845,6.239235,6.13772,6.036206,6.356367,6.6726236,6.98888,7.309041,7.6252975,7.5940623,7.558923,7.5276875,7.4964523,7.461313,8.745861,10.0265045,11.311053,12.591698,13.8762455,12.993851,12.11536,11.23687,10.354475,9.475985,8.968412,8.460839,7.9532676,7.445695,6.9381227,6.899079,6.8561306,6.817086,6.7780423,6.7389984,7.9337454,9.128492,10.323239,11.517986,12.712734,11.783486,10.8542385,9.921086,8.991838,8.062591,6.6687193,5.270943,3.8770714,2.4831998,1.0893283,0.8941081,0.7027924,0.5114767,0.31625658,0.12494087,0.113227665,0.10541886,0.093705654,0.08589685,0.07418364,0.28111696,0.48414588,0.6910792,0.8941081,1.1010414,0.94486535,0.78868926,0.63641757,0.48024148,0.3240654,0.28111696,0.23426414,0.19131571,0.14446288,0.10151446,0.12494087,0.14836729,0.1756981,0.19912452,0.22645533,0.93705654,1.6515622,2.3621633,3.076669,3.78727,4.0527697,4.318269,4.5837684,4.8492675,5.1108627,4.7243266,4.3338866,3.9434462,3.5530062,3.1625657,2.7447948,2.3270237,1.9092526,1.4914817,1.0737107,1.3938715,1.7101282,2.0263848,2.3465457,2.6628022,2.7213683,2.77603,2.8345962,2.893162,2.951728,2.795552,2.6432803,2.4910088,2.338737,2.1864653,1.8038338,1.4172981,1.0307622,0.6481308,0.26159495,0.22645533,0.18741131,0.14836729,0.113227665,0.07418364,0.3318742,0.58566034,0.8394465,1.0932326,1.3509232,1.5929961,1.8350691,2.077142,2.3192148,2.5612879,3.3734035,4.181615,4.9937305,5.801942,6.6140575,6.844417,7.0786815,7.309041,7.5433054,7.773665,8.343708,8.913751,9.483793,10.053836,10.6238785,9.550168,8.476458,7.3988423,6.3251314,5.251421,5.9659266,6.6843367,7.4027467,8.121157,8.835662,8.320281,7.800996,7.2856145,6.7663293,6.250948,6.044015,5.833177,5.6262436,5.4193106,5.212377,5.3295093,5.446641,5.563773,5.6809053,5.801942,5.575486,5.349031,5.12648,4.900025,4.6735697,4.029343,3.3812122,2.7330816,2.084951,1.43682,1.2923572,1.1478943,1.0034313,0.8589685,0.7106012,1.4485333,2.182561,2.9165885,3.6506162,4.388548,6.2743745,8.164105,10.049932,11.935758,13.825488,12.181735,10.534078,8.890324,7.2465706,5.5989127,6.559396,7.5159745,8.472553,9.4291315,10.38571,8.905942,7.422269,5.938596,4.4588275,2.9751544,5.4895897,8.0040245,10.518459,13.036799,15.551234,17.226223,18.905115,20.58401,22.258997,23.937891,20.092054,16.246218,12.404286,8.55845,4.7126136,9.37447,14.036326,18.698183,23.363943,28.025799,23.590399,19.158901,14.727406,10.295909,5.8644123,8.609207,11.354002,14.098797,16.843592,19.588387,18.046146,16.503908,14.96167,13.415526,11.873287,11.678067,11.486752,11.291532,11.096312,10.901091,10.010887,9.120684,8.23048,7.3402762,6.4500723,6.4891167,6.524256,6.5633,6.5984397,6.6374836,5.7668023,4.8961205,4.029343,3.1586614,2.2879796,1.8311646,1.3743496,0.9136301,0.45681506,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.093705654,0.19131571,0.28502136,0.37872702,0.47633708,0.38653582,0.30063897,0.21083772,0.12494087,0.039044023,0.7106012,1.3821584,2.0537157,2.7291772,3.4007344,3.0063896,2.6081407,2.2137961,1.8194515,1.4251068,1.1791295,0.93315214,0.6910792,0.44510186,0.19912452,0.698888,1.1986516,1.698415,2.1981785,2.7018464,2.1630387,1.6281357,1.0932326,0.5583295,0.023426414,0.28111696,0.5349031,0.78868926,1.0463798,1.3001659,1.6359446,1.9756275,2.3114061,2.6510892,2.9868677,3.7287042,4.4705405,5.2162814,5.958118,6.699954,7.000593,7.3012323,7.601871,7.898606,8.1992445,6.930314,5.661383,4.388548,3.1196175,1.8506867,1.8038338,1.7608855,1.7140326,1.6710842,1.6242313,2.077142,2.5300527,2.9829633,3.435874,3.8887846,4.084005,4.279225,4.474445,4.6657605,4.860981,4.4900627,4.1191444,3.7443218,3.3734035,2.998581,2.7916477,2.5808098,2.3699722,2.1591344,1.9482968,1.5617609,1.1713207,0.78088045,0.39044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15617609,0.31625658,0.47243267,0.62860876,0.78868926,0.92534333,1.0619974,1.1986516,1.33921,1.475864,2.358259,3.2445583,4.1308575,5.0132523,5.899552,6.8639393,7.824422,8.78881,9.749292,10.71368,11.108025,11.502369,11.896713,12.291059,12.689307,11.4633255,10.237343,9.01136,7.7892823,6.5633,5.9932575,5.4271193,4.860981,4.290938,3.7247996,4.376835,5.02887,5.6809053,6.336845,6.98888,6.364176,5.743376,5.1186714,4.4978714,3.873167,3.978586,4.0801005,4.181615,4.283129,4.388548,4.041056,3.6935644,3.3460727,2.998581,2.6510892,2.7486992,2.8502135,2.951728,3.049338,3.1508527,2.7565079,2.358259,1.9639144,1.5695697,1.175225,1.097137,1.0190489,0.94096094,0.8667773,0.78868926,0.8902037,0.9917182,1.0932326,1.1986516,1.3001659,1.7296503,2.1591344,2.5886188,3.018103,3.4514916,3.377308,3.3031244,3.232845,3.1586614,3.0883822,0.96438736,0.92924774,0.8980125,0.8667773,0.8316377,0.80040246,0.78868926,0.77307165,0.76135844,0.74964523,0.737932,0.75354964,0.76916724,0.78088045,0.79649806,0.81211567,0.8980125,0.98390937,1.0659018,1.1517987,1.2376955,1.2025559,1.1674163,1.1322767,1.097137,1.0619974,0.95657855,0.8511597,0.74574083,0.6442264,0.5388075,0.46852827,0.39824903,0.3279698,0.25769055,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,0.44119745,0.62860876,0.8199245,1.0112402,1.1986516,1.4641509,1.7257458,1.9873407,2.2489357,2.514435,2.260649,2.0068626,1.7530766,1.5031948,1.2494087,1.6086137,1.9639144,2.3231194,2.67842,3.0376248,3.3460727,3.6584249,3.9668727,4.279225,4.5876727,4.5681505,4.552533,4.5369153,4.5173936,4.5017757,4.31046,4.1191444,3.9317331,3.7404175,3.5491016,3.4319696,3.3148375,3.1977055,3.0805733,2.9634414,3.39683,3.8341231,4.267512,4.7009,5.138193,5.2865605,5.4388323,5.5871997,5.735567,5.8878384,5.4856853,5.083532,4.6813784,4.279225,3.873167,4.0918136,4.31046,4.5291066,4.743849,4.9624953,4.939069,4.9156423,4.8961205,4.872694,4.8492675,4.7516575,4.6540475,4.5564375,4.4588275,4.3612175,4.548629,4.732136,4.9156423,5.1030536,5.2865605,6.3446536,7.4027467,8.460839,9.518932,10.573121,9.659492,8.745861,7.8283267,6.914696,6.001066,6.094772,6.1884775,6.2860875,6.379793,6.473499,5.9346914,5.395884,4.853172,4.3143644,3.775557,3.8224099,3.8692627,3.9161155,3.9668727,4.0137253,4.3143644,4.6110992,4.911738,5.212377,5.5130157,5.3256044,5.138193,4.950782,4.7633705,4.575959,4.6813784,4.7907014,4.8961205,5.0054436,5.1108627,5.3529353,5.591104,5.833177,6.0713453,6.3134184,6.086963,5.8644123,5.6379566,5.4115014,5.1889505,5.001539,4.8180323,4.630621,4.447114,4.263607,4.154284,4.0488653,3.9395418,3.8341231,3.7247996,3.4202564,3.1157131,2.8111696,2.5066261,2.1981785,2.4402514,2.67842,2.920493,3.1586614,3.4007344,3.8067923,4.2167544,4.6228123,5.02887,5.4388323,5.2943697,5.153811,5.009348,4.8687897,4.7243266,4.5447245,4.365122,4.185519,4.0059166,3.8263142,3.7013733,3.5803368,3.4593005,3.3343596,3.213323,3.2562714,3.2992198,3.338264,3.3812122,3.4241607,3.5022488,3.5803368,3.6584249,3.736513,3.8106966,4.068387,4.322173,4.575959,4.83365,5.087436,5.1108627,5.134289,5.153811,5.1772375,5.2006636,5.376362,5.5559645,5.7316628,5.911265,6.086963,6.0518236,6.012779,5.9737353,5.938596,5.899552,6.3836975,6.8639393,7.348085,7.8283267,8.312472,8.082112,7.8517528,7.621393,7.3910336,7.1606736,8.39056,9.6243515,10.8542385,12.084125,13.314012,12.455043,11.596075,10.741011,9.882042,9.023073,8.882515,8.741957,8.597494,8.456935,8.312472,7.941554,7.5667315,7.195813,6.8209906,6.4500723,8.066495,9.686822,11.303245,12.919667,14.53609,12.86891,11.197825,9.526741,7.8556576,6.1884775,5.095245,4.0020123,2.9087796,1.815547,0.7262188,0.61689556,0.5114767,0.40215343,0.29673457,0.18741131,0.1717937,0.15617609,0.14055848,0.12884527,0.113227665,0.30844778,0.5036679,0.698888,0.8941081,1.0893283,0.91753453,0.74574083,0.57785153,0.40605783,0.23816854,0.21864653,0.20302892,0.1835069,0.1678893,0.14836729,0.18741131,0.22645533,0.26159495,0.30063897,0.3357786,1.1127546,1.8858263,2.6628022,3.435874,4.21285,4.185519,4.1581883,4.1308575,4.1035266,4.0761957,3.9668727,3.853645,3.7443218,3.6349986,3.5256753,3.1157131,2.7096553,2.3035975,1.893635,1.4875772,1.7335546,1.9756275,2.2216048,2.4675822,2.7135596,2.9907722,3.2718892,3.5530062,3.8341231,4.1113358,3.9044023,3.6935644,3.4827268,3.2718892,3.0610514,2.522244,1.9834363,1.4407244,0.9019169,0.3631094,0.30063897,0.23816854,0.1756981,0.113227665,0.05075723,0.25769055,0.46462387,0.6715572,0.8784905,1.0893283,1.3704453,1.6515622,1.9365835,2.2177005,2.4988174,3.0532427,3.6037633,4.1581883,4.7087092,5.263134,5.4427366,5.6223392,5.801942,5.9815445,6.1611466,6.7311897,7.297328,7.8634663,8.433509,8.999647,8.187531,7.375416,6.5633,5.7511845,4.939069,5.3841705,5.8292727,6.2743745,6.715572,7.1606736,7.1567693,7.1489606,7.141152,7.1333427,7.125534,6.657006,6.1884775,5.7238536,5.2553253,4.786797,4.743849,4.7009,4.661856,4.618908,4.575959,4.4510183,4.3260775,4.2011366,4.0761957,3.951255,3.435874,2.920493,2.4051118,1.8897307,1.3743496,1.3079748,1.2415999,1.1713207,1.1049459,1.038571,1.4641509,1.893635,2.3192148,2.7486992,3.174279,5.5247293,7.8751793,10.22563,12.576079,14.92653,12.732256,10.541886,8.347612,6.153338,3.9629683,4.6813784,5.395884,6.114294,6.832704,7.551114,6.571109,5.591104,4.6110992,3.631094,2.6510892,6.785851,10.920613,15.055375,19.190138,23.3249,24.183868,25.04674,25.905708,26.764677,27.623646,23.367847,19.115953,14.860155,10.604357,6.348558,13.16174,19.974922,26.788103,33.601284,40.414467,33.644234,26.877905,20.111576,13.341343,6.575013,10.381805,14.184693,17.991486,21.794373,25.601166,23.730957,21.860748,19.99054,18.12033,16.250122,15.344301,14.438479,13.536563,12.630741,11.72492,10.838621,9.956225,9.069926,8.183627,7.3012323,7.211431,7.125534,7.0357327,6.949836,6.8639393,5.794133,4.728231,3.6584249,2.592523,1.5266213,1.2181735,0.9136301,0.60908675,0.30454338,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14055848,0.28502136,0.42557985,0.5700427,0.7106012,0.57394713,0.43729305,0.30063897,0.1639849,0.023426414,0.60127795,1.1791295,1.756981,2.3348327,2.912684,2.6823244,2.4519646,2.2216048,1.9912452,1.7608855,1.4680552,1.1791295,0.8862993,0.59346914,0.30063897,0.60127795,0.9019169,1.1986516,1.4992905,1.7999294,1.4485333,1.0932326,0.7418364,0.39044023,0.039044023,0.42167544,0.80430686,1.1869383,1.5656652,1.9482968,2.3114061,2.6745155,3.0376248,3.4007344,3.7638438,4.40807,5.0522966,5.6965227,6.3407493,6.98888,7.0357327,7.08649,7.137247,7.1880045,7.238762,6.3446536,5.45445,4.560342,3.6662338,2.77603,2.6940374,2.6159496,2.533957,2.455869,2.3738766,3.0610514,3.7443218,4.4314966,5.114767,5.801942,5.8175592,5.833177,5.852699,5.8683167,5.8878384,5.3334136,4.7828927,4.2284675,3.677947,3.1235218,2.87364,2.619854,2.366068,2.1161861,1.8623998,1.4914817,1.116659,0.74574083,0.3709182,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21864653,0.43338865,0.6520352,0.8706817,1.0893283,1.2884527,1.4875772,1.6867018,1.8858263,2.0888553,2.7916477,3.4905357,4.193328,4.8961205,5.5989127,6.426646,7.250475,8.074304,8.898132,9.725866,10.381805,11.033841,11.68978,12.34572,13.001659,12.025558,11.0494585,10.073358,9.101162,8.125061,7.453504,6.785851,6.114294,5.446641,4.775084,5.758993,6.746807,7.7307167,8.714626,9.698535,8.886419,8.070399,7.2543793,6.4383593,5.6262436,5.6848097,5.743376,5.805846,5.8644123,5.9268827,5.309987,4.6930914,4.0801005,3.4632049,2.8502135,3.1000953,3.349977,3.5998588,3.8497405,4.0996222,3.533484,2.9634414,2.397303,1.8311646,1.261122,1.2415999,1.2181735,1.1947471,1.1713207,1.1517987,1.261122,1.3704453,1.4797685,1.5890918,1.698415,2.0810463,2.463678,2.8463092,3.2289407,3.611572,3.39683,3.182088,2.9673457,2.7526035,2.5378613,0.57394713,0.5544251,0.5309987,0.5075723,0.48414588,0.46071947,0.46071947,0.46071947,0.46071947,0.46071947,0.46071947,0.5309987,0.60127795,0.6715572,0.7418364,0.81211567,0.8941081,0.97219616,1.0541886,1.1322767,1.2142692,1.1713207,1.1283722,1.0854238,1.0424755,0.999527,0.8862993,0.76916724,0.6559396,0.5388075,0.42557985,0.37872702,0.3318742,0.28111696,0.23426414,0.18741131,0.21083772,0.23816854,0.26159495,0.28892577,0.31235218,0.5583295,0.80430686,1.0463798,1.2923572,1.5383345,1.7765031,2.0107672,2.2489357,2.4871042,2.7252727,2.3933985,2.0615244,1.7257458,1.3938715,1.0619974,1.397776,1.7335546,2.069333,2.4012074,2.736986,2.9907722,3.2484627,3.5022488,3.7560349,4.0137253,4.0332475,4.056674,4.0801005,4.1035266,4.126953,3.8692627,3.611572,3.3538816,3.096191,2.8385005,2.697942,2.5573835,2.416825,2.2762666,2.135708,2.5534792,2.97125,3.3890212,3.8067923,4.224563,4.4861584,4.7516575,5.0132523,5.2748475,5.5364423,5.169429,4.7985106,4.4275923,4.056674,3.6857557,3.802888,3.9161155,4.0332475,4.1464753,4.263607,4.357313,4.4510183,4.548629,4.6423345,4.73604,4.6696653,4.60329,4.5369153,4.466636,4.4002614,4.5291066,4.661856,4.7907014,4.919547,5.0483923,5.6848097,6.321227,6.9537406,7.590158,8.226576,7.6916723,7.1606736,6.6257706,6.094772,5.563773,5.571582,5.5832953,5.591104,5.602817,5.610626,5.2162814,4.8219366,4.4275923,4.0332475,3.638903,3.8067923,3.970777,4.138666,4.3065557,4.474445,4.5017757,4.5252023,4.548629,4.575959,4.5993857,4.6267166,4.650143,4.6735697,4.7009,4.7243266,4.8492675,4.970304,5.0913405,5.2162814,5.337318,5.395884,5.45445,5.5091114,5.5676775,5.6262436,5.251421,4.8765984,4.5017757,4.123049,3.7482262,3.6467118,3.541293,3.435874,3.330455,3.2250361,3.213323,3.2055142,3.193801,3.1859922,3.174279,2.97125,2.7682211,2.5690966,2.366068,2.1630387,2.4324427,2.7018464,2.97125,3.240654,3.513962,3.736513,3.959064,4.181615,4.4041657,4.6267166,4.6969957,4.7711797,4.841459,4.9156423,4.985922,4.860981,4.732136,4.60329,4.478349,4.349504,4.2323723,4.11524,3.998108,3.8809757,3.7638438,3.7638438,3.767748,3.7716527,3.7716527,3.775557,3.795079,3.814601,3.8341231,3.853645,3.873167,4.0761957,4.279225,4.482254,4.6852827,4.8883114,4.9781127,5.0718184,5.165524,5.2592297,5.349031,5.407597,5.466163,5.520825,5.579391,5.6379566,5.661383,5.688714,5.7121406,5.735567,5.7628975,6.4110284,7.0591593,7.703386,8.351517,8.999647,8.574067,8.144583,7.719003,7.289519,6.8639393,8.039165,9.218294,10.393518,11.572648,12.751778,11.916236,11.080693,10.2451515,9.40961,8.574067,8.796618,9.019169,9.24172,9.464272,9.686822,8.98403,8.277332,7.570636,6.8678436,6.1611466,8.203149,10.241247,12.28325,14.321347,16.36335,13.954333,11.541413,9.132397,6.7233806,4.3143644,3.521771,2.7330816,1.9443923,1.1517987,0.3631094,0.339683,0.31625658,0.29673457,0.27330816,0.24988174,0.23035973,0.21083772,0.19131571,0.1717937,0.14836729,0.3357786,0.5192855,0.7066968,0.8902037,1.0737107,0.8902037,0.7066968,0.5192855,0.3357786,0.14836729,0.16008049,0.1717937,0.1796025,0.19131571,0.19912452,0.24988174,0.30063897,0.3513962,0.39824903,0.44900626,1.2884527,2.1239948,2.9634414,3.7989833,4.6384296,4.318269,3.998108,3.677947,3.357786,3.0376248,3.2094188,3.377308,3.5491016,3.716991,3.8887846,3.4905357,3.0922866,2.6940374,2.2957885,1.901444,2.0732377,2.2450314,2.416825,2.5886188,2.7643168,3.2640803,3.767748,4.271416,4.7711797,5.2748475,5.009348,4.7399445,4.4705405,4.2050414,3.9356375,3.240654,2.5456703,1.8506867,1.1557031,0.46071947,0.37482262,0.28892577,0.19912452,0.113227665,0.023426414,0.1835069,0.3435874,0.5036679,0.6637484,0.8238289,1.1478943,1.4680552,1.7921207,2.1161861,2.436347,2.7330816,3.0259118,3.3226464,3.619381,3.912211,4.041056,4.165997,4.2948427,4.423688,4.548629,5.114767,5.6809053,6.2431393,6.8092775,7.375416,6.824895,6.2743745,5.7238536,5.173333,4.6267166,4.7985106,4.970304,5.142098,5.3138914,5.4856853,5.989353,6.493021,6.996689,7.4964523,8.00012,7.2739015,6.5437784,5.8175592,5.0913405,4.3612175,4.1581883,3.959064,3.7560349,3.5530062,3.349977,3.3265507,3.2992198,3.2757936,3.2484627,3.2250361,2.8424048,2.4597735,2.077142,1.6945106,1.3118792,1.3235924,1.3314011,1.3431144,1.3509232,1.3626363,1.4836729,1.6008049,1.7218413,1.8428779,1.9639144,4.775084,7.5862536,10.401327,13.212498,16.023666,13.286681,10.545791,7.8049,5.0640097,2.3231194,2.803361,3.279698,3.7560349,4.2362766,4.7126136,4.2362766,3.7560349,3.279698,2.803361,2.3231194,8.082112,13.833297,19.588387,25.343475,31.098564,31.141512,31.184462,31.22741,31.270357,31.313307,26.647545,21.981785,17.316025,12.654168,7.988407,16.94901,25.913517,34.874123,43.838627,52.799232,43.69807,34.59691,25.491842,16.39068,7.2856145,12.154405,17.019289,21.884174,26.74906,31.613945,29.415766,27.217588,25.01941,22.821232,20.623053,19.010534,17.394112,15.781594,14.165172,12.548749,11.6702585,10.791768,9.909373,9.030883,8.148487,7.9376497,7.726812,7.5120697,7.3012323,7.08649,5.8214636,4.5564375,3.2914112,2.0263848,0.76135844,0.60908675,0.45681506,0.30454338,0.15227169,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19131571,0.37872702,0.5700427,0.76135844,0.94876975,0.76135844,0.57394713,0.38653582,0.19912452,0.011713207,0.4958591,0.97610056,1.4602464,1.9443923,2.4246337,2.358259,2.2957885,2.2294137,2.1669433,2.1005683,1.7608855,1.4212024,1.0815194,0.7418364,0.39824903,0.4997635,0.60127795,0.698888,0.80040246,0.9019169,0.7301232,0.5583295,0.39044023,0.21864653,0.05075723,0.5583295,1.0698062,1.5812829,2.0888553,2.6003318,2.9868677,3.3734035,3.7638438,4.1503797,4.5369153,5.083532,5.6340523,6.180669,6.727285,7.2739015,7.0747766,6.8756523,6.676528,6.473499,6.2743745,5.758993,5.2436123,4.728231,4.2167544,3.7013733,3.5842414,3.4710135,3.3538816,3.240654,3.1235218,4.041056,4.958591,5.8761253,6.79366,7.7111945,7.551114,7.3910336,7.230953,7.0708723,6.910792,6.180669,5.446641,4.716518,3.9824903,3.2484627,2.9556324,2.6588979,2.366068,2.069333,1.7765031,1.4212024,1.0659018,0.7106012,0.3553006,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.27721256,0.5544251,0.8316377,1.1088502,1.3860629,1.6515622,1.9131571,2.174752,2.436347,2.7018464,3.2211318,3.7404175,4.2597027,4.7789884,5.298274,5.989353,6.676528,7.363703,8.050878,8.738052,9.651682,10.569217,11.482847,12.396477,13.314012,12.587793,11.861574,11.139259,10.413041,9.686822,8.913751,8.140678,7.3715115,6.5984397,5.825368,7.141152,8.460839,9.776623,11.096312,12.412095,11.404759,10.397423,9.390087,8.382751,7.375416,7.3910336,7.4105554,7.426173,7.445695,7.461313,6.578918,5.6965227,4.814128,3.9317331,3.049338,3.4514916,3.8497405,4.251894,4.650143,5.0483923,4.31046,3.5686235,2.8306916,2.0888553,1.3509232,1.3821584,1.4133936,1.4485333,1.4797685,1.5110037,1.6281357,1.7491722,1.8663043,1.9834363,2.1005683,2.436347,2.7682211,3.1039999,3.4397783,3.775557,3.416352,3.0610514,2.7018464,2.3465457,1.9873407,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.31235218,0.43729305,0.5622339,0.6871748,0.81211567,0.8862993,0.96438736,1.038571,1.1127546,1.1869383,1.1361811,1.0893283,1.038571,0.9878138,0.93705654,0.81211567,0.6871748,0.5622339,0.43729305,0.31235218,0.28892577,0.26159495,0.23816854,0.21083772,0.18741131,0.22645533,0.26159495,0.30063897,0.3357786,0.37482262,0.6754616,0.97610056,1.2767396,1.5734742,1.8741131,2.0888553,2.2996929,2.514435,2.7252727,2.9361105,2.5261483,2.1122816,1.698415,1.2884527,0.8745861,1.1869383,1.4992905,1.8116426,2.1239948,2.436347,2.639376,2.8385005,3.0376248,3.2367494,3.435874,3.4983444,3.5608149,3.6232853,3.6857557,3.7482262,3.4241607,3.1000953,2.77603,2.4480603,2.1239948,1.9639144,1.7999294,1.6359446,1.475864,1.3118792,1.7140326,2.1122816,2.514435,2.912684,3.310933,3.6857557,4.0605783,4.4393053,4.814128,5.1889505,4.8492675,4.513489,4.173806,3.8380275,3.4983444,3.513962,3.5256753,3.5373883,3.5491016,3.5608149,3.775557,3.9863946,4.2011366,4.4119744,4.6267166,4.5876727,4.548629,4.513489,4.474445,4.4393053,4.513489,4.5876727,4.661856,4.73604,4.814128,5.024966,5.2358036,5.4505453,5.661383,5.8761253,5.7238536,5.575486,5.423215,5.2748475,5.12648,5.0483923,4.9742084,4.900025,4.825841,4.7516575,4.5017757,4.251894,3.998108,3.7482262,3.4983444,3.78727,4.0761957,4.3612175,4.650143,4.939069,4.689187,4.4393053,4.1894236,3.9356375,3.6857557,3.9239242,4.1620927,4.4002614,4.6384296,4.8765984,5.0132523,5.1499066,5.2865605,5.423215,5.563773,5.4388323,5.3138914,5.1889505,5.0640097,4.939069,4.4119744,3.8887846,3.3616903,2.8385005,2.3114061,2.2879796,2.260649,2.2372224,2.2137961,2.1864653,2.2762666,2.3621633,2.4480603,2.5378613,2.6237583,2.5261483,2.4246337,2.3231194,2.2255092,2.1239948,2.4246337,2.7252727,3.0259118,3.3265507,3.6232853,3.6623292,3.7013733,3.736513,3.775557,3.8106966,4.0996222,4.388548,4.6735697,4.9624953,5.251421,5.173333,5.099149,5.024966,4.950782,4.8765984,4.7633705,4.650143,4.5369153,4.423688,4.3143644,4.2753205,4.2362766,4.2011366,4.1620927,4.123049,4.087909,4.0488653,4.0137253,3.9746814,3.9356375,4.087909,4.2362766,4.388548,4.5369153,4.689187,4.8492675,5.0132523,5.173333,5.337318,5.5013027,5.4388323,5.376362,5.3138914,5.251421,5.1889505,5.2748475,5.3607445,5.4505453,5.5364423,5.6262436,6.4383593,7.250475,8.062591,8.874706,9.686822,9.062118,8.437413,7.812709,7.1880045,6.5633,7.687768,8.812236,9.936704,11.061172,12.185639,11.373524,10.561408,9.749292,8.937177,8.125061,8.710721,9.300286,9.885946,10.475512,11.061172,10.0265045,8.987934,7.9493628,6.910792,5.8761253,8.335898,10.799577,13.263254,15.726933,18.186707,15.035853,11.888905,8.738052,5.5871997,2.436347,1.9482968,1.4641509,0.97610056,0.48805028,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.28892577,0.26159495,0.23816854,0.21083772,0.18741131,0.3631094,0.5388075,0.7106012,0.8862993,1.0619974,0.8628729,0.6637484,0.46071947,0.26159495,0.062470436,0.10151446,0.13665408,0.1756981,0.21083772,0.24988174,0.31235218,0.37482262,0.43729305,0.4997635,0.5622339,1.4641509,2.3621633,3.2640803,4.1620927,5.0640097,4.4510183,3.8380275,3.2250361,2.612045,1.999054,2.4519646,2.900971,3.349977,3.7989833,4.251894,3.8614538,3.474918,3.0883822,2.7018464,2.3114061,2.4129205,2.514435,2.612045,2.7135596,2.8111696,3.5373883,4.263607,4.985922,5.7121406,6.4383593,6.114294,5.786324,5.462259,5.138193,4.814128,3.9629683,3.1118085,2.260649,1.4133936,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.113227665,0.22645533,0.3357786,0.44900626,0.5622339,0.92534333,1.2884527,1.6515622,2.0107672,2.3738766,2.4129205,2.4480603,2.4871042,2.5261483,2.5612879,2.639376,2.7135596,2.787743,2.8619268,2.9361105,3.4983444,4.0605783,4.6267166,5.1889505,5.7511845,5.462259,5.173333,4.8883114,4.5993857,4.3143644,4.21285,4.1113358,4.0137253,3.912211,3.8106966,4.825841,5.8370814,6.8483214,7.8634663,8.874706,7.8868923,6.899079,5.911265,4.9234514,3.9356375,3.5764325,3.213323,2.8502135,2.4871042,2.1239948,2.1981785,2.2762666,2.35045,2.4246337,2.4988174,2.2489357,1.999054,1.7491722,1.4992905,1.2494087,1.33921,1.4251068,1.5110037,1.6008049,1.6867018,1.4992905,1.3118792,1.1244678,0.93705654,0.74964523,4.025439,7.3012323,10.577025,13.848915,17.124708,13.837202,10.549695,7.262188,3.9746814,0.6871748,0.92534333,1.1635119,1.4016805,1.6359446,1.8741131,1.901444,1.9248703,1.9482968,1.9756275,1.999054,9.37447,16.749886,24.125301,31.500717,38.876133,38.099155,37.326084,36.54911,35.77604,34.99906,29.92334,24.85152,19.775797,14.700074,9.6243515,20.73628,31.84821,42.964043,54.07597,65.1879,53.748,42.312008,30.876013,19.436115,8.00012,13.927003,19.849981,25.776863,31.699842,37.626724,35.100574,32.57443,30.048279,27.526035,24.999887,22.67677,20.349745,18.026625,15.699601,13.376482,12.501896,11.623405,10.748819,9.874233,8.999647,8.663869,8.324185,7.988407,7.648724,7.3129454,5.8487945,4.388548,2.9243972,1.4641509,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23816854,0.47633708,0.7106012,0.94876975,1.1869383,0.94876975,0.7106012,0.47633708,0.23816854,0.0,0.38653582,0.77307165,1.1635119,1.5500476,1.9365835,2.0380979,2.135708,2.2372224,2.338737,2.436347,2.0498111,1.6632754,1.2767396,0.8862993,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.698888,1.33921,1.9756275,2.612045,3.2484627,3.6623292,4.0761957,4.4861584,4.900025,5.3138914,5.7628975,6.211904,6.66091,7.113821,7.562827,7.113821,6.66091,6.211904,5.7628975,5.3138914,5.173333,5.036679,4.900025,4.7633705,4.6267166,4.474445,4.3260775,4.173806,4.025439,3.873167,5.024966,6.1767645,7.3246584,8.476458,9.6243515,9.288573,8.94889,8.6131115,8.273428,7.9376497,7.0240197,6.114294,5.2006636,4.2870336,3.3734035,3.0376248,2.7018464,2.3621633,2.0263848,1.6867018,1.3509232,1.0112402,0.6754616,0.3357786,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3357786,0.6754616,1.0112402,1.3509232,1.6867018,2.0107672,2.338737,2.6628022,2.9868677,3.310933,3.6506162,3.9863946,4.3260775,4.661856,5.001539,5.548156,6.098676,6.649197,7.1997175,7.7502384,8.925464,10.100689,11.275913,12.4511385,13.626364,13.150026,12.67369,12.201257,11.72492,11.248583,10.373997,9.499411,8.624825,7.7502384,6.8756523,8.52331,10.174872,11.826434,13.4740925,15.125654,13.923099,12.724447,11.525795,10.323239,9.124588,9.101162,9.073831,9.050405,9.023073,8.999647,7.8517528,6.699954,5.548156,4.4002614,3.2484627,3.7989833,4.349504,4.900025,5.4505453,6.001066,5.087436,4.173806,3.2640803,2.35045,1.43682,1.5266213,1.6125181,1.698415,1.7882162,1.8741131,1.999054,2.1239948,2.2489357,2.3738766,2.4988174,2.787743,3.076669,3.3616903,3.6506162,3.9356375,3.435874,2.9361105,2.436347,1.9365835,1.43682,0.57394713,0.61689556,0.6559396,0.6949836,0.7340276,0.77307165,0.7418364,0.7106012,0.679366,0.6442264,0.61299115,0.6637484,0.7106012,0.76135844,0.81211567,0.8628729,0.8941081,0.92143893,0.95267415,0.98390937,1.0112402,0.97610056,0.93705654,0.9019169,0.8628729,0.8238289,0.7262188,0.62860876,0.5309987,0.43338865,0.3357786,0.32016098,0.30063897,0.28502136,0.26940376,0.24988174,0.28111696,0.31625658,0.3474918,0.37872702,0.41386664,0.6949836,0.97610056,1.261122,1.542239,1.8233559,1.9639144,2.1005683,2.2372224,2.3738766,2.514435,2.1864653,1.8623998,1.5383345,1.2142692,0.8862993,1.1283722,1.3743496,1.6164225,1.8584955,2.1005683,2.3114061,2.5261483,2.736986,2.951728,3.1625657,3.213323,3.2679846,3.3187418,3.3734035,3.4241607,3.1469483,2.8697357,2.592523,2.3153105,2.0380979,1.8506867,1.6632754,1.475864,1.2884527,1.1010414,1.4212024,1.7452679,2.069333,2.3894942,2.7135596,3.0805733,3.4475873,3.814601,4.181615,4.548629,4.3416953,4.1308575,3.9200199,3.7091823,3.4983444,3.49444,3.4905357,3.4866312,3.4788225,3.474918,3.638903,3.8067923,3.970777,4.134762,4.298747,4.357313,4.415879,4.474445,4.5291066,4.5876727,4.646239,4.7087092,4.7672753,4.825841,4.8883114,5.040583,5.196759,5.3529353,5.5091114,5.661383,5.559869,5.4583545,5.35684,5.251421,5.1499066,5.0757227,5.0054436,4.93126,4.860981,4.786797,4.5369153,4.2870336,4.037152,3.78727,3.5373883,3.7482262,3.959064,4.165997,4.376835,4.5876727,4.3729305,4.1581883,3.9434462,3.7287042,3.513962,3.775557,4.041056,4.3065557,4.572055,4.8375545,4.9468775,5.0522966,5.1616197,5.267039,5.376362,5.2592297,5.1460023,5.02887,4.9156423,4.7985106,4.3338866,3.8653584,3.39683,2.9283018,2.463678,2.475391,2.4871042,2.4988174,2.514435,2.5261483,2.5964274,2.6706111,2.7408905,2.815074,2.8892577,2.8267872,2.7682211,2.7057507,2.6471848,2.5886188,2.8111696,3.0376248,3.2640803,3.4866312,3.7130866,3.7911747,3.873167,3.951255,4.0332475,4.1113358,4.369026,4.6228123,4.8765984,5.134289,5.388075,5.3256044,5.267039,5.2084727,5.1460023,5.087436,5.0210614,4.958591,4.892216,4.825841,4.7633705,4.7204223,4.677474,4.6345253,4.591577,4.548629,4.5408196,4.5291066,4.521298,4.5095844,4.5017757,4.6150036,4.728231,4.845363,4.958591,5.0757227,5.196759,5.3138914,5.434928,5.5559645,5.6730967,5.606722,5.5364423,5.466163,5.395884,5.3256044,5.3724575,5.4193106,5.466163,5.5169206,5.563773,6.36808,7.172387,7.9766936,8.781001,9.589212,9.17925,8.769287,8.359325,7.9493628,7.5394006,8.695104,9.850807,11.010414,12.166118,13.325725,12.888432,12.4511385,12.013845,11.576552,11.139259,11.014318,10.889378,10.764437,10.6355915,10.510651,10.053836,9.597021,9.140205,8.683391,8.226576,9.550168,10.87376,12.201257,13.524849,14.848442,12.271536,9.690726,7.1099167,4.5291066,1.9482968,1.5617609,1.1713207,0.78088045,0.39044023,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.23816854,0.22645533,0.21083772,0.19912452,0.18741131,0.39824903,0.60908675,0.8160201,1.0268579,1.2376955,1.2415999,1.2415999,1.2455044,1.2494087,1.2494087,1.1596074,1.0698062,0.98000497,0.8902037,0.80040246,0.92924774,1.0580931,1.1908426,1.319688,1.4485333,1.9834363,2.514435,3.049338,3.5803368,4.1113358,3.7716527,3.4319696,3.0922866,2.7526035,2.4129205,2.8111696,3.213323,3.611572,4.0137253,4.4119744,4.1035266,3.7911747,3.4827268,3.174279,2.8619268,2.9751544,3.0883822,3.2016098,3.310933,3.4241607,3.8614538,4.298747,4.73604,5.173333,5.610626,5.4271193,5.2436123,5.056201,4.872694,4.689187,3.951255,3.2172275,2.4831998,1.7491722,1.0112402,0.8823949,0.75354964,0.62079996,0.49195468,0.3631094,0.5036679,0.6481308,0.78868926,0.93315214,1.0737107,1.3860629,1.698415,2.0107672,2.3231194,2.639376,2.6276627,2.6159496,2.6081407,2.5964274,2.5886188,2.7135596,2.8424048,2.97125,3.096191,3.2250361,3.7208953,4.2167544,4.7087092,5.2045684,5.700427,5.473972,5.2436123,5.017157,4.7907014,4.564246,4.482254,4.4041657,4.322173,4.2440853,4.1620927,5.001539,5.840986,6.6843367,7.523783,8.36323,7.4574084,6.551587,5.645766,4.743849,3.8380275,3.4788225,3.1235218,2.7643168,2.4090161,2.0498111,2.1083772,2.1708477,2.2294137,2.2918842,2.35045,2.2216048,2.0888553,1.9600099,1.8311646,1.698415,1.8663043,2.0341935,2.2020829,2.3699722,2.5378613,2.4441557,2.3543546,2.260649,2.1669433,2.0732377,4.7633705,7.4495993,10.135828,12.825961,15.51219,12.552653,9.593117,6.6335793,3.6740425,0.7106012,0.8706817,1.0268579,1.1869383,1.3431144,1.4992905,1.698415,1.893635,2.0927596,2.2918842,2.4871042,8.761478,15.031949,21.306324,27.576794,33.851166,33.741844,33.636425,33.527103,33.421684,33.31236,29.333775,25.351284,21.372698,17.394112,13.411622,21.43517,29.458715,37.478355,45.501904,53.52545,45.494095,37.466644,29.43529,21.403933,13.376482,16.870922,20.369267,23.86761,27.365955,30.8643,29.505568,28.15074,26.795912,25.441086,24.086258,22.048159,20.006157,17.96806,15.926057,13.887959,12.8767185,11.861574,10.850334,9.839094,8.823949,8.659965,8.495979,8.32809,8.164105,8.00012,6.520352,5.040583,3.5608149,2.0810463,0.60127795,0.48414588,0.3709182,0.25378615,0.14055848,0.023426414,0.023426414,0.019522011,0.015617609,0.015617609,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.27330816,0.5505207,0.8238289,1.1010414,1.3743496,1.1127546,0.8511597,0.58566034,0.3240654,0.062470436,0.359205,0.6559396,0.95657855,1.2533131,1.5500476,1.6632754,1.7804074,1.893635,2.0107672,2.1239948,1.7804074,1.43682,1.0893283,0.74574083,0.39824903,0.46852827,0.5388075,0.60908675,0.679366,0.74964523,0.64032197,0.5309987,0.42167544,0.30844778,0.19912452,0.93315214,1.6710842,2.4051118,3.1391394,3.873167,4.1620927,4.4510183,4.73604,5.024966,5.3138914,5.661383,6.008875,6.356367,6.703859,7.0513506,6.7975645,6.5437784,6.2938967,6.04011,5.786324,5.7707067,5.758993,5.743376,5.727758,5.7121406,5.423215,5.134289,4.841459,4.552533,4.263607,5.173333,6.086963,7.000593,7.914223,8.823949,8.359325,7.8947015,7.4300776,6.9654536,6.5008297,5.9073606,5.3138914,4.7243266,4.1308575,3.5373883,3.240654,2.9478238,2.6510892,2.358259,2.0615244,1.7218413,1.3821584,1.0424755,0.7027924,0.3631094,0.29283017,0.22255093,0.15227169,0.08199245,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.48414588,0.8941081,1.3040704,1.7140326,2.1239948,2.6042364,3.084478,3.5647192,4.044961,4.5252023,4.5369153,4.5447245,4.5564375,4.564246,4.575959,5.138193,5.700427,6.262661,6.824895,7.387129,8.546737,9.702439,10.858143,12.01775,13.173453,12.814248,12.4511385,12.08803,11.72492,11.361811,10.393518,9.421323,8.453031,7.480835,6.5125427,7.890797,9.269051,10.6434,12.021654,13.399908,12.73616,12.068507,11.404759,10.741011,10.073358,9.811763,9.550168,9.288573,9.023073,8.761478,8.043069,7.320754,6.602344,5.883934,5.1616197,5.3060827,5.45445,5.5989127,5.743376,5.8878384,5.036679,4.181615,3.330455,2.4792955,1.6242313,1.6749885,1.7257458,1.7765031,1.8233559,1.8741131,2.0615244,2.2489357,2.436347,2.6237583,2.8111696,2.9165885,3.0220075,3.1274261,3.232845,3.338264,2.9439192,2.5534792,2.1591344,1.7686942,1.3743496,0.96438736,1.0541886,1.1478943,1.2415999,1.3314011,1.4251068,1.3470187,1.2689307,1.1908426,1.116659,1.038571,1.0112402,0.9878138,0.96438736,0.93705654,0.9136301,0.8980125,0.8823949,0.8667773,0.8511597,0.8394465,0.81211567,0.78868926,0.76135844,0.737932,0.7106012,0.6442264,0.57394713,0.5036679,0.43338865,0.3631094,0.3513962,0.3435874,0.3318742,0.3240654,0.31235218,0.339683,0.3670138,0.39434463,0.42167544,0.44900626,0.7145056,0.98000497,1.2455044,1.5110037,1.7765031,1.8389735,1.901444,1.9639144,2.0263848,2.0888553,1.8506867,1.6125181,1.3743496,1.1361811,0.9019169,1.0737107,1.2455044,1.4172981,1.5890918,1.7608855,1.9873407,2.2137961,2.436347,2.6628022,2.8892577,2.9283018,2.97125,3.0141985,3.057147,3.1000953,2.8697357,2.639376,2.4090161,2.1786566,1.9482968,1.737459,1.5266213,1.3118792,1.1010414,0.8862993,1.1322767,1.3782539,1.6242313,1.8663043,2.1122816,2.4714866,2.8306916,3.193801,3.5530062,3.912211,3.8302186,3.7482262,3.6662338,3.5842414,3.4983444,3.4788225,3.455396,3.4319696,3.408543,3.3890212,3.506153,3.6232853,3.7404175,3.8575494,3.9746814,4.126953,4.279225,4.4314966,4.5837684,4.73604,4.7828927,4.825841,4.872694,4.9156423,4.9624953,5.0601053,5.1577153,5.2553253,5.3529353,5.4505453,5.395884,5.3412223,5.2865605,5.2318993,5.173333,5.1030536,5.036679,4.9663997,4.8961205,4.825841,4.575959,4.3260775,4.0761957,3.8263142,3.5764325,3.7091823,3.8419318,3.970777,4.1035266,4.2362766,4.056674,3.8770714,3.697469,3.5178664,3.338264,3.631094,3.9239242,4.2167544,4.50568,4.7985106,4.8765984,4.9546866,5.0327744,5.1108627,5.1889505,5.083532,4.9781127,4.872694,4.7672753,4.661856,4.251894,3.8419318,3.4319696,3.0220075,2.612045,2.6628022,2.7135596,2.7643168,2.8111696,2.8619268,2.920493,2.979059,3.0337205,3.0922866,3.1508527,3.1313305,3.1118085,3.0883822,3.06886,3.049338,3.2016098,3.349977,3.4983444,3.6506162,3.7989833,3.9239242,4.044961,4.165997,4.290938,4.4119744,4.6345253,4.8570766,5.0796275,5.3021784,5.5247293,5.481781,5.434928,5.388075,5.3451266,5.298274,5.282656,5.263134,5.2475166,5.2318993,5.212377,5.165524,5.1186714,5.0718184,5.0210614,4.9742084,4.9937305,5.009348,5.02887,5.044488,5.0640097,5.142098,5.22409,5.3021784,5.3841705,5.462259,5.5403466,5.618435,5.6965227,5.7707067,5.8487945,5.7707067,5.6965227,5.618435,5.5403466,5.462259,5.4700675,5.477876,5.4856853,5.493494,5.5013027,6.297801,7.094299,7.890797,8.691199,9.487698,9.292478,9.097258,8.902037,8.706817,8.511597,9.702439,10.893282,12.084125,13.271063,14.461906,14.399435,14.336966,14.274494,14.212025,14.149553,13.314012,12.4745655,11.639023,10.799577,9.964035,10.085071,10.206107,10.331048,10.452085,10.573121,10.764437,10.951848,11.139259,11.326671,11.514082,9.503315,7.492548,5.481781,3.4710135,1.4641509,1.1713207,0.8784905,0.58566034,0.29283017,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.43338865,0.679366,0.92143893,1.1674163,1.4133936,1.6164225,1.8233559,2.0263848,2.233318,2.436347,2.2216048,2.0029583,1.7843118,1.5656652,1.3509232,1.5461433,1.7452679,1.9443923,2.1396124,2.338737,2.5027218,2.6667068,2.8306916,2.998581,3.1625657,3.096191,3.0259118,2.959537,2.893162,2.8267872,3.174279,3.5256753,3.873167,4.224563,4.575959,4.3416953,4.1113358,3.8770714,3.6467118,3.4124475,3.5373883,3.6623292,3.78727,3.912211,4.037152,4.1894236,4.337791,4.4861584,4.6384296,4.786797,4.743849,4.6969957,4.6540475,4.607195,4.564246,3.9434462,3.3226464,2.7018464,2.0810463,1.4641509,1.3157835,1.1674163,1.0190489,0.8706817,0.7262188,0.8980125,1.0698062,1.2415999,1.4133936,1.5890918,1.8506867,2.1122816,2.3738766,2.639376,2.900971,2.8424048,2.7838387,2.7291772,2.6706111,2.612045,2.7916477,2.97125,3.1508527,3.3343596,3.513962,3.9395418,4.369026,4.794606,5.22409,5.64967,5.481781,5.3138914,5.1460023,4.9781127,4.814128,4.7516575,4.6930914,4.630621,4.572055,4.513489,5.181142,5.8487945,6.5164475,7.1841,7.8517528,7.027924,6.2040954,5.3841705,4.560342,3.736513,3.3851168,3.0337205,2.67842,2.3270237,1.9756275,2.018576,2.0654287,2.1083772,2.15523,2.1981785,2.1903696,2.1786566,2.1708477,2.1591344,2.1513257,2.397303,2.6432803,2.893162,3.1391394,3.3890212,3.3890212,3.3929255,3.39683,3.39683,3.4007344,5.5013027,7.601871,9.698535,11.799104,13.899672,11.268105,8.636538,6.001066,3.3694992,0.737932,0.8160201,0.8941081,0.96829176,1.0463798,1.1244678,1.4953861,1.8663043,2.233318,2.6042364,2.9751544,8.144583,13.314012,18.48344,23.656773,28.826202,29.384531,29.946766,30.505095,31.063425,31.625658,28.740305,25.854952,22.969599,20.084246,17.198893,22.134056,27.065317,31.996576,36.93174,41.863003,37.24019,32.61738,27.994564,23.371752,18.74894,19.818747,20.888552,21.958359,23.028164,24.101875,23.914463,23.730957,23.543545,23.360039,23.176533,21.41955,19.666473,17.909492,16.156416,14.399435,13.251541,12.099743,10.951848,9.80005,8.648251,8.65606,8.663869,8.671678,8.679486,8.687295,7.1880045,5.6926184,4.193328,2.697942,1.1986516,0.96829176,0.7418364,0.5114767,0.28111696,0.05075723,0.046852827,0.039044023,0.03513962,0.031235218,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.31235218,0.62470436,0.93705654,1.2494087,1.5617609,1.2767396,0.9878138,0.698888,0.41386664,0.12494087,0.3318742,0.5388075,0.74574083,0.95657855,1.1635119,1.2923572,1.4212024,1.5539521,1.6827974,1.8116426,1.5110037,1.2064602,0.9058213,0.60127795,0.30063897,0.5388075,0.78088045,1.0190489,1.261122,1.4992905,1.2689307,1.0346665,0.80430686,0.5700427,0.3357786,1.1713207,2.0029583,2.8345962,3.6662338,4.5017757,4.661856,4.825841,4.985922,5.1499066,5.3138914,5.5559645,5.801942,6.0479193,6.2938967,6.5359693,6.481308,6.426646,6.3719845,6.3173227,6.262661,6.36808,6.477403,6.5867267,6.6921453,6.801469,6.36808,5.938596,5.5091114,5.0796275,4.650143,5.3256044,6.001066,6.676528,7.348085,8.023546,7.433982,6.8405128,6.2470436,5.6535745,5.0640097,4.7907014,4.5173936,4.2440853,3.970777,3.7013733,3.4475873,3.193801,2.9439192,2.690133,2.436347,2.096664,1.7530766,1.4094892,1.0659018,0.7262188,0.58566034,0.44510186,0.30454338,0.1639849,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.63251317,1.116659,1.5969005,2.0810463,2.5612879,3.1977055,3.8341231,4.466636,5.1030536,5.735567,5.4193106,5.1030536,4.786797,4.466636,4.1503797,4.7243266,5.298274,5.8761253,6.4500723,7.0240197,8.164105,9.304191,10.444276,11.584361,12.724447,12.4745655,12.224684,11.974802,11.72492,11.475039,10.409137,9.343235,8.281238,7.2153354,6.1494336,7.2543793,8.359325,9.464272,10.569217,11.674163,11.545318,11.416472,11.283723,11.154878,11.0260315,10.526268,10.0265045,9.526741,9.026978,8.52331,8.234385,7.9454584,7.656533,7.363703,7.0747766,6.813182,6.5554914,6.2938967,6.036206,5.774611,4.9820175,4.1894236,3.39683,2.6042364,1.8116426,1.8233559,1.8389735,1.8506867,1.8623998,1.8741131,2.1239948,2.3738766,2.6237583,2.87364,3.1235218,3.049338,2.97125,2.893162,2.815074,2.736986,2.4519646,2.1669433,1.8819219,1.5969005,1.3118792,1.3509232,1.4953861,1.639849,1.7843118,1.9287747,2.0732377,1.9522011,1.8311646,1.7062237,1.5851873,1.4641509,1.3626363,1.261122,1.1635119,1.0619974,0.96438736,0.9019169,0.8433509,0.78088045,0.7223144,0.6637484,0.6481308,0.63641757,0.62470436,0.61299115,0.60127795,0.5583295,0.5153811,0.47243267,0.42948425,0.38653582,0.38653582,0.38263142,0.37872702,0.37872702,0.37482262,0.39824903,0.42167544,0.44119745,0.46462387,0.48805028,0.7340276,0.98390937,1.2298868,1.475864,1.7257458,1.7140326,1.698415,1.6867018,1.6749885,1.6632754,1.5110037,1.3626363,1.2142692,1.0619974,0.9136301,1.0151446,1.116659,1.2181735,1.3235924,1.4251068,1.6632754,1.901444,2.135708,2.3738766,2.612045,2.6432803,2.67842,2.7096553,2.7408905,2.77603,2.592523,2.4090161,2.2294137,2.0459068,1.8623998,1.6242313,1.3860629,1.1517987,0.9136301,0.6754616,0.8433509,1.0112402,1.1791295,1.3431144,1.5110037,1.8663043,2.2177005,2.5690966,2.9243972,3.2757936,3.3187418,3.3655949,3.408543,3.455396,3.4983444,3.4593005,3.4202564,3.3812122,3.338264,3.2992198,3.3694992,3.4397783,3.5100577,3.5803368,3.6506162,3.8965936,4.1464753,4.3924527,4.6384296,4.8883114,4.9156423,4.9468775,4.9781127,5.009348,5.036679,5.0757227,5.1186714,5.1577153,5.196759,5.2358036,5.2318993,5.22409,5.2162814,5.2084727,5.2006636,5.134289,5.0640097,4.997635,4.93126,4.860981,4.6110992,4.3612175,4.1113358,3.8614538,3.611572,3.6662338,3.7208953,3.775557,3.8341231,3.8887846,3.7443218,3.5959544,3.4514916,3.3070288,3.1625657,3.4827268,3.802888,4.123049,4.4432096,4.7633705,4.8102236,4.8570766,4.903929,4.950782,5.001539,4.903929,4.8102236,4.716518,4.618908,4.5252023,4.173806,3.8185053,3.4671092,3.1157131,2.7643168,2.8502135,2.9361105,3.0259118,3.1118085,3.2016098,3.240654,3.2836022,3.3265507,3.3694992,3.4124475,3.4319696,3.4514916,3.4710135,3.49444,3.513962,3.5881457,3.6623292,3.736513,3.8106966,3.8887846,4.0527697,4.2167544,4.380739,4.548629,4.7126136,4.903929,5.0913405,5.282656,5.473972,5.661383,5.6340523,5.602817,5.571582,5.5442514,5.5130157,5.5442514,5.571582,5.602817,5.6340523,5.661383,5.610626,5.5559645,5.505207,5.45445,5.3997884,5.446641,5.4895897,5.5364423,5.579391,5.6262436,5.6691923,5.716045,5.758993,5.805846,5.8487945,5.883934,5.919074,5.9542136,5.989353,6.0244927,5.938596,5.8566036,5.7707067,5.6848097,5.5989127,5.5676775,5.5364423,5.5013027,5.4700675,5.4388323,6.2275214,7.016211,7.8088045,8.597494,9.386183,9.405705,9.4291315,9.448653,9.468176,9.487698,10.709775,11.931853,13.153932,14.376009,15.598087,15.914344,16.226696,16.539047,16.8514,17.163752,15.613705,14.063657,12.513609,10.963562,9.413514,10.116306,10.819098,11.521891,12.220779,12.923572,11.974802,11.0260315,10.073358,9.124588,8.175818,6.735094,5.2943697,3.853645,2.416825,0.97610056,0.78088045,0.58566034,0.39044023,0.19522011,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.46852827,0.74574083,1.0268579,1.3079748,1.5890918,1.9951496,2.4012074,2.8111696,3.2172275,3.6232853,3.279698,2.9361105,2.5886188,2.2450314,1.901444,2.1669433,2.4285383,2.6940374,2.959537,3.2250361,3.0220075,2.8189783,2.6159496,2.416825,2.2137961,2.416825,2.6237583,2.8267872,3.0337205,3.2367494,3.5373883,3.8380275,4.138666,4.4393053,4.73604,4.5837684,4.4275923,4.271416,4.1191444,3.9629683,4.0996222,4.2362766,4.376835,4.513489,4.650143,4.513489,4.376835,4.2362766,4.0996222,3.9629683,4.056674,4.154284,4.2479897,4.3416953,4.4393053,3.9317331,3.4280653,2.9243972,2.416825,1.9131571,1.7491722,1.5812829,1.4172981,1.2533131,1.0893283,1.2884527,1.4914817,1.6945106,1.8975395,2.1005683,2.3114061,2.5261483,2.736986,2.951728,3.1625657,3.057147,2.951728,2.8463092,2.7408905,2.639376,2.8697357,3.1039999,3.3343596,3.5686235,3.7989833,4.1581883,4.521298,4.8805027,5.239708,5.5989127,5.493494,5.3841705,5.278752,5.169429,5.0640097,5.0210614,4.9820175,4.942973,4.903929,4.860981,5.35684,5.852699,6.348558,6.844417,7.336372,6.5984397,5.8566036,5.1186714,4.376835,3.638903,3.2914112,2.9439192,2.5964274,2.2489357,1.901444,1.9287747,1.9600099,1.9912452,2.018576,2.0498111,2.1591344,2.2684577,2.3816853,2.4910088,2.6003318,2.9283018,3.2562714,3.5842414,3.9083066,4.2362766,4.3338866,4.4314966,4.5291066,4.6267166,4.7243266,6.239235,7.7502384,9.261242,10.77615,12.287154,9.983557,7.676055,5.3724575,3.06886,0.76135844,0.76135844,0.75745404,0.75354964,0.75354964,0.74964523,1.2923572,1.8350691,2.377781,2.920493,3.4632049,7.531592,11.596075,15.664462,19.73285,23.801235,25.027218,26.2532,27.483088,28.70907,29.938957,28.146835,26.35862,24.5665,22.778282,20.986162,22.82904,24.671917,26.514795,28.357674,30.200552,28.986282,27.768108,26.55384,25.339571,24.125301,22.76657,21.411741,20.053009,18.694279,17.335546,18.32336,19.30727,20.291178,21.278992,22.262901,20.790941,19.322887,17.850927,16.382872,14.9109125,13.626364,12.337912,11.0494585,9.761005,8.476458,8.65606,8.835662,9.0152645,9.194867,9.37447,7.859562,6.3446536,4.829746,3.3148375,1.7999294,1.456342,1.1088502,0.76526284,0.42167544,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.3513962,0.698888,1.0502841,1.4016805,1.7491722,1.43682,1.1244678,0.81211567,0.4997635,0.18741131,0.30454338,0.42167544,0.5388075,0.6559396,0.77307165,0.92143893,1.0659018,1.2103647,1.3548276,1.4992905,1.2415999,0.98000497,0.71841,0.46071947,0.19912452,0.60908675,1.0190489,1.4290112,1.8389735,2.2489357,1.893635,1.5383345,1.1869383,0.8316377,0.47633708,1.4055848,2.3348327,3.2640803,4.193328,5.12648,5.1616197,5.2006636,5.2358036,5.2748475,5.3138914,5.45445,5.5989127,5.7394714,5.883934,6.0244927,6.168956,6.309514,6.453977,6.5945354,6.7389984,6.969358,7.195813,7.426173,7.656533,7.8868923,7.3168497,6.746807,6.1767645,5.606722,5.036679,5.473972,5.911265,6.348558,6.785851,7.223144,6.504734,5.786324,5.0640097,4.3455997,3.6232853,3.6740425,3.7208953,3.767748,3.814601,3.8614538,3.6506162,3.4436827,3.232845,3.0220075,2.8111696,2.4675822,2.1239948,1.7765031,1.4329157,1.0893283,0.8784905,0.6676528,0.45681506,0.24597734,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.22645533,0.78088045,1.3353056,1.8897307,2.4441557,2.998581,3.7911747,4.579864,5.368553,6.1611466,6.949836,6.3056097,5.661383,5.0132523,4.369026,3.7247996,4.3143644,4.900025,5.4856853,6.0752497,6.66091,7.785378,8.905942,10.03041,11.150972,12.27544,12.138786,11.998228,11.861574,11.72492,11.588266,10.4286585,9.269051,8.105539,6.9459314,5.786324,6.621866,7.453504,8.285142,9.116779,9.948417,10.354475,10.760532,11.166591,11.568744,11.974802,11.23687,10.498938,9.761005,9.026978,8.289046,8.4257,8.566258,8.706817,8.847376,8.987934,8.324185,7.656533,6.9927845,6.329036,5.661383,4.93126,4.1972322,3.4632049,2.7330816,1.999054,1.9756275,1.9482968,1.9248703,1.901444,1.8741131,2.1864653,2.4988174,2.8111696,3.1235218,3.435874,3.1781836,2.9165885,2.6588979,2.397303,2.135708,1.9600099,1.7843118,1.6047094,1.4290112,1.2494087,1.737459,1.9365835,2.1318035,2.330928,2.5261483,2.7252727,2.5573835,2.3894942,2.2216048,2.0537157,1.8858263,1.7140326,1.5383345,1.3626363,1.1869383,1.0112402,0.9058213,0.80430686,0.698888,0.59346914,0.48805028,0.48805028,0.48805028,0.48805028,0.48805028,0.48805028,0.47243267,0.45681506,0.44119745,0.42557985,0.41386664,0.41777104,0.42167544,0.42557985,0.43338865,0.43729305,0.45681506,0.47243267,0.48805028,0.5075723,0.5231899,0.75354964,0.98390937,1.2142692,1.4446288,1.6749885,1.5890918,1.4992905,1.4133936,1.3235924,1.2376955,1.175225,1.1127546,1.0502841,0.9878138,0.92534333,0.95657855,0.9917182,1.0229534,1.0541886,1.0893283,1.33921,1.5890918,1.8389735,2.0888553,2.338737,2.358259,2.3816853,2.4051118,2.4285383,2.4480603,2.3153105,2.1786566,2.0459068,1.9092526,1.7765031,1.5110037,1.2494087,0.9878138,0.7262188,0.46071947,0.5544251,0.6442264,0.7340276,0.8238289,0.9136301,1.2572175,1.6008049,1.9482968,2.2918842,2.639376,2.8111696,2.9829633,3.154757,3.3265507,3.4983444,3.4436827,3.3851168,3.3265507,3.2718892,3.213323,3.2367494,3.2562714,3.279698,3.3031244,3.3265507,3.6662338,4.009821,4.3534083,4.6930914,5.036679,5.0522966,5.067914,5.083532,5.099149,5.1108627,5.095245,5.0757227,5.0601053,5.040583,5.024966,5.0640097,5.1030536,5.1460023,5.185046,5.22409,5.1616197,5.095245,5.02887,4.9663997,4.900025,4.650143,4.4002614,4.1503797,3.900498,3.6506162,3.6271896,3.6037633,3.5842414,3.5608149,3.5373883,3.4280653,3.3187418,3.2094188,3.096191,2.9868677,3.3343596,3.6818514,4.029343,4.376835,4.7243266,4.743849,4.759466,4.7789884,4.794606,4.814128,4.728231,4.6423345,4.5564375,4.474445,4.388548,4.0918136,3.7989833,3.5022488,3.2094188,2.912684,3.0376248,3.1625657,3.2875066,3.4124475,3.5373883,3.5647192,3.59205,3.619381,3.6467118,3.6740425,3.736513,3.795079,3.853645,3.9161155,3.9746814,3.9746814,3.9746814,3.9746814,3.9746814,3.9746814,4.181615,4.388548,4.5993857,4.806319,5.0132523,5.169429,5.3256044,5.4856853,5.6418614,5.801942,5.786324,5.7707067,5.755089,5.7394714,5.7238536,5.801942,5.8800297,5.958118,6.036206,6.114294,6.055728,5.997162,5.938596,5.883934,5.825368,5.8956475,5.969831,6.044015,6.114294,6.1884775,6.196286,6.2079997,6.2158084,6.2275214,6.239235,6.2314262,6.223617,6.2158084,6.2079997,6.2001905,6.1064854,6.016684,5.9229784,5.8292727,5.735567,5.6652875,5.591104,5.520825,5.446641,5.376362,6.1572423,6.9381227,7.7229075,8.503788,9.288573,9.522837,9.757101,9.991365,10.22563,10.4637985,11.717112,12.974329,14.227642,15.480955,16.738173,17.425346,18.112522,18.799696,19.486872,20.174046,17.913397,15.648844,13.388195,11.123642,8.862993,10.143637,11.428185,12.708829,13.993378,15.274021,13.189071,11.100216,9.01136,6.9264097,4.8375545,3.9668727,3.096191,2.2294137,1.358732,0.48805028,0.39044023,0.29283017,0.19522011,0.09761006,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.5036679,0.8160201,1.1322767,1.4485333,1.7608855,2.3738766,2.9829633,3.59205,4.2011366,4.814128,4.3416953,3.8692627,3.39683,2.9243972,2.4480603,2.7838387,3.1157131,3.4475873,3.7794614,4.1113358,3.541293,2.97125,2.4012074,1.8311646,1.261122,1.7413634,2.2177005,2.6940374,3.174279,3.6506162,3.900498,4.1503797,4.4002614,4.650143,4.900025,4.8219366,4.743849,4.6657605,4.591577,4.513489,4.661856,4.814128,4.9624953,5.1108627,5.263134,4.8375545,4.4119744,3.9863946,3.5608149,3.1391394,3.3734035,3.6076677,3.8419318,4.0761957,4.3143644,3.9239242,3.533484,3.1430438,2.7526035,2.3621633,2.1786566,1.999054,1.815547,1.6320401,1.4485333,1.6827974,1.9131571,2.1474214,2.3816853,2.612045,2.77603,2.9361105,3.1000953,3.2640803,3.4241607,3.2718892,3.1196175,2.9673457,2.815074,2.6628022,2.9478238,3.232845,3.5178664,3.802888,4.087909,4.380739,4.6735697,4.9663997,5.2592297,5.548156,5.5013027,5.45445,5.407597,5.3607445,5.3138914,5.2943697,5.270943,5.251421,5.2318993,5.212377,5.5364423,5.8566036,6.180669,6.5008297,6.824895,6.168956,5.5091114,4.853172,4.193328,3.5373883,3.193801,2.854118,2.5105307,2.1669433,1.8233559,1.8389735,1.8545911,1.8702087,1.8858263,1.901444,2.1318035,2.358259,2.5886188,2.8189783,3.049338,3.4593005,3.8653584,4.271416,4.6813784,5.087436,5.278752,5.473972,5.6652875,5.8566036,6.0518236,6.9732623,7.898606,8.823949,9.749292,10.674636,8.699008,6.719476,4.743849,2.7643168,0.78868926,0.7066968,0.62079996,0.5388075,0.45681506,0.37482262,1.0893283,1.8038338,2.5183394,3.2367494,3.951255,6.914696,9.878138,12.845484,15.808925,18.77627,20.669905,22.563541,24.46108,26.354715,28.24835,27.553368,26.858383,26.163399,25.468416,24.773432,23.527927,22.278519,21.033014,19.783606,18.538101,20.728472,22.922745,25.11702,27.30739,29.501663,25.714394,21.931028,18.143757,14.360392,10.573121,12.728352,14.883581,17.03881,19.194042,21.349272,20.166237,18.9793,17.796265,16.609327,15.426293,14.001186,12.576079,11.150972,9.725866,8.300759,8.652155,9.0035515,9.358852,9.710248,10.061645,8.531119,6.996689,5.466163,3.9317331,2.4012074,1.9404879,1.4797685,1.0190489,0.5583295,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.38653582,0.77307165,1.1635119,1.5500476,1.9365835,1.6008049,1.261122,0.92534333,0.58566034,0.24988174,0.27721256,0.30454338,0.3318742,0.359205,0.38653582,0.5466163,0.7066968,0.8667773,1.0268579,1.1869383,0.96829176,0.75354964,0.5349031,0.31625658,0.10151446,0.679366,1.261122,1.8389735,2.4207294,2.998581,2.522244,2.0459068,1.5656652,1.0893283,0.61299115,1.639849,2.6667068,3.6935644,4.7243266,5.7511845,5.661383,5.575486,5.4856853,5.3997884,5.3138914,5.3529353,5.3919797,5.4310236,5.473972,5.5130157,5.852699,6.192382,6.532065,6.871748,7.211431,7.5667315,7.918128,8.269524,8.62092,8.976221,8.265619,7.5550184,6.844417,6.133816,5.423215,5.6262436,5.825368,6.0244927,6.223617,6.426646,5.579391,4.728231,3.8809757,3.0337205,2.1864653,2.5534792,2.9243972,3.2914112,3.6584249,4.025439,3.8575494,3.68966,3.521771,3.3538816,3.1859922,2.8385005,2.4910088,2.1435168,1.796025,1.4485333,1.1713207,0.8902037,0.60908675,0.3318742,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.30063897,0.92924774,1.5539521,2.182561,2.8111696,3.435874,4.380739,5.3256044,6.2743745,7.2192397,8.164105,7.1880045,6.2158084,5.2436123,4.271416,3.2992198,3.900498,4.5017757,5.099149,5.700427,6.3017054,7.406651,8.511597,9.616543,10.721489,11.826434,11.799104,11.775677,11.748346,11.72492,11.701493,10.444276,9.190963,7.9337454,6.6804323,5.423215,5.985449,6.5437784,7.1060123,7.6643414,8.226576,9.163632,10.104593,11.045554,11.986515,12.923572,11.951375,10.975275,9.999174,9.026978,8.050878,8.62092,9.190963,9.761005,10.331048,10.901091,9.8312845,8.761478,7.6916723,6.621866,5.548156,4.8765984,4.2050414,3.533484,2.8619268,2.1864653,2.1239948,2.0615244,1.999054,1.9365835,1.8741131,2.2489357,2.6237583,2.998581,3.3734035,3.7482262,3.3070288,2.8658314,2.4207294,1.979532,1.5383345,1.4680552,1.397776,1.3274968,1.2572175,1.1869383,2.1239948,2.3738766,2.6237583,2.87364,3.1235218,3.3734035,3.1625657,2.951728,2.736986,2.5261483,2.3114061,2.0615244,1.8116426,1.5617609,1.3118792,1.0619974,0.9136301,0.76135844,0.61299115,0.46071947,0.31235218,0.3240654,0.3357786,0.3513962,0.3631094,0.37482262,0.38653582,0.39824903,0.41386664,0.42557985,0.43729305,0.44900626,0.46071947,0.47633708,0.48805028,0.4997635,0.5114767,0.5231899,0.5388075,0.5505207,0.5622339,0.77307165,0.9878138,1.1986516,1.4133936,1.6242313,1.4641509,1.3001659,1.1361811,0.97610056,0.81211567,0.8394465,0.8628729,0.8862993,0.9136301,0.93705654,0.9019169,0.8628729,0.8238289,0.78868926,0.74964523,1.0112402,1.2767396,1.5383345,1.7999294,2.0615244,2.0732377,2.0888553,2.1005683,2.1122816,2.1239948,2.0380979,1.9482968,1.8623998,1.7765031,1.6867018,1.4016805,1.1127546,0.8238289,0.5388075,0.24988174,0.26159495,0.27330816,0.28892577,0.30063897,0.31235218,0.6481308,0.9878138,1.3235924,1.6632754,1.999054,2.2996929,2.6003318,2.900971,3.2016098,3.4983444,3.4241607,3.349977,3.2757936,3.2016098,3.1235218,3.1000953,3.076669,3.049338,3.0259118,2.998581,3.435874,3.873167,4.3143644,4.7516575,5.1889505,5.1889505,5.1889505,5.1889505,5.1889505,5.1889505,5.1108627,5.036679,4.9624953,4.8883114,4.814128,4.900025,4.985922,5.0757227,5.1616197,5.251421,5.1889505,5.12648,5.0640097,5.001539,4.939069,4.689187,4.4393053,4.1894236,3.9356375,3.6857557,3.5881457,3.4866312,3.3890212,3.2875066,3.1859922,3.1118085,3.0376248,2.9634414,2.8892577,2.8111696,3.1859922,3.5608149,3.9356375,4.3143644,4.689187,4.6735697,4.661856,4.650143,4.6384296,4.6267166,4.548629,4.474445,4.4002614,4.3260775,4.251894,4.0137253,3.775557,3.5373883,3.2992198,3.0610514,3.2250361,3.3890212,3.5491016,3.7130866,3.873167,3.8887846,3.900498,3.912211,3.9239242,3.9356375,4.037152,4.138666,4.2362766,4.337791,4.4393053,4.3612175,4.2870336,4.21285,4.138666,4.0605783,4.3143644,4.564246,4.814128,5.0640097,5.3138914,5.4388323,5.563773,5.688714,5.813655,5.938596,5.938596,5.938596,5.938596,5.938596,5.938596,6.0635366,6.1884775,6.3134184,6.4383593,6.5633,6.5008297,6.4383593,6.375889,6.3134184,6.250948,6.348558,6.4500723,6.551587,6.649197,6.7507114,6.7233806,6.699954,6.676528,6.649197,6.6257706,6.575013,6.524256,6.473499,6.426646,6.375889,6.2743745,6.1767645,6.0752497,5.9737353,5.8761253,5.7628975,5.64967,5.5364423,5.423215,5.3138914,6.086963,6.8639393,7.6370106,8.413987,9.187058,9.636065,10.088976,10.537982,10.986988,11.435994,12.724447,14.012899,15.3013525,16.585901,17.874353,18.936352,19.998348,21.06425,22.126247,23.188246,20.21309,17.237936,14.262781,11.287627,8.312472,10.174872,12.037272,13.899672,15.762072,17.624472,14.399435,11.174399,7.9493628,4.7243266,1.4992905,1.1986516,0.9019169,0.60127795,0.30063897,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.5388075,0.8862993,1.2376955,1.5890918,1.9365835,2.7486992,3.5608149,4.376835,5.1889505,6.001066,5.3997884,4.7985106,4.2011366,3.5998588,2.998581,3.4007344,3.7989833,4.2011366,4.5993857,5.001539,4.0605783,3.1235218,2.1864653,1.2494087,0.31235218,1.0619974,1.8116426,2.5612879,3.310933,4.0605783,4.263607,4.462732,4.661856,4.860981,5.0640097,5.0640097,5.0640097,5.0640097,5.0640097,5.0640097,5.22409,5.388075,5.548156,5.7121406,5.8761253,5.1616197,4.4510183,3.736513,3.0259118,2.3114061,2.6862288,3.0610514,3.435874,3.8106966,4.1894236,3.912211,3.638903,3.3616903,3.0883822,2.8111696,2.612045,2.4129205,2.2137961,2.0107672,1.8116426,2.0732377,2.338737,2.6003318,2.8619268,3.1235218,3.2367494,3.349977,3.4632049,3.5764325,3.6857557,3.4866312,3.2875066,3.0883822,2.8892577,2.6862288,3.0259118,3.3616903,3.7013733,4.037152,4.376835,4.5993857,4.825841,5.0483923,5.2748475,5.5013027,5.5130157,5.5247293,5.5364423,5.548156,5.563773,5.563773,5.563773,5.563773,5.563773,5.563773,5.7121406,5.8644123,6.012779,6.1611466,6.3134184,5.735567,5.1616197,4.5876727,4.0137253,3.435874,3.1000953,2.7643168,2.4246337,2.0888553,1.7491722,1.7491722,1.7491722,1.7491722,1.7491722,1.7491722,2.1005683,2.4480603,2.7994564,3.1508527,3.4983444,3.9863946,4.474445,4.9624953,5.4505453,5.938596,6.223617,6.5125427,6.801469,7.08649,7.375416,7.7111945,8.050878,8.386656,8.726339,9.062118,7.4105554,5.7628975,4.1113358,2.463678,0.81211567,0.6481308,0.48805028,0.3240654,0.1639849,0.0,0.8862993,1.7765031,2.6628022,3.5491016,4.4393053,6.3017054,8.164105,10.0265045,11.888905,13.751305,16.312593,18.87388,21.439074,24.00036,26.56165,26.963802,27.362051,27.764204,28.162453,28.560703,24.222912,19.889025,15.551234,11.213444,6.8756523,12.4745655,18.073479,23.676296,29.275208,34.874123,28.662216,22.450314,16.238409,10.0265045,3.8106966,7.137247,10.4637985,13.786445,17.112995,20.435642,19.537628,18.635712,17.7377,16.835783,15.93777,14.376009,12.814248,11.248583,9.686822,8.125061,8.648251,9.175345,9.698535,10.22563,10.748819,9.198771,7.648724,6.098676,4.548629,2.998581,2.4246337,1.8506867,1.2767396,0.698888,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.42557985,0.8511597,1.2767396,1.698415,2.1239948,1.7608855,1.4016805,1.038571,0.6754616,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.1756981,0.3513962,0.5231899,0.698888,0.8745861,0.698888,0.5231899,0.3513962,0.1756981,0.0,0.74964523,1.4992905,2.2489357,2.998581,3.7482262,3.1508527,2.5495746,1.9482968,1.3509232,0.74964523,1.8741131,2.998581,4.126953,5.251421,6.375889,6.1611466,5.950309,5.735567,5.5247293,5.3138914,5.251421,5.1889505,5.12648,5.0640097,5.001539,5.5364423,6.0752497,6.6140575,7.1489606,7.687768,8.164105,8.636538,9.112875,9.589212,10.061645,9.21439,8.36323,7.5120697,6.66091,5.813655,5.774611,5.735567,5.700427,5.661383,5.6262436,4.650143,3.6740425,2.7018464,1.7257458,0.74964523,1.43682,2.1239948,2.8111696,3.4983444,4.1894236,4.0605783,3.9356375,3.8106966,3.6857557,3.5608149,3.213323,2.8619268,2.514435,2.1630387,1.8116426,1.4641509,1.1127546,0.76135844,0.41386664,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.37482262,1.0737107,1.7765031,2.475391,3.174279,3.873167,4.9742084,6.0752497,7.1762915,8.273428,9.37447,8.074304,6.774138,5.473972,4.173806,2.87364,3.4866312,4.0996222,4.7126136,5.3256044,5.938596,7.0240197,8.113348,9.198771,10.2881,11.373524,11.4633255,11.549222,11.639023,11.72492,11.810817,10.4637985,9.112875,7.7619514,6.4110284,5.0640097,5.349031,5.6379566,5.9268827,6.211904,6.5008297,7.9766936,9.448653,10.924518,12.400381,13.8762455,12.661977,11.4516115,10.237343,9.026978,7.812709,8.812236,9.811763,10.81129,11.810817,12.814248,11.338385,9.86252,8.386656,6.910792,5.4388323,4.825841,4.21285,3.5998588,2.9868677,2.3738766,2.2762666,2.174752,2.0732377,1.9756275,1.8741131,2.3114061,2.7486992,3.1859922,3.6232853,4.0605783,3.435874,2.8111696,2.1864653,1.5617609,0.93705654,0.97610056,1.0112402,1.0502841,1.0893283,1.1244678,2.4012074,2.631567,2.8619268,3.0883822,3.3187418,3.5491016,3.2679846,2.9868677,2.7018464,2.4207294,2.135708,1.9600099,1.7843118,1.6047094,1.4290112,1.2494087,1.1439898,1.0346665,0.92924774,0.8199245,0.7106012,0.75354964,0.79649806,0.8394465,0.8823949,0.92534333,0.9058213,0.8862993,0.8667773,0.8433509,0.8238289,0.76916724,0.7106012,0.6520352,0.59346914,0.5388075,0.5388075,0.5388075,0.5388075,0.5388075,0.5388075,0.7106012,0.8862993,1.0619974,1.2376955,1.4133936,1.2767396,1.1361811,0.999527,0.8628729,0.7262188,0.74964523,0.77307165,0.80040246,0.8238289,0.8511597,0.8160201,0.78088045,0.74574083,0.7106012,0.6754616,0.8941081,1.116659,1.3353056,1.5539521,1.7765031,1.8350691,1.893635,1.9561055,2.0146716,2.0732377,1.9834363,1.8897307,1.796025,1.7062237,1.6125181,1.3665408,1.1205635,0.8784905,0.63251317,0.38653582,0.39824903,0.40605783,0.41777104,0.42557985,0.43729305,0.6871748,0.93705654,1.1869383,1.43682,1.6867018,1.9482968,2.2137961,2.475391,2.736986,2.998581,2.9439192,2.8892577,2.8345962,2.7799344,2.7252727,2.7213683,2.7135596,2.7096553,2.7057507,2.7018464,3.0532427,3.408543,3.7638438,4.1191444,4.474445,4.4861584,4.5017757,4.513489,4.5252023,4.5369153,4.4861584,4.4314966,4.380739,4.3260775,4.2753205,4.357313,4.4393053,4.521298,4.60329,4.689187,4.6969957,4.7087092,4.716518,4.728231,4.73604,4.533011,4.3260775,4.123049,3.9161155,3.7130866,3.5959544,3.4788225,3.3616903,3.240654,3.1235218,3.0883822,3.0532427,3.018103,2.9868677,2.951728,3.2640803,3.5803368,3.8965936,4.2089458,4.5252023,4.5095844,4.493967,4.478349,4.466636,4.4510183,4.3846436,4.318269,4.2557983,4.1894236,4.123049,3.9434462,3.7638438,3.5842414,3.4046388,3.2250361,3.416352,3.6037633,3.795079,3.9863946,4.173806,4.173806,4.169902,4.165997,4.165997,4.1620927,4.220659,4.283129,4.3416953,4.4041657,4.462732,4.3729305,4.283129,4.193328,4.1035266,4.0137253,4.1894236,4.369026,4.5447245,4.7243266,4.900025,5.0210614,5.138193,5.2592297,5.380266,5.5013027,5.520825,5.5403466,5.559869,5.579391,5.5989127,5.74728,5.8956475,6.044015,6.1884775,6.336845,6.278279,6.223617,6.165051,6.1064854,6.0518236,6.168956,6.2860875,6.4032197,6.520352,6.6374836,6.6452928,6.6531014,6.66091,6.6687193,6.676528,6.6335793,6.590631,6.547683,6.504734,6.461786,6.395411,6.329036,6.2587566,6.192382,6.126007,6.0713453,6.0205884,5.9659266,5.9151692,5.8644123,6.473499,7.082586,7.6916723,8.300759,8.913751,9.663396,10.416945,11.170495,11.924045,12.67369,14.044135,15.41458,16.785025,18.15547,19.525915,20.295082,21.06425,21.833418,22.60649,23.375656,20.623053,17.87045,15.117846,12.365242,9.612638,10.994797,12.376955,13.759113,15.141272,16.52343,13.458474,10.393518,7.328563,4.263607,1.1986516,1.1439898,1.0893283,1.0346665,0.98000497,0.92534333,0.7418364,0.5544251,0.3709182,0.1835069,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.5583295,0.92924774,1.2962615,1.6671798,2.0380979,2.8306916,3.6232853,4.415879,5.2084727,6.001066,5.3021784,4.60329,3.9083066,3.2094188,2.514435,2.8111696,3.1079042,3.4046388,3.7013733,3.998108,3.2484627,2.4988174,1.7491722,0.999527,0.24988174,0.8511597,1.4485333,2.0498111,2.6510892,3.2484627,3.408543,3.5686235,3.7287042,3.8887846,4.0488653,4.220659,4.396357,4.5681505,4.7399445,4.911738,5.056201,5.2006636,5.349031,5.493494,5.6379566,5.3060827,4.9742084,4.6384296,4.3065557,3.9746814,4.0488653,4.1191444,4.193328,4.263607,4.337791,3.959064,3.5764325,3.1977055,2.8189783,2.436347,2.3738766,2.3114061,2.2489357,2.1864653,2.1239948,2.3543546,2.5808098,2.8072653,3.0337205,3.2640803,3.3538816,3.4436827,3.533484,3.6232853,3.7130866,3.7208953,3.7287042,3.736513,3.7443218,3.7482262,4.0059166,4.2597027,4.513489,4.7711797,5.024966,5.083532,5.138193,5.196759,5.2553253,5.3138914,5.2592297,5.2084727,5.153811,5.1030536,5.0483923,5.181142,5.3138914,5.446641,5.579391,5.7121406,5.8566036,6.001066,6.1494336,6.2938967,6.4383593,5.7980375,5.1616197,4.5252023,3.8887846,3.2484627,2.9439192,2.639376,2.3348327,2.0302892,1.7257458,1.7647898,1.8038338,1.8467822,1.8858263,1.9248703,2.1669433,2.4090161,2.6510892,2.893162,3.1391394,3.5881457,4.041056,4.493967,4.9468775,5.3997884,5.6418614,5.883934,6.126007,6.36808,6.6140575,6.9615493,7.309041,7.656533,8.0040245,8.351517,6.8483214,5.349031,3.8497405,2.35045,0.8511597,0.76916724,0.6910792,0.60908675,0.5309987,0.44900626,1.0698062,1.6906061,2.3114061,2.9283018,3.5491016,5.067914,6.5867267,8.101635,9.620447,11.139259,13.606842,16.07833,18.54591,21.017397,23.488884,23.723148,23.961317,24.199486,24.437654,24.675823,21.130625,17.585428,14.040231,10.495033,6.949836,11.728825,16.503908,21.282896,26.061886,30.83697,25.612879,20.388788,15.160794,9.936704,4.7126136,7.355894,10.003078,12.6463585,15.293544,17.936825,17.261362,16.581997,15.906535,15.227169,14.551707,13.192975,11.838148,10.48332,9.128492,7.773665,8.117252,8.460839,8.804427,9.14411,9.487698,8.19534,6.902983,5.610626,4.318269,3.0259118,2.4480603,1.8741131,1.3001659,0.7262188,0.14836729,0.18741131,0.22645533,0.26159495,0.30063897,0.3357786,0.40605783,0.47633708,0.5466163,0.61689556,0.6871748,1.2064602,1.7218413,2.241127,2.7565079,3.2757936,2.9556324,2.6354716,2.3153105,1.9951496,1.6749885,1.5383345,1.4016805,1.261122,1.1244678,0.9878138,0.999527,1.0112402,1.0268579,1.038571,1.0502841,0.8394465,0.62860876,0.42167544,0.21083772,0.0,0.61299115,1.2259823,1.8389735,2.4480603,3.0610514,2.7018464,2.338737,1.9756275,1.6125181,1.2494087,2.9361105,4.618908,6.3056097,7.988407,9.675109,8.909846,8.144583,7.37932,6.6140575,5.8487945,5.786324,5.7238536,5.661383,5.5989127,5.5364423,5.872221,6.2079997,6.5437784,6.8756523,7.211431,7.558923,7.90251,8.246098,8.59359,8.937177,8.234385,7.531592,6.8287997,6.126007,5.423215,5.298274,5.173333,5.0483923,4.9234514,4.7985106,4.0761957,3.349977,2.6237583,1.901444,1.175225,1.7686942,2.366068,2.959537,3.5569105,4.1503797,3.970777,3.795079,3.619381,3.4397783,3.2640803,2.9361105,2.612045,2.2879796,1.9639144,1.6359446,1.3314011,1.0268579,0.7223144,0.41777104,0.113227665,0.28892577,0.46071947,0.63641757,0.81211567,0.9878138,1.5890918,2.194274,2.795552,3.39683,3.998108,5.0640097,6.1299114,7.195813,8.261715,9.323712,8.187531,7.0513506,5.911265,4.775084,3.638903,4.056674,4.4705405,4.8883114,5.3060827,5.7238536,6.817086,7.910319,9.0035515,10.096785,11.186112,11.478943,11.771772,12.064603,12.357433,12.650263,11.2642,9.878138,8.495979,7.1099167,5.7238536,5.7394714,5.755089,5.7707067,5.786324,5.801942,7.027924,8.253906,9.483793,10.709775,11.935758,10.924518,9.913278,8.898132,7.8868923,6.8756523,7.6643414,8.449126,9.237816,10.0265045,10.81129,9.589212,8.367134,7.1450562,5.9229784,4.7009,4.3260775,3.951255,3.5764325,3.2016098,2.8267872,2.639376,2.4480603,2.260649,2.0732377,1.8858263,2.2020829,2.5183394,2.8306916,3.1469483,3.4632049,2.97125,2.4792955,1.9834363,1.4914817,0.999527,1.0073358,1.0151446,1.0229534,1.0307622,1.038571,2.6745155,2.8853533,3.096191,3.3031244,3.513962,3.7247996,3.3734035,3.018103,2.6667068,2.3153105,1.9639144,1.8584955,1.7530766,1.6476578,1.542239,1.43682,1.3743496,1.3079748,1.2415999,1.1791295,1.1127546,1.1869383,1.2572175,1.3314011,1.4016805,1.475864,1.4212024,1.3704453,1.3157835,1.2650263,1.2142692,1.0854238,0.95657855,0.8316377,0.7027924,0.57394713,0.5622339,0.5505207,0.5388075,0.5231899,0.5114767,0.6481308,0.78868926,0.92534333,1.0619974,1.1986516,1.0893283,0.97610056,0.8628729,0.74964523,0.63641757,0.6637484,0.6871748,0.7106012,0.737932,0.76135844,0.7301232,0.698888,0.6637484,0.63251317,0.60127795,0.77697605,0.95657855,1.1322767,1.3118792,1.4875772,1.5969005,1.7023194,1.8116426,1.9170616,2.0263848,1.9287747,1.8311646,1.7335546,1.6359446,1.5383345,1.3353056,1.1322767,0.92924774,0.7262188,0.5231899,0.5309987,0.5388075,0.5466163,0.5544251,0.5622339,0.7262188,0.8862993,1.0502841,1.2142692,1.3743496,1.6008049,1.8233559,2.0498111,2.2762666,2.4988174,2.463678,2.4285383,2.3933985,2.358259,2.3231194,2.338737,2.3543546,2.3699722,2.3855898,2.4012074,2.6706111,2.9439192,3.2172275,3.4905357,3.7638438,3.78727,3.8106966,3.8380275,3.8614538,3.8887846,3.8575494,3.8263142,3.7989833,3.767748,3.736513,3.814601,3.892689,3.970777,4.0488653,4.126953,4.2089458,4.290938,4.3729305,4.454923,4.5369153,4.376835,4.2167544,4.056674,3.8965936,3.736513,3.6037633,3.4671092,3.3343596,3.1977055,3.0610514,3.06886,3.0727646,3.076669,3.0805733,3.0883822,3.3421683,3.5959544,3.853645,4.1074314,4.3612175,4.3455997,4.3260775,4.31046,4.290938,4.2753205,4.220659,4.165997,4.1113358,4.056674,3.998108,3.8770714,3.7560349,3.631094,3.5100577,3.3890212,3.6037633,3.8224099,4.041056,4.2557983,4.474445,4.4588275,4.4393053,4.423688,4.4041657,4.388548,4.40807,4.4275923,4.447114,4.466636,4.4861584,4.380739,4.279225,4.173806,4.068387,3.9629683,4.068387,4.173806,4.279225,4.380739,4.4861584,4.60329,4.716518,4.83365,4.9468775,5.0640097,5.1030536,5.142098,5.181142,5.22409,5.263134,5.4310236,5.602817,5.7707067,5.9425,6.114294,6.0596323,6.008875,5.9542136,5.903456,5.8487945,5.985449,6.1181984,6.2548523,6.3915067,6.524256,6.5633,6.606249,6.6452928,6.6843367,6.7233806,6.688241,6.6531014,6.621866,6.5867267,6.551587,6.5164475,6.481308,6.446168,6.4110284,6.375889,6.3836975,6.3915067,6.3993154,6.4032197,6.4110284,6.8561306,7.3012323,7.746334,8.191436,8.636538,9.690726,10.748819,11.803008,12.857197,13.911386,15.363823,16.816261,18.268698,19.721136,21.173573,21.653814,22.130152,22.60649,23.086731,23.563068,21.033014,18.502962,15.97291,13.442857,10.912805,11.814721,12.716639,13.618555,14.524376,15.426293,12.521418,9.616543,6.7116675,3.8067923,0.9019169,1.0893283,1.2806439,1.4680552,1.6593709,1.8506867,1.4797685,1.1088502,0.7418364,0.3709182,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.57785153,0.96829176,1.358732,1.7491722,2.135708,2.9087796,3.6818514,4.454923,5.2279944,6.001066,5.2045684,4.4119744,3.6154766,2.8189783,2.0263848,2.2216048,2.416825,2.6081407,2.803361,2.998581,2.436347,1.8741131,1.3118792,0.74964523,0.18741131,0.63641757,1.0893283,1.5383345,1.9873407,2.436347,2.5573835,2.67842,2.7994564,2.9165885,3.0376248,3.3812122,3.7287042,4.0722914,4.415879,4.7633705,4.8883114,5.017157,5.1460023,5.270943,5.3997884,5.446641,5.493494,5.5442514,5.591104,5.6379566,5.407597,5.1772375,4.9468775,4.716518,4.4861584,4.0020123,3.5178664,3.0337205,2.5456703,2.0615244,2.135708,2.2137961,2.2879796,2.3621633,2.436347,2.631567,2.822883,3.0141985,3.2094188,3.4007344,3.4671092,3.533484,3.6037633,3.6701381,3.736513,3.951255,4.165997,4.380739,4.5993857,4.814128,4.985922,5.1577153,5.3295093,5.5013027,5.6730967,5.563773,5.45445,5.3451266,5.2358036,5.12648,5.009348,4.8883114,4.7711797,4.6540475,4.5369153,4.802415,5.067914,5.3334136,5.5989127,5.8644123,6.001066,6.141625,6.282183,6.422742,6.5633,5.860508,5.1616197,4.462732,3.7638438,3.0610514,2.7916477,2.5183394,2.2450314,1.9717231,1.698415,1.7804074,1.8584955,1.9404879,2.018576,2.1005683,2.233318,2.3699722,2.5066261,2.639376,2.77603,3.193801,3.611572,4.029343,4.4432096,4.860981,5.0601053,5.2592297,5.45445,5.6535745,5.8487945,6.2079997,6.5633,6.9225054,7.28171,7.6370106,6.2860875,4.939069,3.5881457,2.2372224,0.8862993,0.8902037,0.8941081,0.8941081,0.8980125,0.9019169,1.2533131,1.6047094,1.9561055,2.3114061,2.6628022,3.8341231,5.009348,6.180669,7.3519893,8.52331,10.901091,13.2788725,15.656653,18.034433,20.412214,20.486399,20.560583,20.63867,20.712854,20.787037,18.034433,15.281831,12.529227,9.776623,7.0240197,10.979179,14.934339,18.889498,22.844658,26.799816,22.563541,18.32336,14.087084,9.850807,5.610626,7.578445,9.542359,11.506273,13.4740925,15.438006,14.981192,14.528281,14.0714655,13.618555,13.16174,12.013845,10.865952,9.718058,8.574067,7.426173,7.5862536,7.746334,7.9064145,8.066495,8.226576,7.1880045,6.153338,5.1186714,4.084005,3.049338,2.475391,1.901444,1.3235924,0.74964523,0.1756981,0.26159495,0.3513962,0.43729305,0.5231899,0.61299115,0.76526284,0.91753453,1.0698062,1.2220778,1.3743496,1.9834363,2.5964274,3.2055142,3.814601,4.423688,4.1464753,3.8692627,3.59205,3.3148375,3.0376248,2.8267872,2.612045,2.4012074,2.1864653,1.9756275,1.8233559,1.6749885,1.5266213,1.3743496,1.2259823,0.98000497,0.7340276,0.48805028,0.24597734,0.0,0.47633708,0.94876975,1.4251068,1.901444,2.3738766,2.2489357,2.1239948,1.999054,1.8741131,1.7491722,3.9942036,6.239235,8.484266,10.729298,12.974329,11.6585455,10.338858,9.023073,7.703386,6.387602,6.3251314,6.262661,6.2001905,6.13772,6.0752497,6.2079997,6.3407493,6.473499,6.606249,6.7389984,6.9537406,7.168483,7.3832245,7.5979667,7.812709,7.2582836,6.703859,6.1494336,5.591104,5.036679,4.825841,4.6110992,4.4002614,4.1894236,3.9746814,3.4983444,3.0259118,2.5495746,2.0732377,1.6008049,2.1044729,2.6042364,3.1079042,3.611572,4.1113358,3.8809757,3.6506162,3.4241607,3.193801,2.9634414,2.6628022,2.3621633,2.0615244,1.7608855,1.4641509,1.2025559,0.94096094,0.6832704,0.42167544,0.1639849,0.44900626,0.737932,1.0268579,1.3118792,1.6008049,2.1044729,2.6081407,3.1157131,3.619381,4.123049,5.153811,6.184573,7.2153354,8.246098,9.276859,8.300759,7.3246584,6.348558,5.376362,4.4002614,4.6228123,4.845363,5.067914,5.290465,5.5130157,6.610153,7.70729,8.804427,9.901564,10.998701,11.498465,11.994324,12.494087,12.989946,13.4858055,12.068507,10.647305,9.226103,7.8088045,6.387602,6.1299114,5.872221,5.6145306,5.35684,5.099149,6.0791545,7.0591593,8.039165,9.019169,9.999174,9.187058,8.374943,7.562827,6.7507114,5.938596,6.5125427,7.08649,7.6643414,8.238289,8.812236,7.843944,6.871748,5.903456,4.93126,3.9629683,3.8263142,3.6857557,3.5491016,3.4124475,3.2757936,2.998581,2.7252727,2.4480603,2.174752,1.901444,2.0927596,2.2840753,2.4792955,2.6706111,2.8619268,2.5027218,2.1435168,1.7843118,1.4212024,1.0619974,1.038571,1.0190489,0.9956226,0.97219616,0.94876975,2.951728,3.1391394,3.330455,3.521771,3.7091823,3.900498,3.4788225,3.0532427,2.631567,2.2098918,1.7882162,1.7530766,1.7218413,1.6906061,1.6593709,1.6242313,1.6008049,1.5812829,1.5578566,1.53443,1.5110037,1.6164225,1.717937,1.8194515,1.9209659,2.0263848,1.9404879,1.8545911,1.7686942,1.6867018,1.6008049,1.4016805,1.2064602,1.0073358,0.80821127,0.61299115,0.58566034,0.5622339,0.5388075,0.5114767,0.48805028,0.58566034,0.6871748,0.78868926,0.8862993,0.9878138,0.9019169,0.81211567,0.7262188,0.63641757,0.5505207,0.57394713,0.60127795,0.62470436,0.6481308,0.6754616,0.6442264,0.61689556,0.58566034,0.5544251,0.5231899,0.659844,0.79649806,0.92924774,1.0659018,1.1986516,1.3548276,1.5110037,1.6632754,1.8194515,1.9756275,1.8741131,1.7686942,1.6671798,1.5656652,1.4641509,1.3040704,1.1439898,0.98390937,0.8238289,0.6637484,0.6676528,0.6715572,0.679366,0.6832704,0.6871748,0.76135844,0.8394465,0.9136301,0.9878138,1.0619974,1.2494087,1.43682,1.6242313,1.8116426,1.999054,1.9834363,1.9717231,1.9561055,1.9404879,1.9248703,1.9600099,1.9951496,2.0302892,2.0654287,2.1005683,2.2918842,2.4792955,2.6706111,2.8619268,3.049338,3.0883822,3.1235218,3.1625657,3.2016098,3.2367494,3.2289407,3.2211318,3.213323,3.2094188,3.2016098,3.2718892,3.3460727,3.416352,3.4905357,3.5608149,3.716991,3.873167,4.029343,4.181615,4.337791,4.220659,4.1074314,3.9942036,3.8770714,3.7638438,3.611572,3.4593005,3.3031244,3.1508527,2.998581,3.0454338,3.0883822,3.135235,3.1781836,3.2250361,3.4202564,3.6154766,3.8106966,4.0059166,4.2011366,4.181615,4.1581883,4.138666,4.1191444,4.0996222,4.056674,4.009821,3.9668727,3.9200199,3.873167,3.8106966,3.7443218,3.6818514,3.6154766,3.5491016,3.795079,4.041056,4.283129,4.5291066,4.775084,4.743849,4.7087092,4.677474,4.646239,4.6110992,4.591577,4.572055,4.552533,4.533011,4.513489,4.3924527,4.271416,4.154284,4.0332475,3.912211,3.9434462,3.978586,4.009821,4.041056,4.0761957,4.185519,4.2948427,4.4041657,4.513489,4.6267166,4.6852827,4.743849,4.806319,4.8648853,4.9234514,5.1186714,5.309987,5.5013027,5.6965227,5.8878384,5.840986,5.794133,5.743376,5.6965227,5.64967,5.801942,5.9542136,6.1064854,6.2587566,6.4110284,6.4852123,6.559396,6.629675,6.703859,6.774138,6.746807,6.719476,6.6921453,6.6648145,6.6374836,6.6335793,6.6335793,6.629675,6.6257706,6.6257706,6.6921453,6.75852,6.8287997,6.8951745,6.9615493,7.2426662,7.523783,7.800996,8.082112,8.36323,9.718058,11.076789,12.435521,13.794253,15.14908,16.683512,18.221846,19.756275,21.290705,22.825136,23.008642,23.196054,23.37956,23.563068,23.750479,21.442978,19.135475,16.827974,14.520472,12.212971,12.634645,13.056321,13.481901,13.903577,14.325252,11.580457,8.835662,6.0908675,3.3460727,0.60127795,1.0346665,1.4680552,1.9053483,2.338737,2.77603,2.2216048,1.6632754,1.1088502,0.5544251,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.59737355,1.0073358,1.4172981,1.8272603,2.2372224,2.9907722,3.7443218,4.493967,5.2475166,6.001066,5.1069584,4.2167544,3.3226464,2.4285383,1.5383345,1.6281357,1.7218413,1.815547,1.9092526,1.999054,1.6242313,1.2494087,0.8745861,0.4997635,0.12494087,0.42557985,0.7262188,1.0268579,1.3235924,1.6242313,1.7062237,1.7843118,1.8663043,1.9443923,2.0263848,2.541766,3.0610514,3.5764325,4.095718,4.6110992,4.7243266,4.83365,4.942973,5.0522966,5.1616197,5.591104,6.016684,6.446168,6.871748,7.3012323,6.7663293,6.2353306,5.704332,5.169429,4.6384296,4.0488653,3.4593005,2.8658314,2.2762666,1.6867018,1.901444,2.1122816,2.3231194,2.5378613,2.7486992,2.9087796,3.0649557,3.2211318,3.3812122,3.5373883,3.5842414,3.6271896,3.6740425,3.716991,3.7638438,4.185519,4.607195,5.02887,5.45445,5.8761253,5.9659266,6.055728,6.1455293,6.2353306,6.3251314,6.0479193,5.7707067,5.493494,5.2162814,4.939069,4.755562,4.572055,4.388548,4.2089458,4.025439,4.423688,4.8219366,5.2162814,5.6145306,6.012779,6.1494336,6.282183,6.4188375,6.551587,6.688241,5.9268827,5.1616197,4.4002614,3.638903,2.87364,2.6354716,2.3933985,2.15523,1.9131571,1.6749885,1.796025,1.9131571,2.0341935,2.15523,2.2762666,2.3035975,2.330928,2.358259,2.3855898,2.4129205,2.795552,3.1781836,3.5608149,3.9434462,4.3260775,4.478349,4.630621,4.7828927,4.9351645,5.087436,5.45445,5.8214636,6.1884775,6.559396,6.9264097,5.7238536,4.5252023,3.3265507,2.1239948,0.92534333,1.0112402,1.0932326,1.1791295,1.2650263,1.3509232,1.43682,1.5188124,1.6047094,1.6906061,1.7765031,2.6042364,3.4280653,4.2557983,5.083532,5.911265,8.1992445,10.48332,12.767395,15.051471,17.335546,17.24965,17.163752,17.073952,16.988054,16.898252,14.938243,12.978233,11.018223,9.058213,7.098203,10.2334385,13.364769,16.4961,19.631334,22.762665,19.514202,16.261835,13.013372,9.761005,6.5125427,7.7970915,9.081639,10.366188,11.650736,12.939189,12.704925,12.470661,12.240301,12.006037,11.775677,10.834716,9.893755,8.956698,8.015738,7.0747766,7.0513506,7.0318284,7.008402,6.984976,6.9615493,6.184573,5.407597,4.630621,3.853645,3.076669,2.4988174,1.9248703,1.3509232,0.77307165,0.19912452,0.3357786,0.47633708,0.61299115,0.74964523,0.8862993,1.1205635,1.358732,1.5929961,1.8272603,2.0615244,2.7643168,3.4671092,4.169902,4.872694,5.575486,5.3412223,5.1069584,4.8687897,4.6345253,4.4002614,4.1113358,3.8263142,3.5373883,3.2484627,2.9634414,2.6510892,2.338737,2.0263848,1.7140326,1.4016805,1.1205635,0.8394465,0.5583295,0.28111696,0.0,0.3357786,0.6754616,1.0112402,1.3509232,1.6867018,1.7999294,1.9131571,2.0263848,2.135708,2.2489357,5.056201,7.859562,10.666827,13.470188,16.273548,14.40334,12.533132,10.666827,8.796618,6.9264097,6.8639393,6.801469,6.7389984,6.676528,6.6140575,6.5437784,6.473499,6.4032197,6.3329406,6.262661,6.348558,6.4305506,6.5164475,6.602344,6.688241,6.278279,5.872221,5.466163,5.056201,4.650143,4.349504,4.0488653,3.7482262,3.4514916,3.1508527,2.9243972,2.7018464,2.475391,2.2489357,2.0263848,2.436347,2.8463092,3.2562714,3.6662338,4.0761957,3.7911747,3.5100577,3.2289407,2.9439192,2.6628022,2.3855898,2.1122816,1.8389735,1.5617609,1.2884527,1.0737107,0.8589685,0.6442264,0.42557985,0.21083772,0.61299115,1.0112402,1.4133936,1.8116426,2.2137961,2.619854,3.0259118,3.435874,3.8419318,4.251894,5.2436123,6.239235,7.2348576,8.23048,9.226103,8.413987,7.601871,6.785851,5.9737353,5.1616197,5.1889505,5.2162814,5.2436123,5.270943,5.298274,6.4032197,7.504261,8.609207,9.710248,10.81129,11.514082,12.216875,12.919667,13.622459,14.325252,12.86891,11.416472,9.96013,8.503788,7.0513506,6.520352,5.989353,5.4583545,4.93126,4.4002614,5.134289,5.8644123,6.5984397,7.328563,8.062591,7.4495993,6.8366084,6.223617,5.610626,5.001539,5.3607445,5.7238536,6.086963,6.4500723,6.813182,6.094772,5.376362,4.661856,3.9434462,3.2250361,3.3265507,3.4241607,3.5256753,3.6232853,3.7247996,3.3616903,2.998581,2.639376,2.2762666,1.9131571,1.9834363,2.0537157,2.1239948,2.194274,2.260649,2.0341935,1.8077383,1.5812829,1.3509232,1.1244678,1.0737107,1.0190489,0.96829176,0.9136301,0.8628729,3.2250361,3.39683,3.5647192,3.736513,3.9044023,4.0761957,3.5842414,3.0883822,2.5964274,2.1044729,1.6125181,1.6515622,1.6906061,1.7335546,1.7725986,1.8116426,1.8311646,1.8506867,1.8741131,1.893635,1.9131571,2.0459068,2.1786566,2.3114061,2.4441557,2.5769055,2.455869,2.338737,2.2216048,2.1044729,1.9873407,1.7218413,1.4524376,1.1869383,0.91753453,0.6481308,0.61299115,0.57394713,0.5388075,0.4997635,0.46071947,0.5231899,0.58566034,0.6481308,0.7106012,0.77307165,0.7106012,0.6481308,0.58566034,0.5231899,0.46071947,0.48805028,0.5114767,0.5388075,0.5622339,0.58566034,0.5583295,0.5309987,0.5036679,0.47633708,0.44900626,0.5427119,0.63641757,0.7262188,0.8199245,0.9136301,1.116659,1.3157835,1.5188124,1.7218413,1.9248703,1.8194515,1.7101282,1.6008049,1.4953861,1.3860629,1.2689307,1.1517987,1.0346665,0.91753453,0.80040246,0.80430686,0.80430686,0.80821127,0.80821127,0.81211567,0.80040246,0.78868926,0.77307165,0.76135844,0.74964523,0.9019169,1.0502841,1.1986516,1.3509232,1.4992905,1.5031948,1.5110037,1.5149081,1.5188124,1.5266213,1.5812829,1.6359446,1.6906061,1.7452679,1.7999294,1.9092526,2.0146716,2.1239948,2.2294137,2.338737,2.3855898,2.436347,2.4871042,2.5378613,2.5886188,2.6042364,2.6159496,2.631567,2.6471848,2.6628022,2.7291772,2.795552,2.8658314,2.9322062,2.998581,3.2289407,3.455396,3.6818514,3.9083066,4.138666,4.068387,3.998108,3.9278288,3.8575494,3.78727,3.619381,3.4475873,3.2757936,3.1079042,2.9361105,3.0220075,3.1079042,3.193801,3.2757936,3.3616903,3.4983444,3.631094,3.767748,3.9044023,4.037152,4.0137253,3.9942036,3.970777,3.9473507,3.9239242,3.8887846,3.853645,3.8185053,3.7833657,3.7482262,3.7443218,3.736513,3.7287042,3.7208953,3.7130866,3.9863946,4.2557983,4.5291066,4.802415,5.0757227,5.02887,4.9781127,4.93126,4.884407,4.8375545,4.7789884,4.716518,4.657952,4.5993857,4.5369153,4.4041657,4.267512,4.1308575,3.998108,3.8614538,3.8224099,3.7833657,3.7443218,3.7013733,3.6623292,3.767748,3.873167,3.978586,4.084005,4.1894236,4.267512,4.3455997,4.4275923,4.50568,4.5876727,4.802415,5.017157,5.2318993,5.446641,5.661383,5.618435,5.579391,5.5364423,5.493494,5.4505453,5.618435,5.7902284,5.958118,6.1299114,6.3017054,6.4032197,6.5086384,6.6140575,6.719476,6.824895,6.805373,6.785851,6.7663293,6.746807,6.7233806,6.754616,6.785851,6.813182,6.844417,6.8756523,7.000593,7.1294384,7.2582836,7.3832245,7.5120697,7.629202,7.7424297,7.8556576,7.9727893,8.086017,9.749292,11.408664,13.068034,14.727406,16.386776,18.003199,19.623526,21.239948,22.85637,24.476698,24.367374,24.25805,24.152632,24.043308,23.937891,21.85294,19.767988,17.683039,15.598087,13.513136,13.45457,13.396004,13.341343,13.282777,13.224211,10.639496,8.054782,5.4700675,2.8853533,0.30063897,0.98000497,1.6593709,2.338737,3.018103,3.7013733,2.959537,2.2216048,1.4797685,0.7418364,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.61689556,1.0463798,1.475864,1.9092526,2.338737,3.06886,3.802888,4.5369153,5.267039,6.001066,5.009348,4.0215344,3.0298162,2.0380979,1.0502841,1.038571,1.0307622,1.0190489,1.0112402,0.999527,0.81211567,0.62470436,0.43729305,0.24988174,0.062470436,0.21083772,0.3631094,0.5114767,0.6637484,0.81211567,0.8511597,0.8941081,0.93315214,0.97219616,1.0112402,1.7023194,2.3933985,3.0805733,3.7716527,4.462732,4.5564375,4.646239,4.7399445,4.83365,4.9234514,5.7316628,6.5398736,7.348085,8.156297,8.960603,8.128965,7.2934237,6.4578815,5.6223392,4.786797,4.0918136,3.39683,2.7018464,2.0068626,1.3118792,1.6632754,2.0107672,2.3621633,2.7135596,3.0610514,3.1859922,3.3070288,3.4280653,3.5530062,3.6740425,3.697469,3.7208953,3.7443218,3.7638438,3.78727,4.415879,5.0483923,5.677001,6.3056097,6.9381227,6.9459314,6.9537406,6.9615493,6.969358,6.9732623,6.5281606,6.086963,5.6418614,5.196759,4.7516575,4.5017757,4.2557983,4.0059166,3.7599394,3.513962,4.041056,4.572055,5.1030536,5.6340523,6.1611466,6.2938967,6.422742,6.551587,6.6843367,6.813182,5.989353,5.1616197,4.337791,3.513962,2.6862288,2.4792955,2.2723622,2.0654287,1.8584955,1.6515622,1.8116426,1.9717231,2.1318035,2.2918842,2.4480603,2.3699722,2.2918842,2.2098918,2.1318035,2.0498111,2.397303,2.7447948,3.0922866,3.4397783,3.78727,3.8965936,4.0020123,4.1113358,4.2167544,4.3260775,4.7009,5.0796275,5.4583545,5.833177,6.211904,5.1616197,4.1113358,3.0610514,2.0107672,0.96438736,1.1283722,1.2962615,1.4641509,1.6320401,1.7999294,1.6164225,1.43682,1.2533131,1.0698062,0.8862993,1.3704453,1.8506867,2.3348327,2.8189783,3.2992198,5.493494,7.6838636,9.878138,12.068507,14.262781,14.012899,13.763018,13.513136,13.263254,13.013372,11.845957,10.67854,9.511124,8.343708,7.1762915,9.483793,11.795199,14.106606,16.414106,18.725513,16.46096,14.200311,11.935758,9.675109,7.4105554,8.015738,8.62092,9.226103,9.8312845,10.436467,10.4286585,10.416945,10.409137,10.397423,10.38571,9.655587,8.921559,8.191436,7.4574084,6.7233806,6.520352,6.3134184,6.1103897,5.903456,5.700427,5.181142,4.661856,4.138666,3.619381,3.1000953,2.5261483,1.9482968,1.3743496,0.80040246,0.22645533,0.41386664,0.60127795,0.78868926,0.97610056,1.1635119,1.4797685,1.796025,2.1161861,2.4324427,2.7486992,3.5451972,4.3416953,5.134289,5.930787,6.7233806,6.532065,6.3407493,6.1494336,5.9542136,5.7628975,5.3997884,5.036679,4.6735697,4.3143644,3.951255,3.474918,2.998581,2.5261483,2.0498111,1.5734742,1.261122,0.94486535,0.62860876,0.31625658,0.0,0.19912452,0.39824903,0.60127795,0.80040246,0.999527,1.3509232,1.698415,2.0498111,2.4012074,2.7486992,6.114294,9.479889,12.845484,16.211079,19.576674,17.152039,14.73131,12.306676,9.885946,7.461313,7.3988423,7.336372,7.2739015,7.211431,7.1489606,6.8756523,6.606249,6.3329406,6.0596323,5.786324,5.743376,5.6965227,5.6535745,5.606722,5.563773,5.3021784,5.040583,4.7828927,4.521298,4.263607,3.873167,3.4866312,3.1000953,2.7135596,2.3231194,2.35045,2.3738766,2.4012074,2.4246337,2.4480603,2.7682211,3.084478,3.4007344,3.7208953,4.037152,3.7013733,3.3655949,3.0337205,2.697942,2.3621633,2.1122816,1.8623998,1.6125181,1.3626363,1.1127546,0.94096094,0.77307165,0.60127795,0.43338865,0.26159495,0.77697605,1.2884527,1.7999294,2.3114061,2.8267872,3.135235,3.4436827,3.7560349,4.0644827,4.376835,5.3334136,6.2938967,7.2543793,8.214863,9.175345,8.52331,7.8751793,7.223144,6.575013,5.9268827,5.758993,5.591104,5.423215,5.2553253,5.087436,6.196286,7.3012323,8.410083,9.518932,10.6238785,11.533605,12.439425,13.349152,14.254972,15.160794,13.673217,12.181735,10.694158,9.202676,7.7111945,6.910792,6.1064854,5.3060827,4.5017757,3.7013733,4.185519,4.6696653,5.153811,5.6418614,6.126007,5.7121406,5.298274,4.8883114,4.474445,4.0605783,4.21285,4.3612175,4.513489,4.661856,4.814128,4.3455997,3.8809757,3.416352,2.951728,2.4871042,2.8267872,3.1625657,3.4983444,3.8380275,4.173806,3.7247996,3.2757936,2.8267872,2.3738766,1.9248703,1.8741131,1.8194515,1.7686942,1.7140326,1.6632754,1.5656652,1.4719596,1.3782539,1.2806439,1.1869383,1.1049459,1.0229534,0.94096094,0.8589685,0.77307165,3.4983444,3.6506162,3.7989833,3.951255,4.0996222,4.251894,3.6857557,3.1235218,2.5612879,1.999054,1.43682,1.5500476,1.6632754,1.7765031,1.8858263,1.999054,2.0615244,2.1239948,2.1864653,2.2489357,2.3114061,2.475391,2.639376,2.7994564,2.9634414,3.1235218,2.9751544,2.8267872,2.6745155,2.5261483,2.3738766,2.0380979,1.698415,1.3626363,1.0268579,0.6871748,0.63641757,0.58566034,0.5388075,0.48805028,0.43729305,0.46071947,0.48805028,0.5114767,0.5388075,0.5622339,0.5231899,0.48805028,0.44900626,0.41386664,0.37482262,0.39824903,0.42557985,0.44900626,0.47633708,0.4997635,0.47633708,0.44900626,0.42557985,0.39824903,0.37482262,0.42557985,0.47633708,0.5231899,0.57394713,0.62470436,0.8745861,1.1244678,1.3743496,1.6242313,1.8741131,1.7608855,1.6515622,1.5383345,1.4251068,1.3118792,1.2376955,1.1635119,1.0893283,1.0112402,0.93705654,0.93705654,0.93705654,0.93705654,0.93705654,0.93705654,0.8394465,0.737932,0.63641757,0.5388075,0.43729305,0.5505207,0.6637484,0.77307165,0.8862993,0.999527,1.0268579,1.0502841,1.0737107,1.1010414,1.1244678,1.1986516,1.2767396,1.3509232,1.4251068,1.4992905,1.5266213,1.5500476,1.5734742,1.6008049,1.6242313,1.6867018,1.7491722,1.8116426,1.8741131,1.9365835,1.9756275,2.0107672,2.0498111,2.0888553,2.1239948,2.1864653,2.2489357,2.3114061,2.3738766,2.436347,2.736986,3.0376248,3.338264,3.638903,3.9356375,3.912211,3.8887846,3.8614538,3.8380275,3.8106966,3.6232853,3.435874,3.2484627,3.0610514,2.87364,2.998581,3.1235218,3.2484627,3.3734035,3.4983444,3.5764325,3.6506162,3.7247996,3.7989833,3.873167,3.8497405,3.8263142,3.7989833,3.775557,3.7482262,3.7247996,3.7013733,3.6740425,3.6506162,3.6232853,3.6740425,3.7247996,3.775557,3.8263142,3.873167,4.173806,4.474445,4.775084,5.0757227,5.376362,5.3138914,5.251421,5.1889505,5.12648,5.0640097,4.9624953,4.860981,4.7633705,4.661856,4.564246,4.4119744,4.263607,4.1113358,3.9629683,3.8106966,3.7013733,3.5881457,3.474918,3.3616903,3.2484627,3.349977,3.4514916,3.5491016,3.6506162,3.7482262,3.8497405,3.951255,4.0488653,4.1503797,4.251894,4.4861584,4.7243266,4.9624953,5.2006636,5.4388323,5.3997884,5.3607445,5.3256044,5.2865605,5.251421,5.4388323,5.6262436,5.813655,6.001066,6.1884775,6.3251314,6.461786,6.5984397,6.7389984,6.8756523,6.8639393,6.8483214,6.8366084,6.824895,6.813182,6.8756523,6.9381227,7.000593,7.0630636,7.125534,7.3129454,7.5003567,7.687768,7.8751793,8.062591,8.011833,7.9610763,7.914223,7.8634663,7.812709,9.776623,11.736633,13.700547,15.664462,17.624472,19.326792,21.025206,22.723621,24.425941,26.124355,25.726107,25.323954,24.925705,24.52355,24.125301,22.262901,20.400501,18.538101,16.675701,14.813302,14.274494,13.735687,13.200784,12.661977,12.123169,9.698535,7.2739015,4.8492675,2.4246337,0.0,0.92534333,1.8506867,2.77603,3.7013733,4.6267166,3.7013733,2.77603,1.8506867,0.92534333,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.63641757,1.0893283,1.5383345,1.9873407,2.436347,3.1508527,3.8614538,4.575959,5.2865605,6.001066,4.911738,3.8263142,2.736986,1.6515622,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.8628729,1.7257458,2.5886188,3.4514916,4.3143644,4.388548,4.462732,4.5369153,4.6110992,4.689187,5.8761253,7.0630636,8.250002,9.43694,10.6238785,9.487698,8.351517,7.211431,6.0752497,4.939069,4.138666,3.338264,2.5378613,1.737459,0.93705654,1.4251068,1.9131571,2.4012074,2.8892577,3.3734035,3.4632049,3.5491016,3.638903,3.7247996,3.8106966,3.8106966,3.8106966,3.8106966,3.8106966,3.8106966,4.650143,5.4856853,6.3251314,7.1606736,8.00012,7.9259367,7.8517528,7.773665,7.699481,7.6252975,7.012306,6.3993154,5.786324,5.173333,4.564246,4.251894,3.9356375,3.6232853,3.310933,2.998581,3.6623292,4.3260775,4.985922,5.64967,6.3134184,6.4383593,6.5633,6.688241,6.813182,6.9381227,6.0518236,5.1616197,4.2753205,3.3890212,2.4988174,2.3231194,2.1513257,1.9756275,1.7999294,1.6242313,1.8233559,2.0263848,2.2255092,2.4246337,2.6237583,2.436347,2.2489357,2.0615244,1.8741131,1.6867018,1.999054,2.3114061,2.6237583,2.9361105,3.2484627,3.310933,3.3734035,3.435874,3.4983444,3.5608149,3.951255,4.337791,4.7243266,5.1108627,5.5013027,4.5993857,3.7013733,2.7994564,1.901444,0.999527,1.2494087,1.4992905,1.7491722,1.999054,2.2489357,1.7999294,1.3509232,0.9019169,0.44900626,0.0,0.13665408,0.27330816,0.41386664,0.5505207,0.6871748,2.787743,4.8883114,6.98888,9.089449,11.186112,10.77615,10.362284,9.948417,9.538455,9.124588,8.749765,8.374943,8.00012,7.6252975,7.250475,8.738052,10.22563,11.713207,13.200784,14.688361,13.411622,12.138786,10.862047,9.589212,8.312472,8.238289,8.164105,8.086017,8.011833,7.9376497,8.148487,8.36323,8.574067,8.78881,8.999647,8.476458,7.9493628,7.426173,6.899079,6.375889,5.989353,5.5989127,5.212377,4.825841,4.4393053,4.173806,3.912211,3.6506162,3.3890212,3.1235218,2.5495746,1.9756275,1.4016805,0.8238289,0.24988174,0.48805028,0.7262188,0.96438736,1.1986516,1.43682,1.8389735,2.2372224,2.639376,3.0376248,3.435874,4.3260775,5.212377,6.098676,6.98888,7.8751793,7.726812,7.57454,7.426173,7.2739015,7.125534,6.688241,6.250948,5.813655,5.376362,4.939069,4.298747,3.6623292,3.0259118,2.3855898,1.7491722,1.4016805,1.0502841,0.698888,0.3513962,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.9019169,1.4875772,2.0732377,2.6628022,3.2484627,7.1762915,11.100216,15.024139,18.95197,22.875893,19.900738,16.925583,13.950429,10.975275,8.00012,7.9376497,7.8751793,7.812709,7.7502384,7.687768,7.211431,6.7389984,6.262661,5.786324,5.3138914,5.138193,4.9624953,4.786797,4.6110992,4.4393053,4.3260775,4.21285,4.0996222,3.9863946,3.873167,3.4007344,2.9243972,2.4480603,1.9756275,1.4992905,1.7765031,2.0498111,2.3231194,2.6003318,2.87364,3.1000953,3.3265507,3.5491016,3.775557,3.998108,3.611572,3.2250361,2.8385005,2.4519646,2.0615244,1.8389735,1.6125181,1.3860629,1.1635119,0.93705654,0.81211567,0.6871748,0.5622339,0.43729305,0.31235218,0.93705654,1.5617609,2.1864653,2.8111696,3.435874,3.6506162,3.8614538,4.0761957,4.2870336,4.5017757,5.423215,6.348558,7.2739015,8.1992445,9.124588,8.636538,8.148487,7.6643414,7.1762915,6.688241,6.3251314,5.9620223,5.5989127,5.2358036,4.8765984,5.989353,7.098203,8.210958,9.323712,10.436467,11.549222,12.661977,13.774731,14.8874855,16.00024,14.473619,12.950902,11.424281,9.901564,8.374943,7.3012323,6.223617,5.1499066,4.0761957,2.998581,3.2367494,3.474918,3.7130866,3.951255,4.1894236,3.9746814,3.7638438,3.5491016,3.338264,3.1235218,3.0610514,2.998581,2.9361105,2.87364,2.8111696,2.6003318,2.3855898,2.174752,1.9639144,1.7491722,2.3231194,2.900971,3.474918,4.0488653,4.6267166,4.087909,3.5491016,3.0141985,2.475391,1.9365835,1.7608855,1.5890918,1.4133936,1.2376955,1.0619974,1.1010414,1.1361811,1.175225,1.2142692,1.2494087,1.1361811,1.0268579,0.9136301,0.80040246,0.6871748,2.8892577,3.049338,3.2094188,3.3655949,3.5256753,3.6857557,3.3538816,3.0220075,2.690133,2.358259,2.0263848,2.1318035,2.233318,2.338737,2.4441557,2.5495746,2.5651922,2.5808098,2.5964274,2.6081407,2.6237583,2.6823244,2.7408905,2.795552,2.854118,2.912684,2.7604125,2.6081407,2.455869,2.3035975,2.1513257,1.8663043,1.5851873,1.3040704,1.0190489,0.737932,0.6832704,0.63251317,0.58175594,0.5270943,0.47633708,0.4958591,0.5192855,0.5427119,0.5661383,0.58566034,0.57394713,0.5583295,0.5427119,0.5270943,0.5114767,0.5036679,0.49195468,0.48414588,0.47243267,0.46071947,0.5036679,0.5427119,0.58175594,0.62079996,0.6637484,0.6442264,0.62079996,0.60127795,0.58175594,0.5622339,0.76526284,0.96829176,1.1713207,1.3743496,1.5734742,1.4875772,1.4016805,1.3118792,1.2259823,1.1361811,1.0619974,0.9878138,0.9136301,0.8394465,0.76135844,0.76526284,0.76916724,0.76916724,0.77307165,0.77307165,0.6910792,0.60908675,0.5270943,0.44510186,0.3631094,0.45291066,0.5427119,0.63251317,0.7223144,0.81211567,0.8316377,0.8511597,0.8706817,0.8941081,0.9136301,0.97610056,1.0424755,1.1088502,1.1713207,1.2376955,1.2650263,1.2923572,1.319688,1.3470187,1.3743496,1.4329157,1.4914817,1.5461433,1.6047094,1.6632754,1.7023194,1.7413634,1.7843118,1.8233559,1.8623998,1.9365835,2.0068626,2.0810463,2.1513257,2.2255092,2.5183394,2.8111696,3.1039999,3.39683,3.6857557,3.6506162,3.611572,3.5764325,3.5373883,3.4983444,3.39683,3.2953155,3.193801,3.0883822,2.9868677,3.1039999,3.2172275,3.3343596,3.4475873,3.5608149,3.5647192,3.5686235,3.5686235,3.5725281,3.5764325,3.638903,3.7052777,3.7716527,3.8341231,3.900498,3.9317331,3.9668727,3.998108,4.029343,4.0605783,4.0996222,4.138666,4.173806,4.21285,4.251894,4.548629,4.845363,5.142098,5.4388323,5.735567,5.7980375,5.8566036,5.919074,5.9776397,6.036206,5.852699,5.6691923,5.481781,5.298274,5.1108627,4.9937305,4.8765984,4.759466,4.6423345,4.5252023,4.4314966,4.3338866,4.240181,4.1464753,4.0488653,4.095718,4.1464753,4.193328,4.240181,4.2870336,4.337791,4.388548,4.4393053,4.4861584,4.5369153,4.7009,4.860981,5.024966,5.1889505,5.349031,5.3724575,5.395884,5.4193106,5.4388323,5.462259,5.610626,5.758993,5.903456,6.0518236,6.2001905,6.36808,6.5359693,6.703859,6.871748,7.0357327,7.039637,7.043542,7.043542,7.0474463,7.0513506,7.043542,7.0357327,7.027924,7.0201154,7.012306,7.3129454,7.6135845,7.914223,8.210958,8.511597,8.6131115,8.718531,8.8200445,8.921559,9.023073,10.9089,12.794726,14.6805525,16.56638,18.448301,20.521538,22.590872,24.660204,26.729538,28.79887,27.807154,26.815435,25.823717,24.828094,23.836376,21.688955,19.541533,17.394112,15.246691,13.09927,12.419904,11.740538,11.061172,10.381805,9.698535,7.7619514,5.8214636,3.8809757,1.9404879,0.0,0.76916724,1.53443,2.3035975,3.06886,3.8380275,3.06886,2.3035975,1.53443,0.76916724,0.0,0.0,0.0,0.0,0.0,0.0,0.10932326,0.21474212,0.3240654,0.42948425,0.5388075,0.9136301,1.2923572,1.6710842,2.0459068,2.4246337,2.9048753,3.3851168,3.8653584,4.3455997,4.825841,4.0332475,3.2445583,2.455869,1.6632754,0.8745861,0.698888,0.5231899,0.3513962,0.1756981,0.0,0.3357786,0.6754616,1.0112402,1.3509232,1.6867018,1.53443,1.3782539,1.2220778,1.0659018,0.9136301,0.8784905,0.8472553,0.8160201,0.78088045,0.74964523,1.4094892,2.069333,2.7291772,3.3890212,4.0488653,4.3416953,4.6345253,4.927356,5.2201858,5.5130157,6.5398736,7.5667315,8.59359,9.6243515,10.651209,9.753197,8.855185,7.957172,7.0591593,6.1611466,5.3256044,4.4861584,3.6506162,2.8111696,1.9756275,2.3075018,2.639376,2.97125,3.3031244,3.638903,3.7013733,3.7638438,3.8263142,3.8887846,3.951255,3.9044023,3.853645,3.8067923,3.7599394,3.7130866,4.3416953,4.9663997,5.5950084,6.223617,6.8483214,6.8561306,6.8639393,6.871748,6.8795567,6.8873653,6.2548523,5.6223392,4.989826,4.357313,3.7247996,3.5256753,3.330455,3.1313305,2.9361105,2.736986,3.2914112,3.8458362,4.4041657,4.958591,5.5130157,5.606722,5.704332,5.7980375,5.891743,5.989353,5.2865605,4.5837684,3.8809757,3.1781836,2.475391,2.338737,2.1981785,2.0615244,1.9248703,1.7882162,1.8897307,1.9912452,2.096664,2.1981785,2.2996929,2.1161861,1.9287747,1.7452679,1.5617609,1.3743496,1.6242313,1.8741131,2.1239948,2.3738766,2.6237583,2.717464,2.8111696,2.900971,2.9946766,3.0883822,3.4241607,3.7638438,4.0996222,4.4393053,4.775084,4.0801005,3.3851168,2.690133,1.9951496,1.3001659,1.4797685,1.6593709,1.8389735,2.018576,2.1981785,1.7608855,1.319688,0.8784905,0.44119745,0.0,0.74574083,1.4914817,2.233318,2.979059,3.7247996,4.825841,5.9268827,7.0240197,8.125061,9.226103,10.186585,11.143164,12.103647,13.06413,14.024612,12.697116,11.369619,10.042123,8.714626,7.387129,8.784905,10.182681,11.580457,12.978233,14.376009,13.224211,12.076316,10.924518,9.776623,8.624825,8.410083,8.19534,7.9805984,7.7658563,7.551114,7.621393,7.6955767,7.7658563,7.8400397,7.914223,7.648724,7.3832245,7.1177254,6.852226,6.5867267,6.196286,5.805846,5.4193106,5.02887,4.6384296,4.376835,4.1113358,3.8497405,3.5881457,3.3265507,2.8814487,2.436347,1.9912452,1.5461433,1.1010414,1.3118792,1.5266213,1.737459,1.9482968,2.1630387,2.5964274,3.0259118,3.4593005,3.892689,4.3260775,4.970304,5.6145306,6.2587566,6.9068875,7.551114,7.4691215,7.3910336,7.309041,7.230953,7.1489606,6.578918,6.008875,5.4388323,4.8687897,4.298747,3.7443218,3.1898966,2.6354716,2.0810463,1.5266213,1.2181735,0.9136301,0.60908675,0.30454338,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.94876975,1.6437533,2.3426414,3.0415294,3.736513,6.75852,9.780528,12.806439,15.828446,18.850454,16.48829,14.126127,11.763964,9.4018,7.0357327,6.883461,6.727285,6.571109,6.4188375,6.262661,5.8761253,5.4856853,5.099149,4.7126136,4.3260775,4.279225,4.2284675,4.181615,4.134762,4.087909,3.9824903,3.8770714,3.7716527,3.6662338,3.5608149,3.1430438,2.7291772,2.3114061,1.893635,1.475864,1.6906061,1.9053483,2.1200905,2.3348327,2.5495746,2.77603,3.0063896,3.232845,3.4593005,3.6857557,3.3343596,2.979059,2.6237583,2.2684577,1.9131571,1.698415,1.4875772,1.2767396,1.0619974,0.8511597,0.7301232,0.60908675,0.48805028,0.3709182,0.24988174,0.9058213,1.5617609,2.2137961,2.8697357,3.5256753,3.6271896,3.7287042,3.8341231,3.9356375,4.037152,4.958591,5.8761253,6.7975645,7.719003,8.636538,8.210958,7.7814736,7.355894,6.9264097,6.5008297,6.278279,6.0596323,5.840986,5.618435,5.3997884,6.2938967,7.1841,8.078208,8.968412,9.86252,10.862047,11.861574,12.861101,13.860628,14.864059,13.431144,12.002132,10.573121,9.14411,7.7111945,6.6687193,5.6262436,4.5837684,3.541293,2.4988174,2.7447948,2.9907722,3.2367494,3.4788225,3.7247996,3.4905357,3.2562714,3.018103,2.7838387,2.5495746,2.4988174,2.4441557,2.3933985,2.338737,2.2879796,2.1122816,1.9365835,1.7608855,1.5890918,1.4133936,1.9443923,2.4714866,3.0024853,3.533484,4.0605783,3.6506162,3.2367494,2.8267872,2.4129205,1.999054,1.9092526,1.8194515,1.7296503,1.639849,1.5500476,1.5461433,1.5461433,1.542239,1.5383345,1.5383345,1.4212024,1.3040704,1.1869383,1.0659018,0.94876975,2.2762666,2.4441557,2.6159496,2.7838387,2.9556324,3.1235218,3.0220075,2.920493,2.8189783,2.7135596,2.612045,2.7096553,2.8072653,2.9048753,3.0024853,3.1000953,3.06886,3.0337205,3.0024853,2.97125,2.9361105,2.8892577,2.8424048,2.795552,2.7486992,2.7018464,2.5456703,2.3894942,2.233318,2.0810463,1.9248703,1.698415,1.4680552,1.2415999,1.0151446,0.78868926,0.7340276,0.679366,0.62079996,0.5661383,0.5114767,0.5309987,0.5544251,0.57394713,0.59346914,0.61299115,0.62079996,0.62860876,0.63641757,0.6442264,0.6481308,0.60518235,0.5583295,0.5153811,0.46852827,0.42557985,0.5309987,0.63641757,0.7418364,0.8433509,0.94876975,0.8589685,0.76916724,0.679366,0.58956474,0.4997635,0.6559396,0.80821127,0.96438736,1.1205635,1.2767396,1.2142692,1.1517987,1.0893283,1.0268579,0.96438736,0.8862993,0.81211567,0.737932,0.6637484,0.58566034,0.59346914,0.59737355,0.60127795,0.60908675,0.61299115,0.5466163,0.48414588,0.41777104,0.3513962,0.28892577,0.3553006,0.42167544,0.48805028,0.5583295,0.62470436,0.64032197,0.6559396,0.6715572,0.6832704,0.698888,0.75354964,0.80821127,0.8667773,0.92143893,0.97610056,1.0034313,1.0346665,1.0659018,1.0932326,1.1244678,1.1791295,1.2298868,1.2806439,1.3353056,1.3860629,1.4290112,1.4719596,1.5149081,1.5578566,1.6008049,1.6827974,1.7647898,1.8467822,1.9287747,2.0107672,2.2957885,2.5808098,2.8658314,3.1508527,3.435874,3.3890212,3.338264,3.2875066,3.2367494,3.1859922,3.1703746,3.1508527,3.135235,3.1157131,3.1000953,3.2055142,3.310933,3.416352,3.521771,3.6232853,3.5569105,3.4866312,3.416352,3.3460727,3.2757936,3.4280653,3.5842414,3.7404175,3.8965936,4.0488653,4.138666,4.2284675,4.318269,4.40807,4.5017757,4.5252023,4.548629,4.575959,4.5993857,4.6267166,4.919547,5.2162814,5.5091114,5.805846,6.098676,6.282183,6.46569,6.649197,6.8287997,7.012306,6.7429028,6.473499,6.2040954,5.930787,5.661383,5.579391,5.493494,5.407597,5.3217,5.2358036,5.1616197,5.083532,5.0054436,4.927356,4.8492675,4.845363,4.841459,4.83365,4.829746,4.825841,4.825841,4.825841,4.825841,4.825841,4.825841,4.911738,5.001539,5.087436,5.173333,5.263134,5.3451266,5.4271193,5.5091114,5.591104,5.6730967,5.7824197,5.891743,5.997162,6.1064854,6.211904,6.4110284,6.606249,6.805373,7.000593,7.1997175,7.2192397,7.2348576,7.2543793,7.269997,7.2856145,7.211431,7.1333427,7.055255,6.9771667,6.899079,7.3129454,7.726812,8.136774,8.550641,8.960603,9.218294,9.47208,9.725866,9.983557,10.237343,12.045081,13.852819,15.660558,17.468296,19.276033,21.716286,24.156536,26.596788,29.033134,31.473387,29.888199,28.306917,26.72173,25.136541,23.551353,21.118912,18.68647,16.254026,13.821584,11.389141,10.565312,9.741484,8.921559,8.097731,7.2739015,5.8214636,4.365122,2.9087796,1.456342,0.0,0.60908675,1.2181735,1.8311646,2.4402514,3.049338,2.4402514,1.8311646,1.2181735,0.60908675,0.0,0.0,0.0,0.0,0.0,0.0,0.1756981,0.3553006,0.5309987,0.7106012,0.8862993,1.1908426,1.4992905,1.8038338,2.1083772,2.4129205,2.6588979,2.9087796,3.154757,3.4007344,3.6506162,3.1586614,2.6667068,2.1708477,1.678893,1.1869383,0.94876975,0.7106012,0.47633708,0.23816854,0.0,0.6754616,1.3509232,2.0263848,2.7018464,3.3734035,3.0649557,2.7565079,2.4441557,2.135708,1.8233559,1.7608855,1.6945106,1.6281357,1.5656652,1.4992905,1.9561055,2.416825,2.87364,3.330455,3.78727,4.298747,4.806319,5.3177958,5.8292727,6.336845,7.2036223,8.074304,8.941081,9.807858,10.674636,10.018696,9.358852,8.702912,8.043069,7.387129,6.5125427,5.6379566,4.7633705,3.8887846,3.0141985,3.1898966,3.3655949,3.5451972,3.7208953,3.900498,3.9356375,3.9746814,4.0137253,4.0488653,4.087909,3.9942036,3.8965936,3.802888,3.7091823,3.611572,4.029343,4.447114,4.8648853,5.282656,5.700427,5.7902284,5.8800297,5.969831,6.0596323,6.1494336,5.4973984,4.845363,4.193328,3.541293,2.8892577,2.803361,2.7213683,2.639376,2.5573835,2.475391,2.9243972,3.3694992,3.8185053,4.263607,4.7126136,4.7789884,4.841459,4.9078336,4.9742084,5.036679,4.521298,4.0020123,3.4866312,2.9673457,2.4480603,2.35045,2.2489357,2.1513257,2.0498111,1.9482968,1.9561055,1.9600099,1.9639144,1.9717231,1.9756275,1.7921207,1.6086137,1.4290112,1.2455044,1.0619974,1.2494087,1.43682,1.6242313,1.8116426,1.999054,2.1239948,2.2450314,2.366068,2.4910088,2.612045,2.900971,3.1859922,3.474918,3.7638438,4.0488653,3.5608149,3.06886,2.5808098,2.0888553,1.6008049,1.7101282,1.8194515,1.9287747,2.0380979,2.1513257,1.7218413,1.2884527,0.8589685,0.42948425,0.0,1.3509232,2.7057507,4.056674,5.4115014,6.7624245,6.8639393,6.9615493,7.0630636,7.1606736,7.262188,9.597021,11.927949,14.258877,16.59371,18.924637,16.644466,14.364296,12.084125,9.803954,7.523783,8.831758,10.139732,11.447707,12.755682,14.063657,13.036799,12.013845,10.986988,9.964035,8.937177,8.581876,8.226576,7.871275,7.5159745,7.1606736,7.094299,7.027924,6.9615493,6.89127,6.824895,6.8209906,6.813182,6.8092775,6.805373,6.801469,6.407124,6.016684,5.6223392,5.2318993,4.8375545,4.575959,4.3143644,4.0488653,3.78727,3.5256753,3.2094188,2.893162,2.5808098,2.2645533,1.9482968,2.135708,2.3231194,2.514435,2.7018464,2.8892577,3.3538816,3.8185053,4.283129,4.747753,5.212377,5.6145306,6.016684,6.4188375,6.8209906,7.223144,7.2153354,7.2036223,7.195813,7.1841,7.1762915,6.473499,5.7707067,5.067914,4.365122,3.6623292,3.1898966,2.717464,2.2450314,1.7725986,1.3001659,1.038571,0.78088045,0.5192855,0.26159495,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.9956226,1.8038338,2.6081407,3.416352,4.224563,6.3446536,8.464745,10.584834,12.704925,14.825015,13.075843,11.326671,9.573594,7.824422,6.0752497,5.8292727,5.579391,5.3334136,5.083532,4.8375545,4.5369153,4.2362766,3.9356375,3.638903,3.338264,3.416352,3.4983444,3.5764325,3.6584249,3.736513,3.638903,3.541293,3.4436827,3.3460727,3.2484627,2.8892577,2.5300527,2.1708477,1.8116426,1.4485333,1.6047094,1.7608855,1.9131571,2.069333,2.2255092,2.455869,2.6862288,2.9165885,3.1430438,3.3734035,3.0532427,2.7291772,2.4090161,2.084951,1.7608855,1.5617609,1.3626363,1.1635119,0.96438736,0.76135844,0.6481308,0.5309987,0.41777104,0.30063897,0.18741131,0.8706817,1.5578566,2.241127,2.9283018,3.611572,3.6037633,3.5959544,3.5881457,3.5842414,3.5764325,4.4900627,5.4036927,6.321227,7.2348576,8.148487,7.7814736,7.4144597,7.0474463,6.6804323,6.3134184,6.2353306,6.1572423,6.0791545,6.001066,5.9268827,6.5984397,7.269997,7.941554,8.6131115,9.288573,10.174872,11.061172,11.951375,12.837675,13.723974,12.388668,11.053363,9.718058,8.386656,7.0513506,6.04011,5.02887,4.0215344,3.0102942,1.999054,2.25284,2.5066261,2.7565079,3.0102942,3.2640803,3.0063896,2.7486992,2.4910088,2.233318,1.9756275,1.9326792,1.8897307,1.8467822,1.8038338,1.7608855,1.6242313,1.4875772,1.3509232,1.2142692,1.0737107,1.5617609,2.0459068,2.5300527,3.0141985,3.4983444,3.213323,2.9243972,2.639376,2.35045,2.0615244,2.05762,2.0537157,2.0459068,2.0420024,2.0380979,1.9951496,1.9522011,1.9092526,1.8663043,1.8233559,1.7023194,1.5812829,1.456342,1.3353056,1.2142692,1.6632754,1.8428779,2.0224805,2.2020829,2.3816853,2.5612879,2.690133,2.8189783,2.9439192,3.0727646,3.2016098,3.2914112,3.3812122,3.4710135,3.5608149,3.6506162,3.5686235,3.4905357,3.408543,3.330455,3.2484627,3.096191,2.9439192,2.7916477,2.639376,2.4871042,2.330928,2.1708477,2.0146716,1.8584955,1.698415,1.5266213,1.3548276,1.183034,1.0112402,0.8394465,0.78088045,0.7223144,0.6637484,0.60908675,0.5505207,0.5661383,0.58566034,0.60127795,0.62079996,0.63641757,0.6676528,0.698888,0.7262188,0.75745404,0.78868926,0.7066968,0.62860876,0.5466163,0.46852827,0.38653582,0.5583295,0.7262188,0.8980125,1.0659018,1.2376955,1.077615,0.91753453,0.75745404,0.59737355,0.43729305,0.5466163,0.6520352,0.76135844,0.8667773,0.97610056,0.93705654,0.9019169,0.8628729,0.8238289,0.78868926,0.7106012,0.63641757,0.5622339,0.48805028,0.41386664,0.42167544,0.42557985,0.43338865,0.44119745,0.44900626,0.40215343,0.3553006,0.30844778,0.26159495,0.21083772,0.25769055,0.30063897,0.3474918,0.39434463,0.43729305,0.44900626,0.45681506,0.46852827,0.47633708,0.48805028,0.5309987,0.57785153,0.62079996,0.6676528,0.7106012,0.74574083,0.77697605,0.80821127,0.8433509,0.8745861,0.92143893,0.96829176,1.0190489,1.0659018,1.1127546,1.1557031,1.2025559,1.2494087,1.2923572,1.33921,1.4290112,1.5227169,1.6164225,1.7062237,1.7999294,2.077142,2.3543546,2.631567,2.9087796,3.1859922,3.1235218,3.0610514,2.998581,2.9361105,2.87364,2.9439192,3.0102942,3.076669,3.1469483,3.213323,3.3070288,3.4007344,3.4983444,3.59205,3.6857557,3.5451972,3.4007344,3.260176,3.1157131,2.9751544,3.2211318,3.4632049,3.7091823,3.9551594,4.2011366,4.3455997,4.493967,4.6423345,4.7907014,4.939069,4.950782,4.9624953,4.9742084,4.985922,5.001539,5.2943697,5.5832953,5.8761253,6.168956,6.461786,6.7663293,7.0708723,7.37932,7.6838636,7.988407,7.633106,7.277806,6.9225054,6.5672045,6.211904,6.1611466,6.1064854,6.055728,6.001066,5.950309,5.891743,5.8292727,5.7707067,5.708236,5.64967,5.591104,5.5364423,5.477876,5.4193106,5.3607445,5.3138914,5.263134,5.212377,5.1616197,5.1108627,5.12648,5.138193,5.1499066,5.1616197,5.173333,5.3177958,5.4583545,5.602817,5.743376,5.8878384,5.9542136,6.0205884,6.0908675,6.1572423,6.223617,6.453977,6.6804323,6.9068875,7.1333427,7.363703,7.394938,7.426173,7.461313,7.492548,7.523783,7.37932,7.230953,7.082586,6.9342184,6.785851,7.3129454,7.8361354,8.36323,8.886419,9.413514,9.8195715,10.22563,10.6355915,11.04165,11.4516115,13.181262,14.9109125,16.640562,18.370213,20.099863,22.911032,25.718298,28.529467,31.340637,34.151806,31.97315,29.794493,27.615837,25.441086,23.262428,20.544964,17.827501,15.110037,12.392572,9.675109,8.710721,7.746334,6.7780423,5.813655,4.8492675,3.8809757,2.9087796,1.9404879,0.96829176,0.0,0.45291066,0.9058213,1.358732,1.8116426,2.260649,1.8116426,1.358732,0.9058213,0.45291066,0.0,0.0,0.0,0.0,0.0,0.0,0.24597734,0.4958591,0.7418364,0.9917182,1.2376955,1.4680552,1.7023194,1.9365835,2.1669433,2.4012074,2.416825,2.4285383,2.4441557,2.4597735,2.475391,2.280171,2.084951,1.8897307,1.6945106,1.4992905,1.1986516,0.9019169,0.60127795,0.30063897,0.0,1.0112402,2.0263848,3.0376248,4.0488653,5.0640097,4.5993857,4.1308575,3.6662338,3.2016098,2.736986,2.639376,2.541766,2.4441557,2.3465457,2.2489357,2.5066261,2.7604125,3.0141985,3.2718892,3.5256753,4.251894,4.9781127,5.708236,6.434455,7.1606736,7.871275,8.577971,9.284669,9.991365,10.698062,10.284196,9.866425,9.448653,9.030883,8.6131115,7.699481,6.785851,5.8761253,4.9624953,4.0488653,4.0722914,4.095718,4.1191444,4.138666,4.1620927,4.173806,4.1894236,4.2011366,4.21285,4.224563,4.084005,3.9395418,3.7989833,3.6545205,3.513962,3.7208953,3.9278288,4.134762,4.3416953,4.548629,4.7243266,4.8961205,5.067914,5.239708,5.4115014,4.7399445,4.068387,3.39683,2.7213683,2.0498111,2.0810463,2.1161861,2.1474214,2.1786566,2.2137961,2.5534792,2.893162,3.232845,3.5725281,3.912211,3.9473507,3.9824903,4.01763,4.0527697,4.087909,3.7560349,3.4241607,3.0883822,2.7565079,2.4246337,2.3621633,2.2996929,2.2372224,2.174752,2.1122816,2.018576,1.9287747,1.8350691,1.7413634,1.6515622,1.4680552,1.2884527,1.1088502,0.92924774,0.74964523,0.8745861,0.999527,1.1244678,1.2494087,1.3743496,1.5266213,1.678893,1.8311646,1.9834363,2.135708,2.3738766,2.612045,2.8502135,3.0883822,3.3265507,3.0415294,2.7565079,2.4714866,2.1864653,1.901444,1.9404879,1.979532,2.018576,2.0615244,2.1005683,1.678893,1.261122,0.8394465,0.42167544,0.0,1.9600099,3.9200199,5.8800297,7.8400397,9.80005,8.898132,8.00012,7.098203,6.2001905,5.298274,9.0035515,12.708829,16.414106,20.119385,23.824663,20.591818,17.358973,14.126127,10.893282,7.6643414,8.878611,10.096785,11.314958,12.533132,13.751305,12.849388,11.951375,11.0494585,10.151445,9.249529,8.75367,8.261715,7.7658563,7.269997,6.774138,6.5672045,6.3602715,6.153338,5.9464045,5.735567,5.9932575,6.2470436,6.5008297,6.75852,7.012306,6.617962,6.223617,5.8292727,5.4310236,5.036679,4.775084,4.513489,4.251894,3.9863946,3.7247996,3.541293,3.3538816,3.1703746,2.9868677,2.7994564,2.9634414,3.1235218,3.2875066,3.4514916,3.611572,4.1113358,4.607195,5.1069584,5.602817,6.098676,6.2587566,6.4188375,6.578918,6.7389984,6.899079,6.9615493,7.0201154,7.0786815,7.141152,7.1997175,6.364176,5.5286336,4.6930914,3.8614538,3.0259118,2.6354716,2.2450314,1.8545911,1.4641509,1.0737107,0.8589685,0.6442264,0.42948425,0.21474212,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,1.0424755,1.9600099,2.8775444,3.795079,4.7126136,5.930787,7.1489606,8.36323,9.581403,10.799577,9.663396,8.52331,7.387129,6.250948,5.1108627,4.7711797,4.4314966,4.0918136,3.7521305,3.4124475,3.2016098,2.9868677,2.77603,2.5612879,2.35045,2.5573835,2.7643168,2.97125,3.1781836,3.3890212,3.2992198,3.2094188,3.1157131,3.0259118,2.9361105,2.6354716,2.330928,2.0302892,1.7257458,1.4251068,1.5188124,1.6164225,1.7101282,1.8038338,1.901444,2.1318035,2.366068,2.5964274,2.8306916,3.0610514,2.7721257,2.4831998,2.194274,1.901444,1.6125181,1.4251068,1.2376955,1.0502841,0.8628729,0.6754616,0.5661383,0.45681506,0.3435874,0.23426414,0.12494087,0.8394465,1.5539521,2.2684577,2.9868677,3.7013733,3.5842414,3.4632049,3.3460727,3.2289407,3.1118085,4.0215344,4.93126,5.840986,6.7507114,7.6643414,7.355894,7.0474463,6.7389984,6.434455,6.126007,6.1884775,6.2548523,6.321227,6.3836975,6.4500723,6.902983,7.355894,7.8088045,8.261715,8.710721,9.487698,10.260769,11.037745,11.810817,12.587793,11.346193,10.108498,8.866898,7.629202,6.387602,5.4115014,4.4314966,3.455396,2.4792955,1.4992905,1.7608855,2.018576,2.280171,2.541766,2.7994564,2.5183394,2.241127,1.9600099,1.678893,1.4016805,1.3665408,1.3353056,1.3040704,1.2689307,1.2376955,1.1361811,1.038571,0.93705654,0.8394465,0.737932,1.1791295,1.6164225,2.05762,2.4988174,2.9361105,2.77603,2.612045,2.4480603,2.2879796,2.1239948,2.2059872,2.2840753,2.366068,2.4441557,2.5261483,2.4441557,2.358259,2.2762666,2.194274,2.1122816,1.9834363,1.8584955,1.7296503,1.6008049,1.475864,1.0502841,1.2415999,1.4290112,1.620327,1.8116426,1.999054,2.358259,2.7135596,3.0727646,3.4280653,3.78727,3.8692627,3.951255,4.0332475,4.1191444,4.2011366,4.0722914,3.9434462,3.8185053,3.68966,3.5608149,3.3031244,3.049338,2.7916477,2.533957,2.2762666,2.1161861,1.9561055,1.796025,1.6359446,1.475864,1.358732,1.2415999,1.1205635,1.0034313,0.8862993,0.8277333,0.76916724,0.7066968,0.6481308,0.58566034,0.60127795,0.61689556,0.63251317,0.6481308,0.6637484,0.7145056,0.76916724,0.8199245,0.8706817,0.92534333,0.80821127,0.6949836,0.58175594,0.46462387,0.3513962,0.58566034,0.8199245,1.0541886,1.2884527,1.5266213,1.2962615,1.0659018,0.8355421,0.60518235,0.37482262,0.43338865,0.4958591,0.5544251,0.61689556,0.6754616,0.6637484,0.6481308,0.63641757,0.62470436,0.61299115,0.5388075,0.46071947,0.38653582,0.31235218,0.23816854,0.24597734,0.25769055,0.26940376,0.27721256,0.28892577,0.25769055,0.22645533,0.19912452,0.1678893,0.13665408,0.16008049,0.1835069,0.20693332,0.22645533,0.24988174,0.25378615,0.26159495,0.26549935,0.26940376,0.27330816,0.30844778,0.3435874,0.37872702,0.41386664,0.44900626,0.48414588,0.5192855,0.5544251,0.58956474,0.62470436,0.6676528,0.7106012,0.75354964,0.79649806,0.8394465,0.8862993,0.93315214,0.98000497,1.0268579,1.0737107,1.1791295,1.2806439,1.3821584,1.4836729,1.5890918,1.8584955,2.1278992,2.397303,2.6667068,2.9361105,2.8619268,2.787743,2.7135596,2.639376,2.5612879,2.7135596,2.8658314,3.018103,3.174279,3.3265507,3.408543,3.49444,3.5803368,3.6662338,3.7482262,3.533484,3.3187418,3.1039999,2.8892577,2.6745155,3.0102942,3.3460727,3.6818514,4.0137253,4.349504,4.5564375,4.759466,4.9663997,5.169429,5.376362,5.376362,5.376362,5.376362,5.376362,5.376362,5.6652875,5.9542136,6.2431393,6.5359693,6.824895,7.2543793,7.6799593,8.109444,8.535024,8.960603,8.52331,8.082112,7.6409154,7.2036223,6.7624245,6.7429028,6.7233806,6.703859,6.6843367,6.66091,6.621866,6.578918,6.5359693,6.493021,6.4500723,6.3407493,6.2314262,6.1181984,6.008875,5.899552,5.801942,5.700427,5.5989127,5.5013027,5.3997884,5.337318,5.2748475,5.212377,5.1499066,5.087436,5.290465,5.493494,5.6965227,5.8956475,6.098676,6.126007,6.153338,6.180669,6.211904,6.239235,6.4969254,6.7507114,7.008402,7.266093,7.523783,7.570636,7.621393,7.6682463,7.715099,7.7619514,7.5433054,7.328563,7.1099167,6.89127,6.676528,7.3129454,7.9493628,8.58578,9.226103,9.86252,10.42085,10.983084,11.541413,12.103647,12.661977,14.313539,15.969006,17.620567,19.27213,20.92369,24.10578,27.283962,30.466051,33.644234,36.82632,34.054195,31.285975,28.51385,25.745628,22.973503,19.971018,16.968533,13.966047,10.963562,7.9610763,6.8561306,5.74728,4.6384296,3.533484,2.4246337,1.9404879,1.456342,0.96829176,0.48414588,0.0,0.29673457,0.58956474,0.8862993,1.1791295,1.475864,1.1791295,0.8862993,0.58956474,0.29673457,0.0,0.0,0.0,0.0,0.0,0.0,0.31625658,0.63641757,0.95267415,1.2689307,1.5890918,1.7491722,1.9092526,2.069333,2.2294137,2.3855898,2.1708477,1.9522011,1.7335546,1.5188124,1.3001659,1.4016805,1.5031948,1.6086137,1.7101282,1.8116426,1.4485333,1.0893283,0.7262188,0.3631094,0.0,1.3509232,2.7018464,4.0488653,5.3997884,6.7507114,6.1299114,5.5091114,4.8883114,4.271416,3.6506162,3.521771,3.3890212,3.260176,3.1313305,2.998581,3.0532427,3.1039999,3.1586614,3.2094188,3.2640803,4.2089458,5.153811,6.098676,7.043542,7.988407,8.535024,9.081639,9.628256,10.178777,10.725393,10.545791,10.370092,10.194394,10.0147915,9.839094,8.886419,7.9376497,6.98888,6.036206,5.087436,4.9546866,4.8219366,4.689187,4.5564375,4.423688,4.4119744,4.4002614,4.388548,4.376835,4.3612175,4.173806,3.9824903,3.7911747,3.6037633,3.4124475,3.408543,3.408543,3.4046388,3.4007344,3.4007344,3.6545205,3.9083066,4.165997,4.4197836,4.6735697,3.9824903,3.2914112,2.5964274,1.9053483,1.2142692,1.358732,1.5070993,1.6554666,1.8038338,1.9482968,2.182561,2.416825,2.6471848,2.8814487,3.1118085,3.1157131,3.1235218,3.1274261,3.1313305,3.1391394,2.9907722,2.8424048,2.6940374,2.5456703,2.4012074,2.3738766,2.35045,2.3231194,2.2996929,2.2762666,2.084951,1.893635,1.7062237,1.5149081,1.3235924,1.1478943,0.96829176,0.79259366,0.61689556,0.43729305,0.4997635,0.5622339,0.62470436,0.6871748,0.74964523,0.93315214,1.116659,1.2962615,1.4797685,1.6632754,1.8506867,2.0380979,2.2255092,2.4129205,2.6003318,2.5183394,2.4402514,2.358259,2.280171,2.1981785,2.1708477,2.1396124,2.1083772,2.0810463,2.0498111,1.639849,1.2298868,0.8199245,0.40996224,0.0,2.5690966,5.134289,7.703386,10.268578,12.837675,10.936231,9.0386915,7.137247,5.2358036,3.338264,8.413987,13.493614,18.569338,23.648964,28.724688,24.539167,20.35365,16.168129,11.986515,7.800996,8.929368,10.053836,11.182208,12.31058,13.438952,12.661977,11.888905,11.111929,10.338858,9.561881,8.929368,8.292951,7.656533,7.0240197,6.387602,6.04011,5.6926184,5.3451266,4.997635,4.650143,5.165524,5.6809053,6.196286,6.7116675,7.223144,6.8287997,6.4305506,6.0323014,5.6340523,5.2358036,4.9742084,4.7126136,4.4510183,4.1894236,3.9239242,3.8692627,3.814601,3.7599394,3.7052777,3.6506162,3.78727,3.9239242,4.0605783,4.2011366,4.337791,4.8687897,5.395884,5.9268827,6.4578815,6.98888,6.9068875,6.8209906,6.7389984,6.657006,6.575013,6.703859,6.8366084,6.9654536,7.094299,7.223144,6.2587566,5.290465,4.322173,3.3538816,2.3855898,2.0810463,1.7725986,1.4641509,1.1557031,0.8511597,0.679366,0.5114767,0.339683,0.1717937,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,1.0893283,2.1161861,3.1469483,4.173806,5.2006636,5.5169206,5.8292727,6.1455293,6.461786,6.774138,6.250948,5.7238536,5.2006636,4.6735697,4.1503797,3.716991,3.2836022,2.854118,2.4207294,1.9873407,1.8623998,1.737459,1.6125181,1.4875772,1.3626363,1.698415,2.0341935,2.366068,2.7018464,3.0376248,2.9556324,2.87364,2.7916477,2.7057507,2.6237583,2.3816853,2.135708,1.8897307,1.6437533,1.4016805,1.43682,1.4680552,1.5031948,1.5383345,1.5734742,1.8116426,2.0459068,2.280171,2.514435,2.7486992,2.4910088,2.233318,1.9756275,1.7218413,1.4641509,1.2884527,1.1127546,0.93705654,0.76135844,0.58566034,0.48414588,0.37872702,0.27330816,0.1678893,0.062470436,0.80821127,1.5539521,2.2957885,3.0415294,3.78727,3.5608149,3.3343596,3.1039999,2.8775444,2.6510892,3.5569105,4.4588275,5.364649,6.27047,7.1762915,6.9264097,6.6804323,6.4305506,6.184573,5.938596,6.1455293,6.3524623,6.559396,6.7663293,6.9732623,7.2075267,7.4417906,7.6721506,7.9064145,8.136774,8.800523,9.464272,10.124115,10.787864,11.4516115,10.303718,9.159728,8.015738,6.871748,5.7238536,4.7789884,3.8341231,2.8892577,1.9443923,0.999527,1.2689307,1.53443,1.8038338,2.069333,2.338737,2.0341935,1.7335546,1.4290112,1.1283722,0.8238289,0.80430686,0.78088045,0.75745404,0.7340276,0.7106012,0.6481308,0.58566034,0.5231899,0.46071947,0.39824903,0.79649806,1.1908426,1.5851873,1.979532,2.3738766,2.338737,2.2996929,2.260649,2.2255092,2.1864653,2.3543546,2.5183394,2.6823244,2.8463092,3.0141985,2.8892577,2.7682211,2.6432803,2.522244,2.4012074,2.2684577,2.135708,2.0029583,1.8702087,1.737459,0.43729305,0.63641757,0.8355421,1.038571,1.2376955,1.43682,2.0263848,2.612045,3.2016098,3.78727,4.376835,4.4510183,4.5252023,4.5993857,4.6735697,4.7516575,4.575959,4.4002614,4.224563,4.0488653,3.873167,3.513962,3.1508527,2.787743,2.4246337,2.0615244,1.901444,1.737459,1.5734742,1.4133936,1.2494087,1.1869383,1.1244678,1.0619974,0.999527,0.93705654,0.8745861,0.81211567,0.74964523,0.6871748,0.62470436,0.63641757,0.6481308,0.6637484,0.6754616,0.6871748,0.76135844,0.8394465,0.9136301,0.9878138,1.0619974,0.9136301,0.76135844,0.61299115,0.46071947,0.31235218,0.61299115,0.9136301,1.2142692,1.5110037,1.8116426,1.5110037,1.2142692,0.9136301,0.61299115,0.31235218,0.3240654,0.3357786,0.3513962,0.3631094,0.37482262,0.38653582,0.39824903,0.41386664,0.42557985,0.43729305,0.3631094,0.28892577,0.21083772,0.13665408,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.22645533,0.26159495,0.30063897,0.3357786,0.37482262,0.41386664,0.44900626,0.48805028,0.5231899,0.5622339,0.61299115,0.6637484,0.7106012,0.76135844,0.81211567,0.92534333,1.038571,1.1517987,1.261122,1.3743496,1.6359446,1.901444,2.1630387,2.4246337,2.6862288,2.6003318,2.514435,2.4246337,2.338737,2.2489357,2.4871042,2.7252727,2.9634414,3.2016098,3.435874,3.513962,3.5881457,3.6623292,3.736513,3.8106966,3.5256753,3.2367494,2.951728,2.6628022,2.3738766,2.7994564,3.2250361,3.6506162,4.0761957,4.5017757,4.7633705,5.024966,5.2865605,5.548156,5.813655,5.801942,5.786324,5.774611,5.7628975,5.7511845,6.036206,6.3251314,6.6140575,6.899079,7.1880045,7.7385254,8.289046,8.835662,9.386183,9.936704,9.413514,8.886419,8.36323,7.8361354,7.3129454,7.3246584,7.336372,7.348085,7.363703,7.375416,7.348085,7.3246584,7.3012323,7.2739015,7.250475,7.08649,6.9264097,6.7624245,6.5984397,6.4383593,6.2860875,6.13772,5.989353,5.8370814,5.688714,5.548156,5.4115014,5.2748475,5.138193,5.001539,5.263134,5.5247293,5.786324,6.0518236,6.3134184,6.3017054,6.2860875,6.2743745,6.262661,6.250948,6.5359693,6.824895,7.113821,7.3988423,7.687768,7.7502384,7.812709,7.8751793,7.9376497,8.00012,7.7111945,7.426173,7.137247,6.8483214,6.5633,7.3129454,8.062591,8.812236,9.561881,10.311526,11.0260315,11.736633,12.4511385,13.16174,13.8762455,15.449719,17.023193,18.600573,20.174046,21.751425,25.300526,28.849628,32.39873,35.951736,39.50084,36.13915,32.773552,29.411861,26.05017,22.688482,19.400974,16.113468,12.825961,9.538455,6.250948,5.001539,3.7482262,2.4988174,1.2494087,0.0,0.0,0.0,0.0,0.0,0.0,0.13665408,0.27330816,0.41386664,0.5505207,0.6871748,0.5505207,0.41386664,0.27330816,0.13665408,0.0,0.0,0.0,0.0,0.0,0.0,0.38653582,0.77307165,1.1635119,1.5500476,1.9365835,2.0263848,2.1122816,2.1981785,2.2879796,2.3738766,1.9248703,1.475864,1.0268579,0.57394713,0.12494087,0.5231899,0.92534333,1.3235924,1.7257458,2.1239948,1.698415,1.2767396,0.8511597,0.42557985,0.0,1.6867018,3.3734035,5.0640097,6.7507114,8.437413,7.6643414,6.8873653,6.114294,5.337318,4.564246,4.4002614,4.2362766,4.0761957,3.912211,3.7482262,3.5998588,3.4514916,3.2992198,3.1508527,2.998581,4.1620927,5.3256044,6.4891167,7.648724,8.812236,9.198771,9.589212,9.975748,10.362284,10.748819,10.81129,10.87376,10.936231,10.998701,11.061172,10.073358,9.089449,8.101635,7.113821,6.126007,5.8370814,5.548156,5.263134,4.9742084,4.689187,4.650143,4.6110992,4.575959,4.5369153,4.5017757,4.263607,4.025439,3.78727,3.5491016,3.310933,3.1000953,2.8892577,2.6745155,2.463678,2.2489357,2.5886188,2.9243972,3.2640803,3.5998588,3.9356375,3.2250361,2.514435,1.7999294,1.0893283,0.37482262,0.63641757,0.9019169,1.1635119,1.4251068,1.6867018,1.8116426,1.9365835,2.0615244,2.1864653,2.3114061,2.2879796,2.260649,2.2372224,2.2137961,2.1864653,2.2255092,2.260649,2.2996929,2.338737,2.3738766,2.3855898,2.4012074,2.4129205,2.4246337,2.436347,2.1513257,1.8623998,1.5734742,1.2884527,0.999527,0.8238289,0.6481308,0.47633708,0.30063897,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.3357786,0.5505207,0.76135844,0.97610056,1.1869383,1.3235924,1.4641509,1.6008049,1.737459,1.8741131,1.999054,2.1239948,2.2489357,2.3738766,2.4988174,2.4012074,2.2996929,2.1981785,2.1005683,1.999054,1.6008049,1.1986516,0.80040246,0.39824903,0.0,3.174279,6.348558,9.526741,12.70102,15.875299,12.974329,10.073358,7.1762915,4.2753205,1.3743496,7.824422,14.274494,20.724567,27.17464,33.624714,28.486519,23.348326,18.214037,13.075843,7.9376497,8.976221,10.010887,11.0494585,12.08803,13.1266,12.4745655,11.826434,11.174399,10.526268,9.874233,9.101162,8.324185,7.551114,6.774138,6.001066,5.5130157,5.024966,4.5369153,4.0488653,3.5608149,4.337791,5.1108627,5.8878384,6.66091,7.437886,7.0357327,6.6374836,6.239235,5.8370814,5.4388323,5.173333,4.911738,4.650143,4.388548,4.123049,4.2011366,4.2753205,4.349504,4.423688,4.5017757,4.6110992,4.7243266,4.8375545,4.950782,5.0640097,5.6262436,6.1884775,6.7507114,7.3129454,7.8751793,7.551114,7.223144,6.899079,6.575013,6.250948,6.4500723,6.649197,6.8483214,7.0513506,7.250475,6.1494336,5.0483923,3.951255,2.8502135,1.7491722,1.5266213,1.3001659,1.0737107,0.8511597,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.0,0.0,0.0,0.0,0.0,0.0,1.1361811,2.2762666,3.4124475,4.548629,5.688714,5.099149,4.513489,3.9239242,3.338264,2.7486992,2.8385005,2.9243972,3.0141985,3.1000953,3.1859922,2.6628022,2.135708,1.6125181,1.0893283,0.5622339,0.5231899,0.48805028,0.44900626,0.41386664,0.37482262,0.8394465,1.3001659,1.7608855,2.2255092,2.6862288,2.612045,2.5378613,2.463678,2.3855898,2.3114061,2.1239948,1.9365835,1.7491722,1.5617609,1.3743496,1.3509232,1.3235924,1.3001659,1.2767396,1.2494087,1.4875772,1.7257458,1.9639144,2.1981785,2.436347,2.2137961,1.9873407,1.7608855,1.5383345,1.3118792,1.1517987,0.9878138,0.8238289,0.6637484,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.77697605,1.5500476,2.3231194,3.1000953,3.873167,3.5373883,3.2016098,2.8619268,2.5261483,2.1864653,3.0883822,3.9863946,4.8883114,5.786324,6.688241,6.5008297,6.3134184,6.126007,5.938596,5.7511845,6.098676,6.4500723,6.801469,7.1489606,7.5003567,7.5120697,7.523783,7.5394006,7.551114,7.562827,8.113348,8.663869,9.21439,9.761005,10.311526,9.261242,8.210958,7.1606736,6.114294,5.0640097,4.1503797,3.2367494,2.3231194,1.4133936,0.4997635,0.77307165,1.0502841,1.3235924,1.6008049,1.8741131,1.5500476,1.2259823,0.9019169,0.57394713,0.24988174,0.23816854,0.22645533,0.21083772,0.19912452,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.41386664,0.76135844,1.1127546,1.4641509,1.8116426,1.901444,1.9873407,2.0732377,2.1630387,2.2489357,2.4988174,2.7486992,2.998581,3.2484627,3.4983444,3.338264,3.174279,3.0141985,2.8502135,2.6862288,2.5495746,2.4129205,2.2762666,2.135708,1.999054,0.5622339,0.7223144,0.8823949,1.0424755,1.2025559,1.3626363,1.815547,2.2723622,2.7291772,3.182088,3.638903,3.68966,3.7443218,3.795079,3.8458362,3.900498,3.7560349,3.611572,3.4632049,3.3187418,3.174279,2.8814487,2.5847144,2.2918842,1.9951496,1.698415,1.5890918,1.475864,1.3626363,1.2494087,1.1361811,1.116659,1.0932326,1.0698062,1.0463798,1.0268579,0.94876975,0.8745861,0.80040246,0.7262188,0.6481308,0.659844,0.6715572,0.679366,0.6910792,0.698888,0.7340276,0.76916724,0.80430686,0.8394465,0.8745861,0.76916724,0.659844,0.5544251,0.44510186,0.3357786,0.62860876,0.92143893,1.2142692,1.5070993,1.7999294,1.542239,1.2845483,1.0268579,0.76916724,0.5114767,0.48414588,0.45291066,0.42167544,0.39434463,0.3631094,0.37872702,0.39434463,0.40605783,0.42167544,0.43729305,0.3631094,0.28892577,0.21083772,0.13665408,0.062470436,0.07027924,0.078088045,0.08589685,0.093705654,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05466163,0.058566034,0.058566034,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.21864653,0.24597734,0.27721256,0.30844778,0.3357786,0.3670138,0.39824903,0.42557985,0.45681506,0.48805028,0.5309987,0.57394713,0.61689556,0.6559396,0.698888,0.79259366,0.8862993,0.97610056,1.0698062,1.1635119,1.3743496,1.5812829,1.7921207,2.0029583,2.2137961,2.1474214,2.0810463,2.018576,1.9522011,1.8858263,2.0927596,2.2957885,2.5027218,2.7057507,2.912684,3.0259118,3.1430438,3.2562714,3.3734035,3.4866312,3.2094188,2.9322062,2.6549935,2.377781,2.1005683,2.4910088,2.8853533,3.2757936,3.6701381,4.0605783,4.388548,4.7126136,5.036679,5.3607445,5.688714,5.6262436,5.5676775,5.5091114,5.446641,5.388075,5.64967,5.911265,6.1767645,6.4383593,6.699954,7.1333427,7.570636,8.0040245,8.441318,8.874706,8.488171,8.101635,7.7111945,7.3246584,6.9381227,6.9732623,7.012306,7.0513506,7.08649,7.125534,7.223144,7.320754,7.4183645,7.5159745,7.6135845,7.57454,7.5394006,7.5003567,7.461313,7.426173,7.195813,6.969358,6.7429028,6.5164475,6.2860875,6.1611466,6.036206,5.911265,5.786324,5.661383,5.891743,6.1221027,6.3524623,6.5828223,6.813182,6.7311897,6.649197,6.5633,6.481308,6.3993154,6.6843367,6.969358,7.2543793,7.5394006,7.824422,7.8361354,7.8517528,7.8634663,7.8751793,7.8868923,7.7229075,7.558923,7.3910336,7.2270484,7.0630636,7.7775693,8.492075,9.20658,9.921086,10.6355915,11.303245,11.966993,12.630741,13.298394,13.962143,15.051471,16.140799,17.234032,18.32336,19.412687,23.531832,27.647072,31.766216,35.88146,40.000603,36.02592,32.05124,28.076557,24.101875,20.12329,17.132517,14.141745,11.147068,8.156297,5.1616197,4.142571,3.1235218,2.1005683,1.0815194,0.062470436,0.07418364,0.08199245,0.093705654,0.10151446,0.113227665,0.32016098,0.5270943,0.7340276,0.94096094,1.1517987,0.92143893,0.6910792,0.46071947,0.23035973,0.0,0.0,0.0,0.0,0.0,0.0,0.3670138,0.7340276,1.1010414,1.4680552,1.8389735,1.8545911,1.8741131,1.8897307,1.9092526,1.9248703,1.5617609,1.1947471,0.8316377,0.46462387,0.10151446,0.42167544,0.7418364,1.0580931,1.3782539,1.698415,1.358732,1.0190489,0.679366,0.339683,0.0,2.0537157,4.1035266,6.1572423,8.210958,10.260769,9.101162,7.9376497,6.774138,5.610626,4.4510183,4.165997,3.8809757,3.5959544,3.310933,3.0259118,2.9361105,2.8463092,2.7565079,2.6667068,2.5769055,3.7013733,4.825841,5.950309,7.0747766,8.1992445,8.738052,9.276859,9.811763,10.350571,10.889378,10.916709,10.947944,10.979179,11.00651,11.037745,10.264673,9.491602,8.718531,7.9493628,7.1762915,6.801469,6.4305506,6.055728,5.6848097,5.3138914,5.173333,5.036679,4.900025,4.7633705,4.6267166,4.388548,4.1503797,3.912211,3.6740425,3.435874,3.1781836,2.9243972,2.6667068,2.4090161,2.1513257,2.3621633,2.5769055,2.787743,2.998581,3.213323,2.7057507,2.2020829,1.698415,1.1908426,0.6871748,0.9058213,1.1283722,1.3470187,1.5656652,1.7882162,1.8038338,1.8233559,1.8389735,1.8584955,1.8741131,1.9404879,2.0068626,2.069333,2.135708,2.1981785,2.3075018,2.416825,2.522244,2.631567,2.736986,2.6042364,2.4714866,2.338737,2.2059872,2.0732377,1.8467822,1.6164225,1.3860629,1.1557031,0.92534333,0.77307165,0.62470436,0.47633708,0.3240654,0.1756981,0.1717937,0.1639849,0.16008049,0.15617609,0.14836729,0.3357786,0.5192855,0.7066968,0.8902037,1.0737107,1.2181735,1.358732,1.5031948,1.6437533,1.7882162,1.9131571,2.0420024,2.1708477,2.2957885,2.4246337,2.2645533,2.1044729,1.9443923,1.7843118,1.6242313,1.3001659,0.97610056,0.6481308,0.3240654,0.0,2.541766,5.0796275,7.621393,10.159255,12.70102,10.545791,8.3944645,6.2431393,4.0918136,1.9365835,7.2465706,12.556558,17.866545,23.176533,28.486519,24.062832,19.643047,15.21936,10.795672,6.375889,7.7541428,9.128492,10.506746,11.885,13.263254,12.201257,11.139259,10.073358,9.01136,7.9493628,8.413987,8.878611,9.343235,9.811763,10.276386,8.941081,7.60968,6.278279,4.9468775,3.611572,4.3338866,5.0522966,5.7707067,6.493021,7.211431,6.89127,6.571109,6.250948,5.930787,5.610626,5.423215,5.2358036,5.0483923,4.860981,4.6735697,4.6696653,4.6657605,4.661856,4.6540475,4.650143,4.73604,4.825841,4.911738,5.001539,5.087436,5.481781,5.872221,6.266566,6.657006,7.0513506,6.75852,6.4695945,6.180669,5.891743,5.5989127,5.735567,5.8761253,6.012779,6.1494336,6.2860875,5.309987,4.3338866,3.3538816,2.377781,1.4016805,1.2181735,1.038571,0.8589685,0.679366,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.0,0.0,0.0,0.0,0.0,0.9097257,1.8194515,2.7291772,3.638903,4.548629,4.084005,3.6154766,3.1469483,2.67842,2.2137961,2.3348327,2.455869,2.5808098,2.7018464,2.8267872,2.3933985,1.9600099,1.5266213,1.0932326,0.6637484,0.7066968,0.75354964,0.79649806,0.8433509,0.8862993,1.1635119,1.43682,1.7140326,1.9873407,2.260649,2.1786566,2.096664,2.0146716,1.9326792,1.8506867,1.698415,1.5500476,1.4016805,1.2494087,1.1010414,1.0932326,1.0893283,1.0854238,1.0815194,1.0737107,1.2533131,1.43682,1.6164225,1.796025,1.9756275,1.7882162,1.6047094,1.4212024,1.2337911,1.0502841,0.93315214,0.8160201,0.698888,0.58175594,0.46071947,0.3709182,0.27721256,0.1835069,0.093705654,0.0,0.737932,1.475864,2.2137961,2.951728,3.6857557,3.4280653,3.174279,2.9165885,2.6588979,2.4012074,3.3187418,4.240181,5.1616197,6.0791545,7.000593,6.813182,6.6257706,6.4383593,6.250948,6.0635366,6.3173227,6.571109,6.8287997,7.082586,7.336372,7.4183645,7.504261,7.5862536,7.6682463,7.7502384,8.066495,8.386656,8.702912,9.019169,9.339331,8.495979,7.656533,6.817086,5.9776397,5.138193,4.3260775,3.513962,2.7018464,1.8858263,1.0737107,1.3274968,1.5812829,1.8311646,2.084951,2.338737,2.0107672,1.6867018,1.3626363,1.038571,0.7106012,0.7027924,0.6910792,0.6832704,0.6715572,0.6637484,0.60908675,0.5544251,0.4958591,0.44119745,0.38653582,0.9136301,1.4407244,1.9717231,2.4988174,3.0259118,3.0220075,3.018103,3.018103,3.0141985,3.0141985,3.2445583,3.4788225,3.7091823,3.9434462,4.173806,3.970777,3.7638438,3.5608149,3.3538816,3.1508527,2.8814487,2.6159496,2.3465457,2.0810463,1.8116426,0.6871748,0.80821127,0.92924774,1.0463798,1.1674163,1.2884527,1.6086137,1.9326792,2.2567444,2.5769055,2.900971,2.9283018,2.959537,2.9907722,3.018103,3.049338,2.9361105,2.8189783,2.7057507,2.5886188,2.475391,2.2489357,2.018576,1.7921207,1.5656652,1.33921,1.2767396,1.2142692,1.1517987,1.0893283,1.0268579,1.0424755,1.0580931,1.077615,1.0932326,1.1127546,1.0268579,0.93705654,0.8511597,0.76135844,0.6754616,0.6832704,0.6910792,0.698888,0.7066968,0.7106012,0.7066968,0.7027924,0.698888,0.6910792,0.6871748,0.62079996,0.5583295,0.49195468,0.42557985,0.3631094,0.6481308,0.93315214,1.2181735,1.5031948,1.7882162,1.5734742,1.358732,1.1439898,0.92924774,0.7106012,0.64032197,0.5661383,0.4958591,0.42167544,0.3513962,0.3670138,0.38653582,0.40215343,0.42167544,0.43729305,0.3631094,0.28892577,0.21083772,0.13665408,0.062470436,0.06637484,0.06637484,0.07027924,0.07418364,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.042948425,0.046852827,0.05075723,0.058566034,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.21083772,0.23426414,0.25378615,0.27721256,0.30063897,0.3240654,0.3435874,0.3670138,0.39044023,0.41386664,0.44900626,0.48414588,0.5192855,0.5544251,0.58566034,0.659844,0.7340276,0.80430686,0.8784905,0.94876975,1.1088502,1.2650263,1.4212024,1.5812829,1.737459,1.6945106,1.6515622,1.6086137,1.5656652,1.5266213,1.698415,1.8702087,2.0420024,2.2137961,2.3855898,2.541766,2.697942,2.854118,3.0063896,3.1625657,2.893162,2.6276627,2.358259,2.0927596,1.8233559,2.1864653,2.5456703,2.9048753,3.2640803,3.6232853,4.0137253,4.4002614,4.786797,5.173333,5.563773,5.45445,5.349031,5.239708,5.134289,5.024966,5.263134,5.5013027,5.735567,5.9737353,6.211904,6.532065,6.852226,7.172387,7.492548,7.812709,7.562827,7.3129454,7.0630636,6.813182,6.5633,6.6257706,6.688241,6.7507114,6.813182,6.8756523,7.094299,7.3168497,7.535496,7.7541428,7.9766936,8.062591,8.148487,8.238289,8.324185,8.413987,8.109444,7.800996,7.4964523,7.191909,6.8873653,6.774138,6.66091,6.551587,6.4383593,6.3251314,6.524256,6.719476,6.918601,7.113821,7.3129454,7.1606736,7.008402,6.8561306,6.703859,6.551587,6.832704,7.113821,7.3988423,7.6799593,7.9610763,7.9259367,7.8868923,7.8517528,7.812709,7.773665,7.7307167,7.6916723,7.648724,7.605776,7.562827,8.242193,8.921559,9.600925,10.284196,10.963562,11.580457,12.197352,12.814248,13.431144,14.051944,14.653222,15.258404,15.863586,16.46877,17.073952,21.759233,26.444517,31.129799,35.815083,40.500366,35.912693,31.32502,26.737347,22.149673,17.562002,14.864059,12.166118,9.468176,6.774138,4.0761957,3.2836022,2.494913,1.7062237,0.9136301,0.12494087,0.14446288,0.1639849,0.1835069,0.20693332,0.22645533,0.5036679,0.78088045,1.0580931,1.3353056,1.6125181,1.2884527,0.96829176,0.6442264,0.3240654,0.0,0.0,0.0,0.0,0.0,0.0,0.3474918,0.6949836,1.0424755,1.3899672,1.737459,1.6867018,1.6320401,1.5812829,1.5266213,1.475864,1.1947471,0.9136301,0.63641757,0.3553006,0.07418364,0.31625658,0.5544251,0.79649806,1.0346665,1.2767396,1.0190489,0.76526284,0.5114767,0.25378615,0.0,2.416825,4.83365,7.2543793,9.671205,12.08803,10.537982,8.987934,7.437886,5.8878384,4.337791,3.9317331,3.521771,3.1157131,2.7057507,2.2996929,2.2684577,2.241127,2.2098918,2.1786566,2.1513257,3.2367494,4.3260775,5.4115014,6.5008297,7.5862536,8.273428,8.960603,9.651682,10.338858,11.0260315,11.022127,11.018223,11.018223,11.014318,11.014318,10.455989,9.897659,9.339331,8.781001,8.226576,7.7658563,7.309041,6.852226,6.395411,5.938596,5.700427,5.462259,5.22409,4.985922,4.7516575,4.513489,4.2753205,4.037152,3.7989833,3.5608149,3.260176,2.9556324,2.6549935,2.3543546,2.0498111,2.135708,2.2255092,2.3114061,2.4012074,2.4871042,2.1903696,1.893635,1.5969005,1.2962615,0.999527,1.1791295,1.3548276,1.53443,1.7101282,1.8858263,1.796025,1.7062237,1.6164225,1.5266213,1.43682,1.5929961,1.7491722,1.901444,2.05762,2.2137961,2.3894942,2.5690966,2.7447948,2.9243972,3.1000953,2.822883,2.5456703,2.2684577,1.9912452,1.7140326,1.5383345,1.3665408,1.1947471,1.0229534,0.8511597,0.7262188,0.60127795,0.47633708,0.3513962,0.22645533,0.21474212,0.20693332,0.19522011,0.1835069,0.1756981,0.3318742,0.48805028,0.6481308,0.80430686,0.96438736,1.1088502,1.2572175,1.4055848,1.5539521,1.698415,1.8311646,1.9600099,2.0888553,2.2216048,2.35045,2.1318035,1.9092526,1.6906061,1.4680552,1.2494087,0.999527,0.74964523,0.4997635,0.24988174,0.0,1.9053483,3.8106966,5.716045,7.621393,9.526741,8.121157,6.715572,5.309987,3.9044023,2.4988174,6.6687193,10.838621,15.008522,19.178425,23.348326,19.643047,15.933866,12.228588,8.519405,4.814128,6.5281606,8.246098,9.964035,11.681972,13.399908,11.924045,10.44818,8.976221,7.5003567,6.0244927,7.7307167,9.433036,11.139259,12.845484,14.551707,12.373051,10.194394,8.015738,5.840986,3.6623292,4.3260775,4.9937305,5.657479,6.321227,6.98888,6.746807,6.5086384,6.266566,6.028397,5.786324,5.6730967,5.563773,5.4505453,5.337318,5.22409,5.138193,5.056201,4.970304,4.884407,4.7985106,4.860981,4.9234514,4.985922,5.0483923,5.1108627,5.3334136,5.5559645,5.7785153,6.001066,6.223617,5.969831,5.716045,5.4583545,5.2045684,4.950782,5.024966,5.099149,5.173333,5.251421,5.3256044,4.4705405,3.6154766,2.7604125,1.9053483,1.0502841,0.9136301,0.78088045,0.6442264,0.5114767,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.6832704,1.3665408,2.0459068,2.7291772,3.4124475,3.0649557,2.717464,2.3699722,2.0224805,1.6749885,1.8311646,1.9912452,2.1474214,2.3035975,2.463678,2.1239948,1.7843118,1.4407244,1.1010414,0.76135844,0.8902037,1.0190489,1.1439898,1.2728351,1.4016805,1.4875772,1.5734742,1.6632754,1.7491722,1.8389735,1.7491722,1.6593709,1.5656652,1.475864,1.3860629,1.2767396,1.1635119,1.0502841,0.93705654,0.8238289,0.8394465,0.8550641,0.8706817,0.8862993,0.9019169,1.0229534,1.1439898,1.2689307,1.3899672,1.5110037,1.3665408,1.2220778,1.077615,0.93315214,0.78868926,0.7145056,0.6442264,0.5700427,0.4958591,0.42557985,0.339683,0.25378615,0.1717937,0.08589685,0.0,0.698888,1.4016805,2.1005683,2.7994564,3.4983444,3.3226464,3.1469483,2.9673457,2.7916477,2.612045,3.5530062,4.493967,5.4310236,6.3719845,7.3129454,7.125534,6.9381227,6.7507114,6.5633,6.375889,6.5359693,6.6960497,6.8561306,7.016211,7.1762915,7.328563,7.480835,7.633106,7.785378,7.9376497,8.023546,8.109444,8.191436,8.277332,8.36323,7.7307167,7.1021075,6.473499,5.840986,5.212377,4.5017757,3.78727,3.076669,2.3621633,1.6515622,1.8819219,2.1083772,2.338737,2.5690966,2.7994564,2.475391,2.1513257,1.8233559,1.4992905,1.175225,1.1674163,1.1596074,1.1517987,1.1439898,1.1361811,1.0541886,0.96829176,0.8823949,0.79649806,0.7106012,1.4172981,2.1239948,2.8267872,3.533484,4.2362766,4.1464753,4.0527697,3.959064,3.8692627,3.775557,3.9902992,4.2050414,4.4197836,4.6345253,4.8492675,4.60329,4.3534083,4.1074314,3.8614538,3.611572,3.213323,2.8189783,2.4207294,2.0224805,1.6242313,0.81211567,0.8941081,0.97219616,1.0541886,1.1322767,1.2142692,1.4016805,1.5929961,1.7843118,1.9717231,2.1630387,2.1708477,2.1786566,2.1864653,2.194274,2.1981785,2.1161861,2.0302892,1.9443923,1.8584955,1.7765031,1.6164225,1.456342,1.2962615,1.1361811,0.97610056,0.96438736,0.94876975,0.93705654,0.92534333,0.9136301,0.96829176,1.0268579,1.0854238,1.1439898,1.1986516,1.1010414,0.999527,0.9019169,0.80040246,0.698888,0.7066968,0.7106012,0.7145056,0.71841,0.7262188,0.679366,0.63641757,0.58956474,0.5466163,0.4997635,0.47633708,0.45681506,0.43338865,0.40996224,0.38653582,0.6637484,0.94096094,1.2181735,1.4992905,1.7765031,1.6008049,1.4290112,1.2572175,1.0854238,0.9136301,0.79649806,0.6832704,0.5661383,0.45291066,0.3357786,0.359205,0.37872702,0.39824903,0.41777104,0.43729305,0.3631094,0.28892577,0.21083772,0.13665408,0.062470436,0.058566034,0.058566034,0.05466163,0.05075723,0.05075723,0.046852827,0.039044023,0.03513962,0.031235218,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.031235218,0.039044023,0.046852827,0.05466163,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.20302892,0.21864653,0.23426414,0.24597734,0.26159495,0.27721256,0.29283017,0.30844778,0.3240654,0.3357786,0.3631094,0.39434463,0.42167544,0.44900626,0.47633708,0.5270943,0.58175594,0.63251317,0.6832704,0.737932,0.8433509,0.94876975,1.0541886,1.1557031,1.261122,1.2415999,1.2220778,1.2025559,1.183034,1.1635119,1.3040704,1.4407244,1.5812829,1.7218413,1.8623998,2.05762,2.25284,2.4480603,2.6432803,2.8385005,2.5808098,2.3231194,2.0654287,1.8077383,1.5500476,1.8780174,2.2059872,2.533957,2.8619268,3.1859922,3.638903,4.087909,4.5369153,4.985922,5.4388323,5.282656,5.12648,4.9742084,4.8180323,4.661856,4.8765984,5.087436,5.298274,5.5130157,5.7238536,5.930787,6.133816,6.3407493,6.5437784,6.7507114,6.6374836,6.524256,6.4110284,6.3017054,6.1884775,6.2743745,6.364176,6.4500723,6.5359693,6.6257706,6.969358,7.309041,7.6526284,7.996216,8.335898,8.550641,8.761478,8.976221,9.187058,9.4018,9.019169,8.636538,8.253906,7.871275,7.4886436,7.387129,7.2856145,7.1880045,7.08649,6.98888,7.152865,7.3168497,7.480835,7.648724,7.812709,7.590158,7.367607,7.1450562,6.9225054,6.699954,6.9810715,7.2582836,7.5394006,7.8205175,8.101635,8.011833,7.9259367,7.8361354,7.7502384,7.6643414,7.7424297,7.824422,7.90251,7.9805984,8.062591,8.706817,9.351044,9.999174,10.6434,11.287627,11.85767,12.427712,12.997755,13.567798,14.13784,14.258877,14.376009,14.4970455,14.618082,14.739119,19.99054,25.24196,30.493382,35.748707,41.00013,35.799465,30.5988,25.398136,20.201378,15.000713,12.595602,10.194394,7.793187,5.388075,2.9868677,2.4285383,1.8663043,1.3079748,0.74574083,0.18741131,0.21864653,0.24597734,0.27721256,0.30844778,0.3357786,0.6832704,1.0307622,1.3782539,1.7257458,2.0732377,1.6593709,1.2455044,0.8316377,0.41386664,0.0,0.0,0.0,0.0,0.0,0.0,0.3279698,0.6559396,0.98390937,1.3118792,1.6359446,1.5149081,1.3938715,1.2689307,1.1478943,1.0268579,0.8316377,0.63641757,0.44119745,0.24597734,0.05075723,0.21083772,0.3709182,0.5309987,0.6910792,0.8511597,0.679366,0.5114767,0.339683,0.1717937,0.0,2.7838387,5.563773,8.347612,11.131451,13.911386,11.974802,10.0382185,8.101635,6.1611466,4.224563,3.6935644,3.1664703,2.6354716,2.1044729,1.5734742,1.6047094,1.6359446,1.6632754,1.6945106,1.7257458,2.77603,3.8263142,4.8765984,5.9268827,6.9732623,7.812709,8.648251,9.487698,10.323239,11.162686,11.127546,11.092407,11.057267,11.022127,10.986988,10.6434,10.303718,9.96013,9.616543,9.276859,8.734148,8.191436,7.648724,7.1060123,6.5633,6.223617,5.8878384,5.548156,5.212377,4.8765984,4.6384296,4.4002614,4.1620927,3.9239242,3.6857557,3.338264,2.9907722,2.6432803,2.2957885,1.9482968,1.9131571,1.8741131,1.8389735,1.7999294,1.7608855,1.6710842,1.5812829,1.4914817,1.4016805,1.3118792,1.4485333,1.5812829,1.717937,1.8506867,1.9873407,1.7882162,1.5929961,1.3938715,1.1986516,0.999527,1.2455044,1.4914817,1.7335546,1.979532,2.2255092,2.4714866,2.7213683,2.9673457,3.213323,3.4632049,3.0415294,2.6159496,2.194274,1.7725986,1.3509232,1.2337911,1.1205635,1.0034313,0.8902037,0.77307165,0.6754616,0.57394713,0.47633708,0.37482262,0.27330816,0.26159495,0.24597734,0.23035973,0.21474212,0.19912452,0.3318742,0.46071947,0.58956474,0.71841,0.8511597,1.0034313,1.1557031,1.3079748,1.4602464,1.6125181,1.7452679,1.8780174,2.0107672,2.1435168,2.2762666,1.9951496,1.7140326,1.43682,1.1557031,0.8745861,0.698888,0.5231899,0.3513962,0.1756981,0.0,1.2689307,2.541766,3.8106966,5.0796275,6.348558,5.6926184,5.036679,4.376835,3.7208953,3.0610514,6.0908675,9.120684,12.154405,15.18422,18.214037,15.21936,12.228588,9.2339115,6.2431393,3.2484627,5.3060827,7.363703,9.421323,11.478943,13.536563,11.650736,9.761005,7.8751793,5.989353,4.0996222,7.043542,9.991365,12.935285,15.879204,18.823124,15.801116,12.779109,9.757101,6.735094,3.7130866,4.322173,4.93126,5.5442514,6.153338,6.7624245,6.602344,6.4422636,6.282183,6.1221027,5.9620223,5.9268827,5.8878384,5.8487945,5.813655,5.774611,5.610626,5.446641,5.278752,5.114767,4.950782,4.985922,5.024966,5.0640097,5.099149,5.138193,5.1889505,5.2436123,5.2943697,5.349031,5.3997884,5.181142,4.958591,4.7399445,4.521298,4.298747,4.3143644,4.3260775,4.337791,4.349504,4.3612175,3.631094,2.8970666,2.1630387,1.4329157,0.698888,0.60908675,0.5192855,0.42948425,0.339683,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.45681506,0.9097257,1.3665408,1.8194515,2.2762666,2.0459068,1.8194515,1.5929961,1.3665408,1.1361811,1.3314011,1.5227169,1.7140326,1.9092526,2.1005683,1.8506867,1.6047094,1.358732,1.1088502,0.8628729,1.0737107,1.2806439,1.4914817,1.7023194,1.9131571,1.8116426,1.7140326,1.6125181,1.5110037,1.4133936,1.3157835,1.2181735,1.1205635,1.0229534,0.92534333,0.8511597,0.77307165,0.698888,0.62470436,0.5505207,0.58566034,0.62079996,0.6559396,0.6910792,0.7262188,0.78868926,0.8550641,0.92143893,0.98390937,1.0502841,0.94486535,0.8394465,0.7340276,0.62860876,0.5231899,0.4958591,0.46852827,0.44119745,0.41386664,0.38653582,0.30844778,0.23426414,0.15617609,0.078088045,0.0,0.6637484,1.3235924,1.9873407,2.6510892,3.310933,3.213323,3.1157131,3.018103,2.9243972,2.8267872,3.7833657,4.743849,5.704332,6.6648145,7.6252975,7.437886,7.250475,7.0630636,6.8756523,6.688241,6.7507114,6.817086,6.883461,6.9459314,7.012306,7.2348576,7.4574084,7.6799593,7.90251,8.125061,7.9766936,7.8283267,7.6838636,7.535496,7.387129,6.969358,6.547683,6.126007,5.708236,5.2865605,4.6735697,4.0605783,3.4514916,2.8385005,2.2255092,2.4324427,2.639376,2.8463092,3.0532427,3.2640803,2.9361105,2.612045,2.2879796,1.9639144,1.6359446,1.6320401,1.6281357,1.6242313,1.6164225,1.6125181,1.4992905,1.3821584,1.2689307,1.1517987,1.038571,1.9209659,2.803361,3.6857557,4.5681505,5.4505453,5.267039,5.083532,4.903929,4.7204223,4.5369153,4.73604,4.93126,5.1303844,5.3256044,5.5247293,5.2358036,4.9468775,4.6540475,4.365122,4.0761957,3.5491016,3.018103,2.4910088,1.9639144,1.43682,0.93705654,0.97610056,1.0190489,1.0580931,1.097137,1.1361811,1.1947471,1.2533131,1.3118792,1.3665408,1.4251068,1.4094892,1.3938715,1.3782539,1.3665408,1.3509232,1.2962615,1.2415999,1.1869383,1.1283722,1.0737107,0.98390937,0.8902037,0.79649806,0.7066968,0.61299115,0.6481308,0.6871748,0.7262188,0.76135844,0.80040246,0.8980125,0.9956226,1.0932326,1.1908426,1.2884527,1.175225,1.0619974,0.94876975,0.8394465,0.7262188,0.7262188,0.7301232,0.7340276,0.7340276,0.737932,0.6520352,0.5661383,0.48414588,0.39824903,0.31235218,0.3318742,0.3513962,0.3709182,0.39434463,0.41386664,0.6832704,0.95267415,1.2220778,1.4914817,1.7608855,1.6320401,1.5031948,1.3743496,1.2415999,1.1127546,0.95657855,0.79649806,0.64032197,0.48414588,0.3240654,0.3474918,0.3709182,0.39434463,0.41386664,0.43729305,0.3631094,0.28892577,0.21083772,0.13665408,0.062470436,0.05466163,0.046852827,0.039044023,0.031235218,0.023426414,0.023426414,0.019522011,0.015617609,0.015617609,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.023426414,0.031235218,0.042948425,0.05075723,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.19522011,0.20302892,0.21083772,0.21864653,0.22645533,0.23426414,0.23816854,0.24597734,0.25378615,0.26159495,0.28111696,0.30063897,0.3240654,0.3435874,0.3631094,0.39434463,0.42557985,0.46071947,0.49195468,0.5231899,0.57785153,0.62860876,0.6832704,0.7340276,0.78868926,0.78868926,0.79259366,0.79649806,0.79649806,0.80040246,0.9058213,1.0151446,1.1205635,1.2298868,1.33921,1.5734742,1.8077383,2.0420024,2.2762666,2.514435,2.2645533,2.018576,1.7686942,1.5227169,1.2767396,1.5695697,1.8663043,2.1591344,2.455869,2.7486992,3.2640803,3.775557,4.2870336,4.7985106,5.3138914,5.1108627,4.9078336,4.704805,4.5017757,4.298747,4.4861584,4.6735697,4.860981,5.0483923,5.2358036,5.3256044,5.4193106,5.5091114,5.5989127,5.688714,5.7121406,5.735567,5.7628975,5.786324,5.813655,5.9268827,6.036206,6.1494336,6.262661,6.375889,6.8405128,7.3051367,7.7697606,8.234385,8.699008,9.0386915,9.37447,9.714153,10.049932,10.38571,9.928895,9.468176,9.007456,8.546737,8.086017,8.00012,7.914223,7.824422,7.7385254,7.648724,7.7814736,7.914223,8.046973,8.179723,8.312472,8.019642,7.726812,7.433982,7.141152,6.8483214,7.1294384,7.406651,7.6838636,7.9610763,8.238289,8.101635,7.9610763,7.824422,7.687768,7.551114,7.7541428,7.9532676,8.156297,8.359325,8.562354,9.171441,9.780528,10.393518,11.002605,11.611692,12.134882,12.658072,13.181262,13.704452,14.223738,13.860628,13.493614,13.130505,12.763491,12.400381,18.221846,24.039404,29.860868,35.67843,41.499893,35.686237,29.876486,24.062832,18.249176,12.439425,10.331048,8.2226715,6.114294,4.0059166,1.901444,1.5695697,1.2415999,0.9097257,0.58175594,0.24988174,0.28892577,0.3318742,0.3709182,0.40996224,0.44900626,0.8667773,1.2845483,1.7023194,2.1200905,2.5378613,2.0302892,1.5227169,1.0151446,0.5075723,0.0,0.0,0.0,0.0,0.0,0.0,0.30844778,0.61689556,0.92143893,1.2298868,1.5383345,1.3431144,1.1517987,0.96048295,0.76916724,0.57394713,0.46462387,0.3553006,0.24597734,0.13665408,0.023426414,0.10541886,0.1835069,0.26549935,0.3435874,0.42557985,0.339683,0.25378615,0.1717937,0.08589685,0.0,3.1469483,6.2938967,9.440845,12.591698,15.738646,13.411622,11.088503,8.761478,6.4383593,4.1113358,3.4593005,2.8072653,2.15523,1.5031948,0.8511597,0.94096094,1.0307622,1.1205635,1.2103647,1.3001659,2.3114061,3.3265507,4.337791,5.349031,6.364176,7.3519893,8.335898,9.323712,10.311526,11.29934,11.232965,11.166591,11.096312,11.029937,10.963562,10.834716,10.705871,10.58093,10.452085,10.323239,9.698535,9.069926,8.441318,7.816613,7.1880045,6.7507114,6.3134184,5.8761253,5.4388323,5.001539,4.7633705,4.5252023,4.2870336,4.0488653,3.8106966,3.4202564,3.0259118,2.6354716,2.241127,1.8506867,1.6867018,1.5266213,1.3626363,1.1986516,1.038571,1.1557031,1.2728351,1.3899672,1.5070993,1.6242313,1.717937,1.8116426,1.901444,1.9951496,2.0888553,1.7843118,1.475864,1.1713207,0.8667773,0.5622339,0.8980125,1.2337911,1.5656652,1.901444,2.2372224,2.5534792,2.87364,3.1898966,3.506153,3.8263142,3.2562714,2.690133,2.1239948,1.5539521,0.9878138,0.92924774,0.8706817,0.8160201,0.75745404,0.698888,0.62470436,0.5505207,0.47633708,0.39824903,0.3240654,0.30454338,0.28502136,0.26549935,0.24597734,0.22645533,0.3279698,0.42948425,0.5309987,0.63641757,0.737932,0.8941081,1.0541886,1.2103647,1.3665408,1.5266213,1.6593709,1.796025,1.9287747,2.0654287,2.1981785,1.8584955,1.5188124,1.1791295,0.8394465,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.63641757,1.2689307,1.9053483,2.541766,3.174279,3.2640803,3.3538816,3.4436827,3.533484,3.6232853,5.5169206,7.406651,9.296382,11.186112,13.075843,10.795672,8.519405,6.2431393,3.9668727,1.6867018,4.084005,6.481308,8.878611,11.275913,13.673217,11.373524,9.073831,6.774138,4.474445,2.174752,6.3602715,10.545791,14.73131,18.916828,23.098444,19.233086,15.363823,11.498465,7.629202,3.7638438,4.318269,4.872694,5.4271193,5.9815445,6.5359693,6.4578815,6.375889,6.297801,6.2158084,6.13772,6.1767645,6.211904,6.250948,6.2860875,6.3251314,6.0791545,5.833177,5.591104,5.3451266,5.099149,5.1108627,5.12648,5.138193,5.1499066,5.1616197,5.044488,4.927356,4.8102236,4.6930914,4.575959,4.388548,4.2050414,4.0215344,3.8341231,3.6506162,3.5998588,3.5491016,3.4983444,3.4514916,3.4007344,2.7916477,2.1786566,1.5695697,0.96048295,0.3513962,0.30454338,0.26159495,0.21474212,0.1717937,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.22645533,0.45681506,0.6832704,0.9097257,1.1361811,1.0307622,0.92143893,0.8160201,0.7066968,0.60127795,0.8277333,1.0541886,1.2806439,1.5110037,1.737459,1.5812829,1.4290112,1.2728351,1.116659,0.96438736,1.2533131,1.5461433,1.8389735,2.1318035,2.4246337,2.135708,1.8506867,1.5617609,1.2767396,0.9878138,0.8823949,0.77697605,0.6715572,0.5661383,0.46071947,0.42557985,0.38653582,0.3513962,0.31235218,0.27330816,0.3318742,0.38653582,0.44119745,0.4958591,0.5505207,0.5583295,0.5661383,0.57394713,0.58175594,0.58566034,0.5231899,0.45681506,0.39434463,0.3279698,0.26159495,0.28111696,0.29673457,0.31625658,0.3318742,0.3513962,0.28111696,0.21083772,0.14055848,0.07027924,0.0,0.62470436,1.2494087,1.8741131,2.4988174,3.1235218,3.1079042,3.0883822,3.0727646,3.0532427,3.0376248,4.01763,4.997635,5.9776397,6.957645,7.9376497,7.7502384,7.562827,7.375416,7.1880045,7.000593,6.969358,6.9381227,6.910792,6.8795567,6.8483214,7.141152,7.433982,7.726812,8.019642,8.312472,7.9337454,7.551114,7.172387,6.79366,6.4110284,6.2040954,5.9932575,5.7824197,5.571582,5.3607445,4.8492675,4.337791,3.8263142,3.310933,2.7994564,2.9868677,3.1703746,3.3538816,3.541293,3.7247996,3.4007344,3.076669,2.7486992,2.4246337,2.1005683,2.096664,2.096664,2.0927596,2.0888553,2.0888553,1.9443923,1.796025,1.6515622,1.5070993,1.3626363,2.4207294,3.4827268,4.5408196,5.602817,6.66091,6.3915067,6.1181984,5.84489,5.571582,5.298274,5.481781,5.661383,5.840986,6.0205884,6.2001905,5.8683167,5.5364423,5.2006636,4.8687897,4.5369153,3.8809757,3.2211318,2.5651922,1.9092526,1.2494087,1.0619974,1.0619974,1.0619974,1.0619974,1.0619974,1.0619974,0.9878138,0.9136301,0.8394465,0.76135844,0.6871748,0.6481308,0.61299115,0.57394713,0.5388075,0.4997635,0.47633708,0.44900626,0.42557985,0.39824903,0.37482262,0.3513962,0.3240654,0.30063897,0.27330816,0.24988174,0.3357786,0.42557985,0.5114767,0.60127795,0.6871748,0.8238289,0.96438736,1.1010414,1.2376955,1.3743496,1.2494087,1.1244678,0.999527,0.8745861,0.74964523,0.74964523,0.74964523,0.74964523,0.74964523,0.74964523,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.18741131,0.24988174,0.31235218,0.37482262,0.43729305,0.698888,0.96438736,1.2259823,1.4875772,1.7491722,1.6632754,1.5734742,1.4875772,1.4016805,1.3118792,1.1127546,0.9136301,0.7106012,0.5114767,0.31235218,0.3357786,0.3631094,0.38653582,0.41386664,0.43729305,0.3631094,0.28892577,0.21083772,0.13665408,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,0.26159495,0.27330816,0.28892577,0.30063897,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.3357786,0.3631094,0.38653582,0.41386664,0.43729305,0.5114767,0.58566034,0.6637484,0.737932,0.81211567,1.0893283,1.3626363,1.6359446,1.9131571,2.1864653,1.9482968,1.7140326,1.475864,1.2376955,0.999527,1.261122,1.5266213,1.7882162,2.0498111,2.3114061,2.8892577,3.4632049,4.037152,4.6110992,5.1889505,4.939069,4.689187,4.4393053,4.1894236,3.9356375,4.0996222,4.263607,4.423688,4.5876727,4.7516575,4.7243266,4.7009,4.6735697,4.650143,4.6267166,4.786797,4.950782,5.1108627,5.2748475,5.4388323,5.575486,5.7121406,5.8487945,5.989353,6.126007,6.7116675,7.3012323,7.8868923,8.476458,9.062118,9.526741,9.987461,10.44818,10.912805,11.373524,10.838621,10.299813,9.761005,9.226103,8.687295,8.6131115,8.538928,8.460839,8.386656,8.312472,8.413987,8.511597,8.6131115,8.710721,8.812236,8.449126,8.086017,7.726812,7.363703,7.000593,7.2739015,7.551114,7.824422,8.101635,8.374943,8.187531,8.00012,7.812709,7.6252975,7.437886,7.7619514,8.086017,8.413987,8.738052,9.062118,9.636065,10.213917,10.787864,11.361811,11.935758,12.412095,12.888432,13.360865,13.837202,14.313539,13.462379,12.611219,11.763964,10.912805,10.061645,16.449247,22.83685,29.224451,35.612053,41.999657,35.576912,29.150267,22.723621,16.300879,9.874233,8.062591,6.250948,4.4393053,2.6237583,0.81211567,0.7106012,0.61299115,0.5114767,0.41386664,0.31235218,0.3631094,0.41386664,0.46071947,0.5114767,0.5622339,1.0502841,1.5383345,2.0263848,2.514435,2.998581,2.4012074,1.7999294,1.1986516,0.60127795,0.0,0.0,0.0,0.0,0.0,0.0,0.28892577,0.57394713,0.8628729,1.1517987,1.43682,1.175225,0.9136301,0.6481308,0.38653582,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.513962,7.0240197,10.537982,14.051944,17.562002,14.848442,12.138786,9.425227,6.7116675,3.998108,3.2250361,2.4519646,1.6749885,0.9019169,0.12494087,0.27330816,0.42557985,0.57394713,0.7262188,0.8745861,1.8506867,2.8267872,3.7989833,4.775084,5.7511845,6.8873653,8.023546,9.163632,10.299813,11.435994,11.338385,11.23687,11.139259,11.037745,10.936231,11.0260315,11.111929,11.20173,11.287627,11.373524,10.662923,9.948417,9.237816,8.52331,7.812709,7.2739015,6.7389984,6.2001905,5.661383,5.12648,4.8883114,4.650143,4.4119744,4.173806,3.9356375,3.4983444,3.0610514,2.6237583,2.1864653,1.7491722,1.4641509,1.175225,0.8862993,0.60127795,0.31235218,0.63641757,0.96438736,1.2884527,1.6125181,1.9365835,1.9873407,2.0380979,2.0888553,2.135708,2.1864653,1.7765031,1.3626363,0.94876975,0.5388075,0.12494087,0.5505207,0.97610056,1.4016805,1.8233559,2.2489357,2.639376,3.0259118,3.4124475,3.7989833,4.1894236,3.474918,2.7643168,2.0498111,1.33921,0.62470436,0.62470436,0.62470436,0.62470436,0.62470436,0.62470436,0.57394713,0.5231899,0.47633708,0.42557985,0.37482262,0.3513962,0.3240654,0.30063897,0.27330816,0.24988174,0.3240654,0.39824903,0.47633708,0.5505207,0.62470436,0.78868926,0.94876975,1.1127546,1.2767396,1.43682,1.5734742,1.7140326,1.8506867,1.9873407,2.1239948,1.7257458,1.3235924,0.92534333,0.5231899,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.8394465,1.6749885,2.514435,3.349977,4.1894236,4.939069,5.688714,6.4383593,7.1880045,7.9376497,6.375889,4.814128,3.2484627,1.6867018,0.12494087,2.8619268,5.5989127,8.335898,11.076789,13.813775,11.100216,8.386656,5.6730967,2.9634414,0.24988174,5.677001,11.100216,16.52343,21.95055,27.373764,22.66115,17.948538,13.235924,8.52331,3.8106966,4.3143644,4.814128,5.3138914,5.813655,6.3134184,6.3134184,6.3134184,6.3134184,6.3134184,6.3134184,6.426646,6.5359693,6.649197,6.7624245,6.8756523,6.551587,6.223617,5.899552,5.575486,5.251421,5.2358036,5.22409,5.212377,5.2006636,5.1889505,4.900025,4.6110992,4.3260775,4.037152,3.7482262,3.5998588,3.4514916,3.2992198,3.1508527,2.998581,2.8892577,2.77603,2.6628022,2.5495746,2.436347,1.9482968,1.4641509,0.97610056,0.48805028,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.3240654,0.58566034,0.8511597,1.1127546,1.3743496,1.3118792,1.2494087,1.1869383,1.1244678,1.0619974,1.43682,1.8116426,2.1864653,2.5612879,2.9361105,2.463678,1.9873407,1.5110037,1.038571,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.3240654,0.27330816,0.22645533,0.1756981,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.58566034,1.175225,1.7608855,2.35045,2.9361105,2.998581,3.0610514,3.1235218,3.1859922,3.2484627,4.251894,5.251421,6.250948,7.250475,8.250002,8.062591,7.8751793,7.687768,7.5003567,7.3129454,7.1880045,7.0630636,6.9381227,6.813182,6.688241,7.0513506,7.4105554,7.773665,8.136774,8.499884,7.8868923,7.2739015,6.66091,6.0518236,5.4388323,5.4388323,5.4388323,5.4388323,5.4388323,5.4388323,5.024966,4.6110992,4.2011366,3.78727,3.3734035,3.5373883,3.7013733,3.8614538,4.025439,4.1894236,3.8614538,3.5373883,3.213323,2.8892577,2.5612879,2.5612879,2.5612879,2.5612879,2.5612879,2.5612879,2.3855898,2.2137961,2.0380979,1.8623998,1.6867018,2.9243972,4.1620927,5.3997884,6.6374836,7.8751793,7.5120697,7.1489606,6.785851,6.426646,6.0635366,6.223617,6.387602,6.551587,6.7116675,6.8756523,6.5008297,6.126007,5.7511845,5.376362,5.001539,4.21285,3.4241607,2.639376,1.8506867,1.0619974,1.6242313,1.5188124,1.4094892,1.3040704,1.1947471,1.0893283,1.0580931,1.0268579,0.9956226,0.96829176,0.93705654,0.8706817,0.80821127,0.7418364,0.679366,0.61299115,0.59737355,0.58175594,0.5661383,0.5544251,0.5388075,0.5192855,0.4958591,0.47633708,0.45681506,0.43729305,0.5622339,0.6871748,0.81211567,0.93705654,1.0619974,1.1322767,1.2025559,1.2728351,1.3431144,1.4133936,1.2572175,1.1010414,0.94876975,0.79259366,0.63641757,0.62860876,0.62079996,0.61689556,0.60908675,0.60127795,0.5075723,0.41386664,0.3240654,0.23035973,0.13665408,0.23426414,0.3318742,0.42948425,0.5270943,0.62470436,0.78478485,0.94486535,1.1049459,1.2650263,1.4251068,1.3509232,1.2767396,1.1986516,1.1244678,1.0502841,0.8902037,0.7301232,0.5700427,0.40996224,0.24988174,0.29673457,0.339683,0.38653582,0.42948425,0.47633708,0.39044023,0.30454338,0.21864653,0.13665408,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.042948425,0.03513962,0.027330816,0.019522011,0.011713207,0.027330816,0.042948425,0.058566034,0.07418364,0.08589685,0.10932326,0.13274968,0.15617609,0.1756981,0.19912452,0.20302892,0.20693332,0.20693332,0.21083772,0.21083772,0.20693332,0.19912452,0.19131571,0.1835069,0.1756981,0.1835069,0.19522011,0.20693332,0.21474212,0.22645533,0.23816854,0.24988174,0.26159495,0.27330816,0.28892577,0.28892577,0.29283017,0.29673457,0.29673457,0.30063897,0.3240654,0.3435874,0.3670138,0.39044023,0.41386664,0.48024148,0.5466163,0.61689556,0.6832704,0.74964523,0.98390937,1.2142692,1.4485333,1.678893,1.9131571,1.7413634,1.5656652,1.3938715,1.2220778,1.0502841,1.2533131,1.4602464,1.6632754,1.8702087,2.0732377,2.5612879,3.049338,3.5373883,4.025439,4.513489,4.3455997,4.181615,4.01763,3.853645,3.6857557,3.8419318,3.998108,4.154284,4.3065557,4.462732,4.513489,4.5681505,4.618908,4.6735697,4.7243266,4.814128,4.900025,4.985922,5.0757227,5.1616197,5.2553253,5.349031,5.4388323,5.532538,5.6262436,6.2197127,6.813182,7.4105554,8.0040245,8.601398,8.956698,9.308095,9.663396,10.018696,10.373997,9.971844,9.56969,9.167537,8.765383,8.36323,8.331994,8.300759,8.273428,8.242193,8.210958,8.253906,8.296855,8.339804,8.382751,8.4257,8.289046,8.148487,8.011833,7.8751793,7.7385254,7.9766936,8.218767,8.456935,8.699008,8.937177,8.804427,8.671678,8.538928,8.406178,8.273428,8.644346,9.0152645,9.386183,9.753197,10.124115,10.612165,11.100216,11.588266,12.076316,12.564366,12.939189,13.314012,13.688834,14.063657,14.438479,13.946525,13.450665,12.958711,12.466757,11.974802,17.999294,24.019882,30.044374,36.064964,42.085552,35.303604,28.521658,21.739712,14.957765,8.175818,7.043542,5.9151692,4.786797,3.6545205,2.5261483,2.3035975,2.0810463,1.8584955,1.6359446,1.4133936,1.2181735,1.0268579,0.8355421,0.6442264,0.44900626,0.8433509,1.2337911,1.6281357,2.018576,2.4129205,2.1200905,1.8272603,1.53443,1.2415999,0.94876975,0.8238289,0.698888,0.57394713,0.44900626,0.3240654,0.48805028,0.6559396,0.8199245,0.98390937,1.1517987,0.94096094,0.7301232,0.5192855,0.30844778,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,3.2055142,6.3134184,9.421323,12.529227,15.637131,13.200784,10.768341,8.331994,5.8956475,3.4632049,2.8189783,2.1786566,1.53443,0.8941081,0.24988174,0.5231899,0.80040246,1.0737107,1.3509232,1.6242313,2.7252727,3.8263142,4.9234514,6.0244927,7.125534,7.812709,8.499884,9.187058,9.874233,10.561408,10.545791,10.534078,10.518459,10.502842,10.487225,10.471607,10.455989,10.444276,10.4286585,10.413041,9.917182,9.421323,8.929368,8.433509,7.9376497,7.551114,7.168483,6.7819467,6.3993154,6.012779,5.5989127,5.1889505,4.775084,4.3612175,3.951255,3.5725281,3.193801,2.8189783,2.4402514,2.0615244,1.8038338,1.5461433,1.2884527,1.0307622,0.77307165,1.0268579,1.2767396,1.5266213,1.7765031,2.0263848,2.0224805,2.018576,2.018576,2.0146716,2.0107672,1.6749885,1.33921,0.999527,0.6637484,0.3240654,0.63641757,0.94486535,1.2533131,1.5656652,1.8741131,2.2177005,2.5612879,2.900971,3.2445583,3.5881457,3.0024853,2.416825,1.8311646,1.2494087,0.6637484,0.6481308,0.63251317,0.61689556,0.60127795,0.58566034,0.5661383,0.5466163,0.5270943,0.5075723,0.48805028,0.44119745,0.39824903,0.3513962,0.30844778,0.26159495,0.3513962,0.44119745,0.5309987,0.62079996,0.7106012,0.8433509,0.97610056,1.1088502,1.2415999,1.3743496,1.5890918,1.7999294,2.0107672,2.2255092,2.436347,2.069333,1.698415,1.3274968,0.95657855,0.58566034,0.46852827,0.3513962,0.23426414,0.11713207,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.698888,1.3626363,2.0263848,2.6862288,3.349977,3.951255,4.548629,5.1499066,5.7511845,6.348558,5.099149,3.8497405,2.6003318,1.3509232,0.10151446,2.494913,4.8883114,7.2856145,9.679013,12.076316,9.8195715,7.5667315,5.309987,3.0532427,0.80040246,6.0596323,11.318862,16.581997,21.841227,27.100456,22.692387,18.284315,13.8762455,9.468176,5.0640097,5.2358036,5.4115014,5.5871997,5.7628975,5.938596,6.086963,6.239235,6.387602,6.5359693,6.688241,6.617962,6.547683,6.477403,6.407124,6.336845,6.1611466,5.9815445,5.805846,5.6262436,5.4505453,5.407597,5.364649,5.3217,5.278752,5.2358036,5.0601053,4.884407,4.704805,4.5291066,4.349504,4.1581883,3.9668727,3.7716527,3.5803368,3.3890212,3.2211318,3.0532427,2.8853533,2.717464,2.5495746,2.0380979,1.5305257,1.0190489,0.5114767,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.26159495,0.46852827,0.679366,0.8902037,1.1010414,1.0502841,0.999527,0.94876975,0.9019169,0.8511597,1.1517987,1.4485333,1.7491722,2.0498111,2.35045,1.9717231,1.5890918,1.2103647,0.8316377,0.44900626,0.359205,0.26940376,0.1796025,0.08980125,0.0,0.0,0.0,0.0,0.0,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.27330816,0.23426414,0.19131571,0.15227169,0.113227665,0.093705654,0.078088045,0.058566034,0.042948425,0.023426414,0.07418364,0.12103647,0.1678893,0.21474212,0.26159495,0.21083772,0.15617609,0.10541886,0.05075723,0.0,0.4958591,0.9956226,1.4914817,1.9912452,2.4871042,2.612045,2.736986,2.8619268,2.9868677,3.1118085,3.9824903,4.853172,5.7238536,6.590631,7.461313,7.4144597,7.367607,7.320754,7.2739015,7.223144,7.039637,6.8561306,6.6687193,6.4852123,6.3017054,6.688241,7.0786815,7.4691215,7.859562,8.250002,7.70729,7.164578,6.621866,6.0791545,5.5364423,5.579391,5.6223392,5.6652875,5.708236,5.7511845,5.4388323,5.1303844,4.8219366,4.5095844,4.2011366,4.40807,4.6150036,4.8219366,5.02887,5.2358036,4.892216,4.548629,4.2011366,3.8575494,3.513962,3.6623292,3.8106966,3.9629683,4.1113358,4.263607,4.0059166,3.7521305,3.4983444,3.240654,2.9868677,4.0020123,5.017157,6.0323014,7.0474463,8.062591,7.715099,7.367607,7.0201154,6.6726236,6.3251314,6.3056097,6.2860875,6.266566,6.2431393,6.223617,5.989353,5.755089,5.520825,5.2865605,5.0483923,4.318269,3.5842414,2.854118,2.1200905,1.3860629,2.1864653,1.9717231,1.756981,1.542239,1.3274968,1.1127546,1.1283722,1.1439898,1.1557031,1.1713207,1.1869383,1.0932326,1.0034313,0.9097257,0.8160201,0.7262188,0.71841,0.7145056,0.7106012,0.7066968,0.698888,0.6832704,0.6715572,0.6559396,0.64032197,0.62470436,0.78868926,0.94876975,1.1127546,1.2767396,1.43682,1.4407244,1.4407244,1.4446288,1.4485333,1.4485333,1.2650263,1.0815194,0.8941081,0.7106012,0.5231899,0.5114767,0.4958591,0.48024148,0.46462387,0.44900626,0.39044023,0.3318742,0.26940376,0.21083772,0.14836729,0.28111696,0.41386664,0.5466163,0.679366,0.81211567,0.8706817,0.92924774,0.98390937,1.0424755,1.1010414,1.038571,0.97610056,0.9136301,0.8511597,0.78868926,0.6676528,0.5466163,0.42557985,0.30844778,0.18741131,0.25378615,0.31625658,0.38263142,0.44900626,0.5114767,0.41777104,0.3240654,0.22645533,0.13274968,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.08589685,0.07027924,0.05466163,0.039044023,0.023426414,0.042948425,0.058566034,0.078088045,0.093705654,0.113227665,0.13274968,0.15227169,0.1717937,0.19131571,0.21083772,0.21864653,0.22255093,0.22645533,0.23426414,0.23816854,0.22255093,0.20693332,0.19131571,0.1756981,0.1639849,0.1717937,0.1756981,0.1835069,0.19131571,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,0.26159495,0.26940376,0.27330816,0.27721256,0.28111696,0.28892577,0.30844778,0.3279698,0.3474918,0.3670138,0.38653582,0.44900626,0.5075723,0.5661383,0.62860876,0.6871748,0.8784905,1.0659018,1.2572175,1.4485333,1.6359446,1.5305257,1.4212024,1.3157835,1.2064602,1.1010414,1.2494087,1.3938715,1.542239,1.6906061,1.8389735,2.2372224,2.639376,3.0376248,3.435874,3.8380275,3.7560349,3.677947,3.5959544,3.5178664,3.435874,3.5842414,3.7326086,3.8809757,4.029343,4.173806,4.3065557,4.435401,4.564246,4.6930914,4.825841,4.8375545,4.8492675,4.860981,4.8765984,4.8883114,4.9351645,4.9820175,5.02887,5.0757227,5.12648,5.727758,6.329036,6.9342184,7.535496,8.136774,8.386656,8.632633,8.878611,9.128492,9.37447,9.108971,8.839567,8.574067,8.304664,8.039165,8.050878,8.066495,8.082112,8.097731,8.113348,8.097731,8.082112,8.066495,8.050878,8.039165,8.125061,8.210958,8.300759,8.386656,8.476458,8.679486,8.886419,9.089449,9.296382,9.499411,9.421323,9.343235,9.269051,9.190963,9.112875,9.526741,9.940608,10.358379,10.772245,11.186112,11.588266,11.986515,12.388668,12.786918,13.189071,13.462379,13.735687,14.012899,14.286208,14.56342,14.426766,14.294017,14.157363,14.020708,13.887959,19.545437,25.202917,30.860395,36.517876,42.175354,35.034203,27.896954,20.755802,13.614651,6.473499,6.028397,5.579391,5.134289,4.6852827,4.2362766,3.892689,3.5491016,3.2016098,2.8580225,2.514435,2.077142,1.6437533,1.2064602,0.77307165,0.3357786,0.63641757,0.93315214,1.2298868,1.5266213,1.8233559,1.8389735,1.8545911,1.8702087,1.8858263,1.901444,1.6515622,1.4016805,1.1517987,0.9019169,0.6481308,0.6910792,0.7340276,0.77697605,0.8199245,0.8628729,0.7066968,0.5466163,0.39044023,0.23426414,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,2.900971,5.606722,8.308568,11.010414,13.712261,11.553126,9.397896,7.238762,5.083532,2.9243972,2.416825,1.9053483,1.3938715,0.8862993,0.37482262,0.77697605,1.175225,1.5734742,1.9756275,2.3738766,3.5998588,4.825841,6.0518236,7.2739015,8.499884,8.738052,8.976221,9.21439,9.448653,9.686822,9.757101,9.82738,9.897659,9.967939,10.0382185,9.921086,9.803954,9.686822,9.565785,9.448653,9.171441,8.894228,8.617016,8.339804,8.062591,7.8283267,7.5979667,7.363703,7.1333427,6.899079,6.3134184,5.7238536,5.138193,4.548629,3.9629683,3.6467118,3.3265507,3.0102942,2.6940374,2.3738766,2.1474214,1.9209659,1.6906061,1.4641509,1.2376955,1.4133936,1.5890918,1.7608855,1.9365835,2.1122816,2.05762,2.0029583,1.9482968,1.893635,1.8389735,1.5734742,1.3118792,1.0502841,0.78868926,0.5231899,0.71841,0.9136301,1.1088502,1.3040704,1.4992905,1.796025,2.096664,2.3933985,2.690133,2.9868677,2.5300527,2.0732377,1.6164225,1.1557031,0.698888,0.6715572,0.64032197,0.60908675,0.58175594,0.5505207,0.5583295,0.5700427,0.58175594,0.58956474,0.60127795,0.5349031,0.46852827,0.40605783,0.339683,0.27330816,0.37872702,0.48414588,0.58956474,0.6949836,0.80040246,0.9019169,1.0034313,1.1088502,1.2103647,1.3118792,1.6008049,1.8858263,2.174752,2.463678,2.7486992,2.4090161,2.069333,1.7296503,1.3899672,1.0502841,0.8394465,0.62860876,0.42167544,0.21083772,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.5622339,1.0502841,1.5383345,2.0263848,2.514435,2.9634414,3.4124475,3.8614538,4.3143644,4.7633705,3.8263142,2.8892577,1.9482968,1.0112402,0.07418364,2.1278992,4.181615,6.2314262,8.285142,10.338858,8.538928,6.7429028,4.9468775,3.1469483,1.3509232,6.446168,11.541413,16.636658,21.731903,26.823244,22.723621,18.620094,14.516567,10.413041,6.3134184,6.1611466,6.012779,5.8644123,5.7121406,5.563773,5.8644123,6.1611466,6.461786,6.7624245,7.0630636,6.8092775,6.559396,6.3056097,6.0518236,5.801942,5.7707067,5.7394714,5.708236,5.6809053,5.64967,5.579391,5.505207,5.4310236,5.3607445,5.2865605,5.2201858,5.153811,5.083532,5.017157,4.950782,4.716518,4.478349,4.2440853,4.009821,3.775557,3.5530062,3.330455,3.1079042,2.8853533,2.6628022,2.1318035,1.5969005,1.0659018,0.5309987,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.19522011,0.3513962,0.5114767,0.6676528,0.8238289,0.78868926,0.74964523,0.7106012,0.6754616,0.63641757,0.8628729,1.0893283,1.3118792,1.5383345,1.7608855,1.475864,1.1908426,0.9058213,0.62079996,0.3357786,0.26940376,0.20302892,0.13665408,0.06637484,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.21864653,0.19131571,0.16008049,0.12884527,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.08199245,0.113227665,0.14836729,0.1796025,0.21083772,0.1717937,0.12884527,0.08589685,0.042948425,0.0,0.40605783,0.8160201,1.2220778,1.6281357,2.0380979,2.2255092,2.4129205,2.6003318,2.787743,2.9751544,3.716991,4.454923,5.196759,5.9346914,6.676528,6.7663293,6.860035,6.9537406,7.043542,7.137247,6.89127,6.649197,6.4032197,6.1572423,5.911265,6.329036,6.746807,7.164578,7.5823493,8.00012,7.5276875,7.055255,6.5828223,6.1103897,5.6379566,5.7238536,5.805846,5.891743,5.9776397,6.0635366,5.8566036,5.645766,5.4388323,5.2318993,5.024966,5.278752,5.5286336,5.7824197,6.036206,6.2860875,5.9229784,5.5559645,5.192855,4.825841,4.462732,4.7633705,5.0640097,5.3607445,5.661383,5.9620223,5.6262436,5.2943697,4.958591,4.6228123,4.2870336,5.0796275,5.872221,6.6648145,7.4574084,8.250002,7.918128,7.5862536,7.2543793,6.918601,6.5867267,6.3836975,6.180669,5.9815445,5.7785153,5.575486,5.481781,5.3841705,5.290465,5.196759,5.099149,4.423688,3.7443218,3.06886,2.3894942,1.7140326,2.7486992,2.4285383,2.1044729,1.7843118,1.4602464,1.1361811,1.1986516,1.2572175,1.3157835,1.3782539,1.43682,1.3157835,1.1986516,1.077615,0.95657855,0.8394465,0.8433509,0.8472553,0.8511597,0.8589685,0.8628729,0.8511597,0.8433509,0.8316377,0.8238289,0.81211567,1.0112402,1.2142692,1.4133936,1.6125181,1.8116426,1.7491722,1.6827974,1.6164225,1.5539521,1.4875772,1.2728351,1.0580931,0.8433509,0.62860876,0.41386664,0.39044023,0.3670138,0.3435874,0.3240654,0.30063897,0.27330816,0.24597734,0.21864653,0.19131571,0.1639849,0.3318742,0.4958591,0.6637484,0.8316377,0.999527,0.95657855,0.9097257,0.8667773,0.8199245,0.77307165,0.7262188,0.6754616,0.62470436,0.57394713,0.5231899,0.44510186,0.3631094,0.28502136,0.20693332,0.12494087,0.21083772,0.29673457,0.37872702,0.46462387,0.5505207,0.44510186,0.339683,0.23426414,0.12884527,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.12884527,0.10541886,0.08199245,0.058566034,0.039044023,0.058566034,0.078088045,0.09761006,0.11713207,0.13665408,0.15617609,0.1717937,0.19131571,0.20693332,0.22645533,0.23426414,0.23816854,0.24597734,0.25378615,0.26159495,0.23816854,0.21864653,0.19522011,0.1717937,0.14836729,0.15617609,0.16008049,0.1639849,0.1717937,0.1756981,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24597734,0.25378615,0.26159495,0.26940376,0.27330816,0.29283017,0.30844778,0.3279698,0.3435874,0.3631094,0.41386664,0.46852827,0.5192855,0.57394713,0.62470436,0.77307165,0.92143893,1.0659018,1.2142692,1.3626363,1.319688,1.2767396,1.2337911,1.1908426,1.1517987,1.2415999,1.3314011,1.4212024,1.5110037,1.6008049,1.9131571,2.2255092,2.5378613,2.8502135,3.1625657,3.1664703,3.174279,3.1781836,3.182088,3.1859922,3.3265507,3.4671092,3.6076677,3.7482262,3.8887846,4.095718,4.3026514,4.5095844,4.716518,4.9234514,4.860981,4.7985106,4.73604,4.6735697,4.6110992,4.6150036,4.618908,4.618908,4.6228123,4.6267166,5.2358036,5.84489,6.453977,7.0630636,7.676055,7.816613,7.9532676,8.093826,8.234385,8.374943,8.242193,8.109444,7.9766936,7.843944,7.7111945,7.773665,7.832231,7.890797,7.9532676,8.011833,7.941554,7.8673706,7.793187,7.7229075,7.648724,7.9610763,8.273428,8.58578,8.898132,9.21439,9.382278,9.554072,9.721962,9.893755,10.061645,10.0382185,10.018696,9.99527,9.971844,9.948417,10.409137,10.869856,11.330575,11.791295,12.24811,12.564366,12.8767185,13.189071,13.501423,13.813775,13.985569,14.161267,14.336966,14.512663,14.688361,14.9109125,15.133463,15.356014,15.578565,15.801116,21.091581,26.38595,31.676416,36.970783,42.26125,34.764797,27.268345,19.767988,12.271536,4.775084,5.009348,5.2436123,5.481781,5.716045,5.950309,5.481781,5.0132523,4.548629,4.0801005,3.611572,2.9361105,2.2567444,1.5812829,0.9019169,0.22645533,0.42557985,0.62860876,0.8316377,1.0346665,1.2376955,1.5617609,1.8819219,2.2059872,2.5261483,2.8502135,2.475391,2.1005683,1.7257458,1.3509232,0.97610056,0.8941081,0.8160201,0.7340276,0.6559396,0.57394713,0.46852827,0.3631094,0.26159495,0.15617609,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,2.5964274,4.8961205,7.191909,9.491602,11.787391,9.909373,8.027451,6.1455293,4.267512,2.3855898,2.0107672,1.6320401,1.2533131,0.8784905,0.4997635,1.0268579,1.5500476,2.0732377,2.6003318,3.1235218,4.474445,5.825368,7.1762915,8.52331,9.874233,9.663396,9.448653,9.237816,9.023073,8.812236,8.968412,9.120684,9.276859,9.433036,9.589212,9.366661,9.148014,8.929368,8.706817,8.488171,8.4257,8.367134,8.308568,8.246098,8.187531,8.109444,8.027451,7.9493628,7.8673706,7.7892823,7.0240197,6.262661,5.5013027,4.73604,3.9746814,3.716991,3.4593005,3.2016098,2.9439192,2.6862288,2.4910088,2.2918842,2.096664,1.8975395,1.698415,1.7999294,1.901444,1.999054,2.1005683,2.1981785,2.0927596,1.9834363,1.8780174,1.7686942,1.6632754,1.475864,1.2884527,1.1010414,0.9136301,0.7262188,0.80430686,0.8862993,0.96438736,1.0463798,1.1244678,1.3782539,1.6281357,1.8819219,2.135708,2.3855898,2.05762,1.7257458,1.397776,1.0659018,0.737932,0.6910792,0.6481308,0.60127795,0.5583295,0.5114767,0.5544251,0.59346914,0.63251317,0.6715572,0.7106012,0.62860876,0.5427119,0.45681506,0.3709182,0.28892577,0.40605783,0.5270943,0.6481308,0.76916724,0.8862993,0.96048295,1.0307622,1.1049459,1.1791295,1.2494087,1.6125181,1.9756275,2.338737,2.7018464,3.0610514,2.7526035,2.4441557,2.1318035,1.8233559,1.5110037,1.2103647,0.9058213,0.60518235,0.30063897,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.42557985,0.737932,1.0502841,1.3626363,1.6749885,1.9756275,2.2762666,2.5769055,2.87364,3.174279,2.5495746,1.9248703,1.3001659,0.6754616,0.05075723,1.7608855,3.4710135,5.181142,6.89127,8.601398,7.2582836,5.919074,4.579864,3.240654,1.901444,6.8287997,11.760059,16.69132,21.618675,26.549934,22.750952,18.955873,15.15689,11.361811,7.562827,7.08649,6.6140575,6.13772,5.661383,5.1889505,5.6379566,6.086963,6.5359693,6.98888,7.437886,7.000593,6.5672045,6.133816,5.6965227,5.263134,5.380266,5.4973984,5.6145306,5.7316628,5.8487945,5.74728,5.645766,5.5442514,5.4388323,5.337318,5.380266,5.423215,5.466163,5.5091114,5.548156,5.270943,4.9937305,4.716518,4.4393053,4.1620927,3.8848803,3.6076677,3.330455,3.0532427,2.77603,2.2216048,1.6632754,1.1088502,0.5544251,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.12884527,0.23426414,0.339683,0.44510186,0.5505207,0.5231899,0.4997635,0.47633708,0.44900626,0.42557985,0.57394713,0.7262188,0.8745861,1.0268579,1.175225,0.98390937,0.79649806,0.60518235,0.41386664,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.1678893,0.14836729,0.12884527,0.10932326,0.08589685,0.08589685,0.08199245,0.078088045,0.078088045,0.07418364,0.093705654,0.10932326,0.12884527,0.14446288,0.1639849,0.12884527,0.09761006,0.06637484,0.031235218,0.0,0.31625658,0.63641757,0.95267415,1.2689307,1.5890918,1.8389735,2.0888553,2.338737,2.5886188,2.8385005,3.4475873,4.056674,4.6657605,5.278752,5.8878384,6.1181984,6.3524623,6.5867267,6.817086,7.0513506,6.746807,6.4383593,6.133816,5.8292727,5.5247293,5.969831,6.4149327,6.860035,7.3051367,7.7502384,7.348085,6.9459314,6.5437784,6.141625,5.735567,5.8644123,5.9932575,6.1181984,6.2470436,6.375889,6.27047,6.165051,6.0596323,5.9542136,5.8487945,6.1494336,6.446168,6.7429028,7.039637,7.336372,6.9537406,6.5672045,6.180669,5.7980375,5.4115014,5.8644123,6.3134184,6.7624245,7.211431,7.6643414,7.2465706,6.832704,6.4188375,6.001066,5.5871997,6.1572423,6.727285,7.297328,7.8673706,8.437413,8.121157,7.800996,7.4847393,7.168483,6.8483214,6.46569,6.0791545,5.6965227,5.309987,4.9234514,4.970304,5.0132523,5.0601053,5.1030536,5.1499066,4.5291066,3.9044023,3.2836022,2.6588979,2.0380979,3.310933,2.8814487,2.4519646,2.0224805,1.5929961,1.1635119,1.2689307,1.3743496,1.475864,1.5812829,1.6867018,1.5383345,1.3938715,1.2455044,1.097137,0.94876975,0.96438736,0.98000497,0.9956226,1.0112402,1.0268579,1.0190489,1.0151446,1.0112402,1.0034313,0.999527,1.2376955,1.475864,1.7140326,1.9482968,2.1864653,2.0537157,1.9209659,1.7882162,1.6593709,1.5266213,1.2806439,1.0346665,0.78868926,0.5466163,0.30063897,0.26940376,0.23816854,0.21083772,0.1796025,0.14836729,0.15617609,0.16008049,0.1639849,0.1717937,0.1756981,0.37872702,0.58175594,0.78088045,0.98390937,1.1869383,1.038571,0.8941081,0.74574083,0.59737355,0.44900626,0.41386664,0.37482262,0.3357786,0.30063897,0.26159495,0.22255093,0.1835069,0.14055848,0.10151446,0.062470436,0.1678893,0.27330816,0.37872702,0.48414588,0.58566034,0.47243267,0.359205,0.24207294,0.12884527,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.1717937,0.14055848,0.10932326,0.078088045,0.05075723,0.07418364,0.093705654,0.11713207,0.14055848,0.1639849,0.1756981,0.19131571,0.20693332,0.22255093,0.23816854,0.24597734,0.25769055,0.26940376,0.27721256,0.28892577,0.25769055,0.22645533,0.19912452,0.1678893,0.13665408,0.14055848,0.14055848,0.14446288,0.14836729,0.14836729,0.1639849,0.1756981,0.18741131,0.19912452,0.21083772,0.22255093,0.23426414,0.24207294,0.25378615,0.26159495,0.27721256,0.29283017,0.30844778,0.3240654,0.3357786,0.38263142,0.42557985,0.47243267,0.5192855,0.5622339,0.6676528,0.77307165,0.8784905,0.98390937,1.0893283,1.1088502,1.1322767,1.1557031,1.1791295,1.1986516,1.2337911,1.2650263,1.2962615,1.3314011,1.3626363,1.5890918,1.8116426,2.0380979,2.260649,2.4871042,2.5769055,2.6667068,2.7565079,2.8463092,2.9361105,3.06886,3.2016098,3.3343596,3.4671092,3.5998588,3.8848803,4.169902,4.454923,4.7399445,5.024966,4.8883114,4.7516575,4.6110992,4.474445,4.337791,4.2948427,4.251894,4.2089458,4.165997,4.126953,4.743849,5.3607445,5.9776397,6.5945354,7.211431,7.2465706,7.277806,7.309041,7.3441806,7.375416,7.37932,7.37932,7.3832245,7.3832245,7.387129,7.492548,7.5979667,7.703386,7.8088045,7.914223,7.7814736,7.6526284,7.523783,7.3910336,7.262188,7.800996,8.335898,8.874706,9.413514,9.948417,10.085071,10.221725,10.354475,10.491129,10.6238785,10.6590185,10.690253,10.721489,10.756628,10.787864,11.291532,11.799104,12.302772,12.806439,13.314012,13.536563,13.763018,13.985569,14.212025,14.438479,14.512663,14.586847,14.661031,14.739119,14.813302,15.391153,15.97291,16.55076,17.132517,17.714273,22.641628,27.568985,32.49634,37.423695,42.35105,34.495396,26.639736,18.784079,10.928422,3.076669,3.9942036,4.911738,5.8292727,6.746807,7.6643414,7.0708723,6.481308,5.891743,5.3021784,4.7126136,3.7911747,2.87364,1.9522011,1.0307622,0.113227665,0.21864653,0.3279698,0.43338865,0.5427119,0.6481308,1.2806439,1.9092526,2.541766,3.1703746,3.7989833,3.2992198,2.7994564,2.2996929,1.7999294,1.3001659,1.097137,0.8941081,0.6910792,0.48805028,0.28892577,0.23426414,0.1835069,0.12884527,0.078088045,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,2.2918842,4.185519,6.0791545,7.968885,9.86252,8.261715,6.657006,5.056201,3.4514916,1.8506867,1.6047094,1.358732,1.116659,0.8706817,0.62470436,1.2767396,1.9248703,2.5769055,3.2250361,3.873167,5.349031,6.824895,8.300759,9.776623,11.248583,10.588739,9.924991,9.261242,8.601398,7.9376497,8.175818,8.4178915,8.65606,8.898132,9.136301,8.81614,8.492075,8.171914,7.8478484,7.523783,7.6838636,7.8400397,7.996216,8.156297,8.312472,8.386656,8.456935,8.531119,8.601398,8.675582,7.7385254,6.801469,5.8644123,4.9234514,3.9863946,3.7911747,3.59205,3.39683,3.1977055,2.998581,2.8306916,2.6667068,2.4988174,2.330928,2.1630387,2.1864653,2.2137961,2.2372224,2.260649,2.2879796,2.1278992,1.9678187,1.8077383,1.6476578,1.4875772,1.3743496,1.261122,1.1517987,1.038571,0.92534333,0.8902037,0.8550641,0.8199245,0.78478485,0.74964523,0.95657855,1.1635119,1.3743496,1.5812829,1.7882162,1.5851873,1.3821584,1.1791295,0.97610056,0.77307165,0.7145056,0.6559396,0.59346914,0.5349031,0.47633708,0.5466163,0.61689556,0.6832704,0.75354964,0.8238289,0.71841,0.61689556,0.5114767,0.40605783,0.30063897,0.43338865,0.5700427,0.7066968,0.8394465,0.97610056,1.0190489,1.0580931,1.1010414,1.1439898,1.1869383,1.6242313,2.0615244,2.4988174,2.9361105,3.3734035,3.096191,2.815074,2.533957,2.2567444,1.9756275,1.5812829,1.1869383,0.78868926,0.39434463,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.28892577,0.42557985,0.5622339,0.698888,0.8394465,0.9878138,1.1361811,1.2884527,1.43682,1.5890918,1.2767396,0.96438736,0.6481308,0.3357786,0.023426414,1.3938715,2.7604125,4.126953,5.493494,6.8639393,5.9815445,5.099149,4.2167544,3.3343596,2.4480603,7.2153354,11.978706,16.745981,21.509352,26.276627,22.782187,19.29165,15.797212,12.306676,8.812236,8.011833,7.211431,6.4110284,5.610626,4.814128,5.4115014,6.012779,6.6140575,7.211431,7.812709,7.195813,6.578918,5.958118,5.3412223,4.7243266,4.989826,5.2553253,5.520825,5.786324,6.0518236,5.919074,5.786324,5.6535745,5.520825,5.388075,5.5403466,5.6926184,5.84489,5.997162,6.1494336,5.8292727,5.5091114,5.1889505,4.8687897,4.548629,4.2167544,3.8848803,3.5530062,3.2211318,2.8892577,2.3114061,1.7335546,1.1557031,0.57785153,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.06637484,0.11713207,0.1717937,0.22255093,0.27330816,0.26159495,0.24988174,0.23816854,0.22645533,0.21083772,0.28892577,0.3631094,0.43729305,0.5114767,0.58566034,0.49195468,0.39824903,0.30063897,0.20693332,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.113227665,0.10541886,0.093705654,0.08589685,0.07418364,0.078088045,0.08589685,0.08980125,0.093705654,0.10151446,0.10151446,0.10541886,0.10932326,0.10932326,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.22645533,0.45681506,0.6832704,0.9097257,1.1361811,1.4485333,1.7608855,2.0732377,2.3855898,2.7018464,3.1781836,3.6584249,4.138666,4.618908,5.099149,5.473972,5.84489,6.2158084,6.590631,6.9615493,6.5984397,6.2314262,5.8683167,5.5013027,5.138193,5.610626,6.083059,6.5554914,7.027924,7.5003567,7.168483,6.8366084,6.5008297,6.168956,5.8370814,6.008875,6.1767645,6.348558,6.5164475,6.688241,6.6843367,6.6843367,6.6804323,6.676528,6.676528,7.016211,7.3597984,7.703386,8.043069,8.386656,7.9805984,7.578445,7.172387,6.7663293,6.364176,6.9615493,7.562827,8.164105,8.761478,9.362757,8.866898,8.371038,7.8790836,7.3832245,6.8873653,7.2348576,7.5823493,7.929841,8.277332,8.624825,8.324185,8.019642,7.719003,7.4144597,7.113821,6.5437784,5.9776397,5.4115014,4.841459,4.2753205,4.4588275,4.646239,4.829746,5.0132523,5.2006636,4.630621,4.0644827,3.4983444,2.9283018,2.3621633,3.873167,3.338264,2.7994564,2.260649,1.7257458,1.1869383,1.33921,1.4875772,1.6359446,1.7882162,1.9365835,1.7608855,1.5890918,1.4133936,1.2376955,1.0619974,1.0893283,1.1127546,1.1361811,1.1635119,1.1869383,1.1869383,1.1869383,1.1869383,1.1869383,1.1869383,1.4641509,1.737459,2.0107672,2.2879796,2.5612879,2.3621633,2.1630387,1.9639144,1.7608855,1.5617609,1.2884527,1.0112402,0.737932,0.46071947,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.42557985,0.6637484,0.9019169,1.1361811,1.3743496,1.1244678,0.8745861,0.62470436,0.37482262,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,0.26159495,0.27330816,0.28892577,0.30063897,0.31235218,0.27330816,0.23816854,0.19912452,0.1639849,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,0.26159495,0.27330816,0.28892577,0.30063897,0.31235218,0.3513962,0.38653582,0.42557985,0.46071947,0.4997635,0.5622339,0.62470436,0.6871748,0.74964523,0.81211567,0.9019169,0.9878138,1.0737107,1.1635119,1.2494087,1.2259823,1.1986516,1.175225,1.1517987,1.1244678,1.261122,1.4016805,1.5383345,1.6749885,1.8116426,1.9873407,2.1630387,2.338737,2.514435,2.6862288,2.8111696,2.9361105,3.0610514,3.1859922,3.310933,3.6740425,4.037152,4.4002614,4.7633705,5.12648,4.911738,4.7009,4.4861584,4.2753205,4.0605783,3.9746814,3.8887846,3.7989833,3.7130866,3.6232853,4.251894,4.8765984,5.5013027,6.126007,6.7507114,6.676528,6.5984397,6.524256,6.4500723,6.375889,6.5125427,6.649197,6.785851,6.9264097,7.0630636,7.211431,7.363703,7.5120697,7.6643414,7.812709,7.6252975,7.437886,7.250475,7.0630636,6.8756523,7.6370106,8.398369,9.163632,9.924991,10.686349,10.787864,10.889378,10.986988,11.088503,11.186112,11.275913,11.361811,11.4516115,11.537509,11.623405,12.173926,12.724447,13.274967,13.825488,14.376009,14.512663,14.649317,14.785972,14.92653,15.063184,15.035853,15.012426,14.989,14.96167,14.938243,15.875299,16.812357,17.749413,18.68647,19.623526,24.187773,28.748114,33.31236,37.876606,42.436947,34.22599,26.011127,17.800169,9.589212,1.3743496,2.9751544,4.575959,6.1767645,7.773665,9.37447,8.663869,7.9493628,7.238762,6.524256,5.813655,4.650143,3.4866312,2.3231194,1.1635119,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.999527,1.9365835,2.87364,3.8106966,4.7516575,4.126953,3.4983444,2.87364,2.2489357,1.6242313,1.3001659,0.97610056,0.6481308,0.3240654,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,1.9873407,3.474918,4.9624953,6.4500723,7.9376497,6.6140575,5.2865605,3.9629683,2.639376,1.3118792,1.1986516,1.0893283,0.97610056,0.8628729,0.74964523,1.5266213,2.2996929,3.076669,3.8497405,4.6267166,6.223617,7.824422,9.425227,11.0260315,12.626837,11.514082,10.401327,9.288573,8.175818,7.0630636,7.387129,7.7111945,8.039165,8.36323,8.687295,8.261715,7.8361354,7.4105554,6.98888,6.5633,6.9381227,7.3129454,7.687768,8.062591,8.437413,8.663869,8.886419,9.112875,9.339331,9.561881,8.449126,7.336372,6.223617,5.1108627,3.998108,3.8614538,3.7247996,3.5881457,3.4514916,3.310933,3.174279,3.0376248,2.900971,2.7643168,2.6237583,2.5769055,2.5261483,2.475391,2.4246337,2.3738766,2.1630387,1.9482968,1.737459,1.5266213,1.3118792,1.2767396,1.2376955,1.1986516,1.1635119,1.1244678,0.97610056,0.8238289,0.6754616,0.5231899,0.37482262,0.5388075,0.698888,0.8628729,1.0268579,1.1869383,1.1127546,1.038571,0.96438736,0.8862993,0.81211567,0.737932,0.6637484,0.58566034,0.5114767,0.43729305,0.5388075,0.63641757,0.737932,0.8394465,0.93705654,0.81211567,0.6871748,0.5622339,0.43729305,0.31235218,0.46071947,0.61299115,0.76135844,0.9136301,1.0619974,1.0737107,1.0893283,1.1010414,1.1127546,1.1244678,1.6359446,2.1513257,2.6628022,3.174279,3.6857557,3.435874,3.1859922,2.9361105,2.6862288,2.436347,1.9482968,1.4641509,0.97610056,0.48805028,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0268579,2.0498111,3.076669,4.0996222,5.12648,4.7009,4.2753205,3.8497405,3.4241607,2.998581,7.601871,12.201257,16.800642,21.400028,25.999414,22.813423,19.623526,16.437534,13.251541,10.061645,8.937177,7.812709,6.688241,5.563773,4.4393053,5.1889505,5.938596,6.688241,7.437886,8.187531,7.387129,6.5867267,5.786324,4.985922,4.1894236,4.5993857,5.0132523,5.423215,5.8370814,6.250948,6.086963,5.9268827,5.7628975,5.5989127,5.4388323,5.700427,5.9620223,6.223617,6.4891167,6.7507114,6.387602,6.0244927,5.661383,5.298274,4.939069,4.548629,4.1620927,3.775557,3.3890212,2.998581,2.4012074,1.7999294,1.1986516,0.60127795,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.13665408,0.27330816,0.41386664,0.5505207,0.6871748,1.0619974,1.43682,1.8116426,2.1864653,2.5612879,2.912684,3.2640803,3.611572,3.9629683,4.3143644,4.825841,5.337318,5.8487945,6.364176,6.8756523,6.4500723,6.0244927,5.5989127,5.173333,4.7516575,5.251421,5.7511845,6.250948,6.7507114,7.250475,6.98888,6.7233806,6.461786,6.2001905,5.938596,6.1494336,6.364176,6.575013,6.785851,7.000593,7.098203,7.1997175,7.3012323,7.3988423,7.5003567,7.8868923,8.273428,8.663869,9.050405,9.43694,9.01136,8.58578,8.164105,7.7385254,7.3129454,8.062591,8.812236,9.561881,10.311526,11.061172,10.487225,9.913278,9.339331,8.761478,8.187531,8.312472,8.437413,8.562354,8.687295,8.812236,8.52331,8.238289,7.9493628,7.6643414,7.375416,6.6257706,5.8761253,5.12648,4.376835,3.6232853,3.951255,4.2753205,4.5993857,4.9234514,5.251421,4.73604,4.224563,3.7130866,3.2016098,2.6862288,3.1391394,2.7135596,2.2918842,1.8702087,1.4485333,1.0268579,1.1635119,1.3001659,1.43682,1.5734742,1.7140326,1.5461433,1.3821584,1.2181735,1.0541886,0.8862993,0.9136301,0.93705654,0.96438736,0.9878138,1.0112402,1.0463798,1.0815194,1.116659,1.1517987,1.1869383,1.3860629,1.5812829,1.7804074,1.9756275,2.174752,1.999054,1.8194515,1.6437533,1.4641509,1.2884527,1.0580931,0.8316377,0.60518235,0.37872702,0.14836729,0.13274968,0.113227665,0.09761006,0.078088045,0.062470436,0.10151446,0.14055848,0.1835069,0.22255093,0.26159495,0.49195468,0.7223144,0.95267415,1.183034,1.4133936,1.1557031,0.8980125,0.64032197,0.38263142,0.12494087,0.10151446,0.078088045,0.058566034,0.03513962,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.10151446,0.20693332,0.30844778,0.40996224,0.5114767,0.42557985,0.3357786,0.24988174,0.1639849,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.058566034,0.10151446,0.14836729,0.19131571,0.23816854,0.20693332,0.1756981,0.14836729,0.11713207,0.08589685,0.10932326,0.13274968,0.15617609,0.1756981,0.19912452,0.21864653,0.23816854,0.26159495,0.28111696,0.30063897,0.29283017,0.28502136,0.27721256,0.26940376,0.26159495,0.23426414,0.20302892,0.1717937,0.14055848,0.113227665,0.10932326,0.10932326,0.10541886,0.10151446,0.10151446,0.113227665,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,0.26159495,0.27330816,0.28892577,0.3240654,0.3631094,0.39824903,0.43729305,0.47633708,0.5388075,0.60518235,0.6715572,0.7340276,0.80040246,0.8941081,0.9917182,1.0854238,1.1791295,1.2767396,1.2806439,1.2845483,1.2884527,1.2962615,1.3001659,1.4016805,1.5031948,1.6086137,1.7101282,1.8116426,1.9443923,2.077142,2.2098918,2.3426414,2.475391,2.6081407,2.7447948,2.8814487,3.0141985,3.1508527,3.5647192,3.978586,4.396357,4.8102236,5.22409,4.997635,4.7711797,4.5408196,4.3143644,4.087909,3.9942036,3.8965936,3.802888,3.7091823,3.611572,4.0918136,4.5681505,5.044488,5.520825,6.001066,5.958118,5.919074,5.8800297,5.840986,5.801942,5.919074,6.036206,6.153338,6.27047,6.387602,6.5633,6.7429028,6.918601,7.098203,7.2739015,7.0630636,6.8561306,6.6452928,6.434455,6.223617,6.9810715,7.734621,8.488171,9.245625,9.999174,10.09288,10.186585,10.276386,10.370092,10.4637985,10.487225,10.510651,10.537982,10.561408,10.588739,11.373524,12.158309,12.943093,13.727879,14.512663,14.528281,14.543899,14.555612,14.571229,14.586847,14.582942,14.579038,14.571229,14.567325,14.56342,15.629322,16.69913,17.76503,18.830933,19.900738,22.83685,25.769054,28.705166,31.641275,34.573483,27.881336,21.185287,14.489237,7.793187,1.1010414,2.3816853,3.6584249,4.939069,6.2197127,7.5003567,7.0240197,6.5437784,6.067441,5.591104,5.1108627,4.0918136,3.06886,2.0459068,1.0229534,0.0,0.13665408,0.26940376,0.40605783,0.5388075,0.6754616,1.3274968,1.979532,2.631567,3.2836022,3.9356375,3.408543,2.8814487,2.3543546,1.8272603,1.3001659,1.038571,0.78088045,0.5192855,0.26159495,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18741131,0.37482262,0.5622339,0.74964523,0.93705654,2.194274,3.4514916,4.7087092,5.9659266,7.223144,6.0518236,4.8765984,3.7013733,2.5261483,1.3509232,2.1786566,3.0102942,3.8419318,4.6696653,5.5013027,5.376362,5.251421,5.12648,5.001539,4.8765984,6.17286,7.4691215,8.769287,10.065549,11.361811,10.48332,9.600925,8.722435,7.843944,6.9615493,7.1099167,7.2582836,7.406651,7.551114,7.699481,7.363703,7.0240197,6.688241,6.348558,6.012779,6.356367,6.703859,7.0474463,7.3910336,7.7385254,7.9064145,8.074304,8.238289,8.406178,8.574067,7.6838636,6.7897553,5.8956475,5.0054436,4.1113358,3.959064,3.802888,3.6467118,3.49444,3.338264,3.174279,3.0141985,2.8502135,2.6862288,2.5261483,2.494913,2.463678,2.436347,2.4051118,2.3738766,2.1708477,1.9639144,1.7608855,1.5539521,1.3509232,1.3157835,1.2806439,1.2455044,1.2103647,1.175225,1.038571,0.9058213,0.76916724,0.63641757,0.4997635,0.62470436,0.74964523,0.8745861,0.999527,1.1244678,1.0424755,0.96048295,0.8784905,0.79649806,0.7106012,0.6637484,0.61689556,0.5700427,0.5231899,0.47633708,0.5583295,0.6442264,0.7301232,0.8160201,0.9019169,0.78868926,0.6754616,0.5622339,0.44900626,0.3357786,0.5153811,0.6910792,0.8706817,1.0463798,1.2259823,1.1713207,1.116659,1.0580931,1.0034313,0.94876975,1.3782539,1.8116426,2.241127,2.6706111,3.1000953,2.9087796,2.7213683,2.5300527,2.338737,2.1513257,1.8741131,1.6008049,1.3235924,1.0502841,0.77307165,0.6481308,0.5231899,0.39824903,0.27330816,0.14836729,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.113227665,0.20693332,0.29673457,0.38653582,0.47633708,0.5661383,0.659844,0.75354964,0.8433509,0.93705654,1.8194515,2.7018464,3.5842414,4.466636,5.349031,4.8492675,4.3455997,3.8419318,3.338264,2.8385005,6.7702336,10.701966,14.633699,18.569338,22.50107,20.006157,17.511244,15.016331,12.521418,10.0265045,8.921559,7.8205175,6.715572,5.6145306,4.513489,5.1772375,5.840986,6.5086384,7.172387,7.8361354,7.066968,6.297801,5.5286336,4.755562,3.9863946,4.3065557,4.6267166,4.9468775,5.267039,5.5871997,5.4310236,5.278752,5.1225758,4.9663997,4.814128,4.93126,5.0483923,5.165524,5.282656,5.3997884,5.1303844,4.860981,4.591577,4.318269,4.0488653,3.7208953,3.3890212,3.0610514,2.7291772,2.4012074,1.9209659,1.4407244,0.96048295,0.48024148,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05466163,0.058566034,0.06637484,0.07027924,0.07418364,0.093705654,0.10932326,0.12884527,0.14446288,0.1639849,0.14055848,0.12103647,0.10151446,0.08199245,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.12103647,0.24597734,0.3670138,0.48805028,0.61299115,0.98000497,1.3470187,1.7140326,2.0810463,2.4480603,2.7994564,3.1508527,3.4983444,3.8497405,4.2011366,4.591577,4.985922,5.376362,5.7707067,6.1611466,5.9346914,5.708236,5.481781,5.251421,5.024966,5.5013027,5.9737353,6.4500723,6.9264097,7.3988423,7.1762915,6.949836,6.7233806,6.5008297,6.2743745,6.5437784,6.813182,7.08649,7.355894,7.6252975,7.793187,7.9649806,8.136774,8.304664,8.476458,8.663869,8.85128,9.0386915,9.226103,9.413514,9.269051,9.128492,8.98403,8.843472,8.699008,9.058213,9.413514,9.772718,10.131924,10.487225,9.921086,9.358852,8.792714,8.226576,7.6643414,7.746334,7.8283267,7.910319,7.9923115,8.074304,7.9220324,7.7697606,7.617489,7.465217,7.3129454,6.5008297,5.6926184,4.884407,4.0722914,3.2640803,3.4788225,3.6935644,3.9083066,4.123049,4.337791,3.9356375,3.5373883,3.1391394,2.736986,2.338737,2.4012074,2.0927596,1.7843118,1.475864,1.1713207,0.8628729,0.9878138,1.1127546,1.2376955,1.3626363,1.4875772,1.3314011,1.1791295,1.0229534,0.8667773,0.7106012,0.737932,0.76135844,0.78868926,0.81211567,0.8394465,0.9058213,0.97610056,1.0463798,1.116659,1.1869383,1.3079748,1.4290112,1.5461433,1.6671798,1.7882162,1.6320401,1.475864,1.3235924,1.1674163,1.0112402,0.8316377,0.6520352,0.47243267,0.29283017,0.113227665,0.113227665,0.11713207,0.12103647,0.12103647,0.12494087,0.1678893,0.21083772,0.25378615,0.29673457,0.3357786,0.5583295,0.78088045,1.0034313,1.2259823,1.4485333,1.1869383,0.92143893,0.6559396,0.39044023,0.12494087,0.10541886,0.08589685,0.06637484,0.046852827,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,0.3513962,0.30063897,0.24988174,0.19912452,0.14836729,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.06637484,0.10541886,0.14446288,0.1835069,0.22645533,0.20302892,0.1796025,0.15617609,0.13665408,0.113227665,0.13274968,0.15227169,0.1717937,0.19131571,0.21083772,0.23816854,0.26940376,0.29673457,0.3240654,0.3513962,0.3240654,0.29673457,0.26940376,0.23816854,0.21083772,0.19131571,0.1678893,0.14446288,0.12103647,0.10151446,0.093705654,0.08980125,0.08589685,0.078088045,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,0.26159495,0.30063897,0.3357786,0.37482262,0.41386664,0.44900626,0.5192855,0.58566034,0.6520352,0.71841,0.78868926,0.8902037,0.9917182,1.0932326,1.1986516,1.3001659,1.3353056,1.3704453,1.4055848,1.4407244,1.475864,1.542239,1.6086137,1.678893,1.7452679,1.8116426,1.901444,1.9912452,2.0810463,2.1708477,2.260649,2.4090161,2.5534792,2.697942,2.8424048,2.9868677,3.455396,3.9239242,4.388548,4.8570766,5.3256044,5.083532,4.841459,4.5993857,4.3534083,4.1113358,4.009821,3.9083066,3.8067923,3.7013733,3.5998588,3.9317331,4.2597027,4.591577,4.919547,5.251421,5.2436123,5.239708,5.2358036,5.2318993,5.22409,5.3217,5.4193106,5.5169206,5.6145306,5.7121406,5.919074,6.1221027,6.329036,6.532065,6.7389984,6.504734,6.2743745,6.04011,5.805846,5.575486,6.321227,7.0708723,7.816613,8.566258,9.311999,9.397896,9.483793,9.565785,9.651682,9.737579,9.698535,9.663396,9.6243515,9.589212,9.550168,10.569217,11.588266,12.611219,13.630268,14.649317,14.543899,14.434575,14.329156,14.219833,14.114414,14.126127,14.141745,14.157363,14.17298,14.188598,15.383345,16.581997,17.780647,18.9793,20.174046,21.482021,22.789995,24.097971,25.405945,26.71392,21.536682,16.359446,11.178304,6.001066,0.8238289,1.7843118,2.7447948,3.7052777,4.6657605,5.6262436,5.3841705,5.138193,4.8961205,4.6540475,4.4119744,3.5295796,2.6471848,1.7647898,0.8823949,0.0,0.25769055,0.5153811,0.77307165,1.0307622,1.2884527,1.6554666,2.0224805,2.3894942,2.7565079,3.1235218,2.6940374,2.2645533,1.8350691,1.4055848,0.97610056,0.78088045,0.58566034,0.39044023,0.19522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.27330816,0.5505207,0.8238289,1.1010414,1.3743496,2.4012074,3.4280653,4.4588275,5.4856853,6.5125427,5.4856853,4.462732,3.435874,2.4129205,1.3860629,3.1586614,4.93126,6.703859,8.476458,10.249056,9.226103,8.1992445,7.1762915,6.1494336,5.12648,6.1181984,7.113821,8.109444,9.105066,10.100689,9.452558,8.804427,8.156297,7.5081654,6.8639393,6.832704,6.801469,6.774138,6.7429028,6.7116675,6.461786,6.211904,5.9620223,5.7121406,5.462259,5.7785153,6.0908675,6.407124,6.7233806,7.0357327,7.1489606,7.2582836,7.367607,7.47693,7.5862536,6.914696,6.2431393,5.571582,4.8961205,4.224563,4.0527697,3.8809757,3.7091823,3.533484,3.3616903,3.174279,2.9868677,2.7994564,2.612045,2.4246337,2.416825,2.4051118,2.3933985,2.3855898,2.3738766,2.1786566,1.979532,1.7843118,1.5851873,1.3860629,1.3548276,1.3235924,1.2884527,1.2572175,1.2259823,1.1049459,0.98390937,0.8667773,0.74574083,0.62470436,0.7106012,0.80040246,0.8862993,0.97610056,1.0619974,0.97219616,0.8823949,0.79259366,0.7027924,0.61299115,0.59346914,0.57394713,0.5544251,0.5309987,0.5114767,0.58175594,0.6520352,0.7223144,0.79259366,0.8628729,0.76135844,0.6637484,0.5622339,0.46071947,0.3631094,0.5661383,0.77307165,0.97610056,1.183034,1.3860629,1.2650263,1.1439898,1.0190489,0.8980125,0.77307165,1.1244678,1.4680552,1.8194515,2.1669433,2.514435,2.3816853,2.25284,2.1239948,1.9912452,1.8623998,1.7999294,1.737459,1.6749885,1.6125181,1.5500476,1.261122,0.97610056,0.6871748,0.39824903,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.23035973,0.40996224,0.58956474,0.76916724,0.94876975,1.1361811,1.319688,1.5031948,1.6906061,1.8741131,2.6159496,3.3538816,4.095718,4.83365,5.575486,4.9937305,4.415879,3.8341231,3.2562714,2.6745155,5.938596,9.20658,12.470661,15.734741,18.998821,17.198893,15.395058,13.591225,11.791295,9.987461,8.905942,7.8283267,6.746807,5.6691923,4.5876727,5.169429,5.74728,6.329036,6.9068875,7.4886436,6.746807,6.008875,5.267039,4.5291066,3.78727,4.0137253,4.2440853,4.4705405,4.6969957,4.9234514,4.7789884,4.630621,4.482254,4.3338866,4.1894236,4.1581883,4.1308575,4.1035266,4.0761957,4.0488653,3.873167,3.6935644,3.5178664,3.338264,3.1625657,2.8892577,2.6159496,2.3465457,2.0732377,1.7999294,1.4407244,1.0815194,0.71841,0.359205,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.046852827,0.058566034,0.06637484,0.078088045,0.08589685,0.10932326,0.13274968,0.15617609,0.1756981,0.19912452,0.1717937,0.14446288,0.11713207,0.08980125,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.10932326,0.21474212,0.3240654,0.42948425,0.5388075,0.8980125,1.2572175,1.6164225,1.9756275,2.338737,2.6862288,3.0376248,3.3890212,3.736513,4.087909,4.3612175,4.630621,4.903929,5.1772375,5.4505453,5.4193106,5.388075,5.3607445,5.3295093,5.298274,5.7511845,6.2001905,6.649197,7.098203,7.551114,7.363703,7.1762915,6.98888,6.801469,6.6140575,6.9381227,7.266093,7.5940623,7.9220324,8.250002,8.488171,8.730244,8.968412,9.2104845,9.448653,9.43694,9.425227,9.413514,9.4018,9.386183,9.526741,9.6673,9.807858,9.948417,10.088976,10.053836,10.018696,9.983557,9.948417,9.913278,9.358852,8.800523,8.246098,7.6916723,7.137247,7.1762915,7.2192397,7.2582836,7.297328,7.336372,7.320754,7.3012323,7.2856145,7.266093,7.250475,6.379793,5.5091114,4.6384296,3.7716527,2.900971,3.0063896,3.1118085,3.213323,3.3187418,3.4241607,3.1391394,2.8502135,2.5612879,2.2762666,1.9873407,1.6632754,1.4680552,1.2767396,1.0854238,0.8941081,0.698888,0.81211567,0.92534333,1.038571,1.1517987,1.261122,1.116659,0.97219616,0.8277333,0.6832704,0.5388075,0.5622339,0.58566034,0.61299115,0.63641757,0.6637484,0.76916724,0.8706817,0.97610056,1.0815194,1.1869383,1.2298868,1.2728351,1.3157835,1.358732,1.4016805,1.2689307,1.1361811,1.0034313,0.8706817,0.737932,0.60518235,0.47243267,0.339683,0.20693332,0.07418364,0.09761006,0.12103647,0.14055848,0.1639849,0.18741131,0.23426414,0.27721256,0.3240654,0.3670138,0.41386664,0.62860876,0.8433509,1.0580931,1.2728351,1.4875772,1.2142692,0.94096094,0.6715572,0.39824903,0.12494087,0.10932326,0.08980125,0.07418364,0.05466163,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.058566034,0.113227665,0.1717937,0.23035973,0.28892577,0.27330816,0.26159495,0.24988174,0.23816854,0.22645533,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.07418364,0.10932326,0.14055848,0.1756981,0.21083772,0.19912452,0.1835069,0.1678893,0.15227169,0.13665408,0.15617609,0.1717937,0.19131571,0.20693332,0.22645533,0.26159495,0.29673457,0.3318742,0.3631094,0.39824903,0.3513962,0.30454338,0.25769055,0.21083772,0.1639849,0.14836729,0.13274968,0.11713207,0.10151446,0.08589685,0.078088045,0.07418364,0.06637484,0.058566034,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.27330816,0.31235218,0.3513962,0.38653582,0.42557985,0.4958591,0.5661383,0.63641757,0.7066968,0.77307165,0.8862993,0.9956226,1.1049459,1.2142692,1.3235924,1.3899672,1.456342,1.5188124,1.5851873,1.6515622,1.6827974,1.7140326,1.7491722,1.7804074,1.8116426,1.8584955,1.9092526,1.9561055,2.0029583,2.0498111,2.2059872,2.358259,2.514435,2.6706111,2.8267872,3.3460727,3.8653584,4.3846436,4.903929,5.423215,5.169429,4.911738,4.6540475,4.396357,4.138666,4.029343,3.9161155,3.8067923,3.697469,3.5881457,3.7716527,3.951255,4.134762,4.318269,4.5017757,4.5291066,4.560342,4.591577,4.618908,4.650143,4.728231,4.806319,4.884407,4.958591,5.036679,5.270943,5.5013027,5.735567,5.9659266,6.2001905,5.9464045,5.688714,5.434928,5.181142,4.9234514,5.6652875,6.4032197,7.1450562,7.8868923,8.624825,8.702912,8.781001,8.859089,8.933272,9.01136,8.913751,8.812236,8.710721,8.6131115,8.511597,9.768814,11.022127,12.2793455,13.532659,14.785972,14.555612,14.329156,14.098797,13.868437,13.638077,13.673217,13.708356,13.743496,13.778636,13.813775,15.141272,16.46877,17.796265,19.123762,20.45126,20.131098,19.810938,19.490776,19.170614,18.850454,15.188125,11.5297,7.871275,4.2089458,0.5505207,1.1908426,1.8311646,2.4714866,3.1118085,3.7482262,3.7443218,3.736513,3.7287042,3.7208953,3.7130866,2.97125,2.2294137,1.4836729,0.7418364,0.0,0.37872702,0.76135844,1.1400855,1.5188124,1.901444,1.9834363,2.0654287,2.1474214,2.2294137,2.3114061,1.979532,1.6476578,1.3157835,0.98390937,0.6481308,0.5192855,0.39044023,0.26159495,0.12884527,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3631094,0.7262188,1.0893283,1.4485333,1.8116426,2.6081407,3.408543,4.2050414,5.001539,5.801942,4.9234514,4.0488653,3.174279,2.2996929,1.4251068,4.138666,6.8561306,9.56969,12.28325,15.000713,13.075843,11.150972,9.226103,7.3012323,5.376362,6.067441,6.75852,7.453504,8.144583,8.835662,8.421796,8.007929,7.5940623,7.1762915,6.7624245,6.5554914,6.348558,6.141625,5.930787,5.7238536,5.563773,5.3997884,5.2358036,5.0757227,4.911738,5.196759,5.481781,5.7668023,6.0518236,6.336845,6.3915067,6.4422636,6.4969254,6.547683,6.5984397,6.1455293,5.6965227,5.2436123,4.7907014,4.337791,4.1464753,3.959064,3.767748,3.5764325,3.3890212,3.174279,2.9634414,2.7486992,2.5378613,2.3231194,2.3348327,2.3465457,2.3543546,2.366068,2.3738766,2.1864653,1.9951496,1.8038338,1.6164225,1.4251068,1.3938715,1.3665408,1.3353056,1.3040704,1.2767396,1.1713207,1.0659018,0.96048295,0.8550641,0.74964523,0.80040246,0.8511597,0.9019169,0.94876975,0.999527,0.9019169,0.80430686,0.7066968,0.60908675,0.5114767,0.5192855,0.5270943,0.5349031,0.5427119,0.5505207,0.60518235,0.659844,0.7145056,0.76916724,0.8238289,0.737932,0.6481308,0.5622339,0.47633708,0.38653582,0.62079996,0.8511597,1.0854238,1.3157835,1.5500476,1.358732,1.1713207,0.98000497,0.78868926,0.60127795,0.8667773,1.1283722,1.3938715,1.6593709,1.9248703,1.8545911,1.7843118,1.7140326,1.6437533,1.5734742,1.7257458,1.8741131,2.0263848,2.174752,2.3231194,1.8741131,1.4251068,0.97610056,0.5231899,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.3435874,0.61689556,0.8862993,1.1557031,1.4251068,1.7023194,1.979532,2.2567444,2.533957,2.8111696,3.408543,4.0059166,4.60329,5.2006636,5.801942,5.142098,4.4861584,3.8263142,3.1703746,2.514435,5.1108627,7.70729,10.303718,12.90405,15.500477,14.391626,13.2788725,12.170022,11.061172,9.948417,8.894228,7.8361354,6.7780423,5.7199492,4.661856,5.1577153,5.6535745,6.1494336,6.6413884,7.137247,6.426646,5.716045,5.009348,4.298747,3.5881457,3.7208953,3.8575494,3.9942036,4.126953,4.263607,4.123049,3.9824903,3.8419318,3.7013733,3.5608149,3.3890212,3.2172275,3.0454338,2.87364,2.7018464,2.6159496,2.5300527,2.4441557,2.358259,2.2762666,2.0615244,1.8467822,1.6281357,1.4133936,1.1986516,0.96048295,0.71841,0.48024148,0.23816854,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.039044023,0.05466163,0.07027924,0.08589685,0.10151446,0.12884527,0.15617609,0.1835069,0.21083772,0.23816854,0.20302892,0.1678893,0.13274968,0.09761006,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.093705654,0.1835069,0.27721256,0.3709182,0.46071947,0.8160201,1.1674163,1.5188124,1.8741131,2.2255092,2.5769055,2.9243972,3.2757936,3.6232853,3.9746814,4.126953,4.279225,4.4314966,4.5837684,4.73604,4.903929,5.0718184,5.239708,5.407597,5.575486,6.001066,6.426646,6.8483214,7.2739015,7.699481,7.551114,7.3988423,7.250475,7.098203,6.949836,7.336372,7.719003,8.105539,8.488171,8.874706,9.183154,9.495506,9.803954,10.116306,10.424754,10.213917,9.999174,9.788337,9.573594,9.362757,9.784432,10.206107,10.631687,11.053363,11.475039,11.045554,10.619974,10.194394,9.76491,9.339331,8.792714,8.246098,7.703386,7.1567693,6.6140575,6.610153,6.606249,6.606249,6.602344,6.5984397,6.715572,6.8366084,6.9537406,7.0708723,7.1880045,6.2587566,5.3256044,4.396357,3.4671092,2.5378613,2.533957,2.5261483,2.522244,2.5183394,2.514435,2.338737,2.1630387,1.9873407,1.8116426,1.6359446,0.92534333,0.8472553,0.76916724,0.6910792,0.61689556,0.5388075,0.63641757,0.737932,0.8394465,0.93705654,1.038571,0.9019169,0.76916724,0.63251317,0.4958591,0.3631094,0.38653582,0.41386664,0.43729305,0.46071947,0.48805028,0.62860876,0.76916724,0.9058213,1.0463798,1.1869383,1.1517987,1.116659,1.0815194,1.0463798,1.0112402,0.9019169,0.79259366,0.6832704,0.57394713,0.46071947,0.37872702,0.29283017,0.20693332,0.12103647,0.039044023,0.078088045,0.12103647,0.1639849,0.20693332,0.24988174,0.29673457,0.3435874,0.39434463,0.44119745,0.48805028,0.6949836,0.9019169,1.1088502,1.3157835,1.5266213,1.2455044,0.96438736,0.6832704,0.40605783,0.12494087,0.10932326,0.093705654,0.078088045,0.06637484,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.19912452,0.22645533,0.24988174,0.27330816,0.30063897,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.078088045,0.10932326,0.14055848,0.1717937,0.19912452,0.19131571,0.1835069,0.1756981,0.1717937,0.1639849,0.1756981,0.19131571,0.20693332,0.22255093,0.23816854,0.28111696,0.3240654,0.3631094,0.40605783,0.44900626,0.38263142,0.31625658,0.24597734,0.1796025,0.113227665,0.10541886,0.09761006,0.08980125,0.08199245,0.07418364,0.06637484,0.05466163,0.046852827,0.03513962,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.19912452,0.21083772,0.24988174,0.28892577,0.3240654,0.3631094,0.39824903,0.47243267,0.5466163,0.61689556,0.6910792,0.76135844,0.8784905,0.9956226,1.116659,1.2337911,1.3509232,1.4446288,1.5383345,1.6359446,1.7296503,1.8233559,1.8233559,1.8194515,1.8194515,1.815547,1.8116426,1.8194515,1.8233559,1.8272603,1.8311646,1.8389735,2.0029583,2.1669433,2.330928,2.4988174,2.6628022,3.2367494,3.8067923,4.380739,4.950782,5.5247293,5.251421,4.9781127,4.7087092,4.435401,4.1620927,4.044961,3.9278288,3.8106966,3.6935644,3.5764325,3.611572,3.6467118,3.6818514,3.7130866,3.7482262,3.814601,3.8809757,3.9434462,4.009821,4.0761957,4.1308575,4.1894236,4.2479897,4.3065557,4.3612175,4.6228123,4.884407,5.142098,5.4036927,5.661383,5.3841705,5.1069584,4.829746,4.552533,4.2753205,5.009348,5.7394714,6.473499,7.2036223,7.9376497,8.007929,8.078208,8.148487,8.218767,8.289046,8.125061,7.9610763,7.800996,7.6370106,7.47693,8.964508,10.455989,11.943566,13.435048,14.92653,14.571229,14.219833,13.868437,13.513136,13.16174,13.216402,13.271063,13.325725,13.384291,13.438952,14.895294,16.351637,17.811884,19.268225,20.724567,18.77627,16.831879,14.883581,12.935285,10.986988,8.843472,6.703859,4.560342,2.416825,0.27330816,0.59346914,0.9136301,1.2337911,1.5539521,1.8741131,2.1005683,2.330928,2.5573835,2.7838387,3.0141985,2.4090161,1.8077383,1.2064602,0.60127795,0.0,0.5036679,1.0034313,1.5070993,2.0107672,2.514435,2.3114061,2.1083772,1.9053483,1.7023194,1.4992905,1.2650263,1.0307622,0.79649806,0.5583295,0.3240654,0.26159495,0.19522011,0.12884527,0.06637484,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.44900626,0.9019169,1.3509232,1.7999294,2.2489357,2.8189783,3.3851168,3.951255,4.521298,5.087436,4.3612175,3.638903,2.912684,2.1864653,1.4641509,5.1186714,8.777096,12.435521,16.093946,19.748466,16.925583,14.098797,11.275913,8.449126,5.6262436,6.016684,6.4032197,6.79366,7.1841,7.57454,7.3910336,7.211431,7.027924,6.844417,6.66091,6.278279,5.891743,5.5091114,5.1225758,4.73604,4.661856,4.5876727,4.513489,4.4393053,4.3612175,4.618908,4.872694,5.12648,5.3841705,5.6379566,5.6340523,5.6262436,5.6223392,5.618435,5.610626,5.380266,5.1460023,4.9156423,4.6813784,4.4510183,4.2440853,4.0332475,3.8263142,3.619381,3.4124475,3.174279,2.9361105,2.7018464,2.463678,2.2255092,2.2567444,2.2840753,2.3153105,2.3465457,2.3738766,2.194274,2.0107672,1.8272603,1.6437533,1.4641509,1.43682,1.4055848,1.3782539,1.3509232,1.3235924,1.2337911,1.1439898,1.0541886,0.96438736,0.8745861,0.8862993,0.9019169,0.9136301,0.92534333,0.93705654,0.8316377,0.7262188,0.62079996,0.5192855,0.41386664,0.44900626,0.48414588,0.5192855,0.5544251,0.58566034,0.62860876,0.6676528,0.7066968,0.74574083,0.78868926,0.7106012,0.63641757,0.5622339,0.48805028,0.41386664,0.6715572,0.93315214,1.1908426,1.4524376,1.7140326,1.456342,1.1986516,0.94096094,0.6832704,0.42557985,0.60908675,0.78868926,0.97219616,1.1557031,1.33921,1.3274968,1.3157835,1.3079748,1.2962615,1.2884527,1.6515622,2.0107672,2.3738766,2.736986,3.1000953,2.4871042,1.8741131,1.261122,0.6481308,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.46071947,0.8199245,1.1791295,1.5383345,1.901444,2.2684577,2.639376,3.0102942,3.3812122,3.7482262,4.2050414,4.661856,5.114767,5.571582,6.0244927,5.290465,4.5564375,3.8185053,3.084478,2.35045,4.279225,6.2079997,8.140678,10.069453,11.998228,11.584361,11.166591,10.748819,10.331048,9.913278,8.878611,7.843944,6.8092775,5.7707067,4.73604,5.1460023,5.5559645,5.9659266,6.375889,6.785851,6.1064854,5.4271193,4.747753,4.068387,3.3890212,3.4280653,3.4710135,3.513962,3.5569105,3.5998588,3.4671092,3.3343596,3.2016098,3.06886,2.9361105,2.619854,2.3035975,1.9834363,1.6671798,1.3509232,1.358732,1.3665408,1.3743496,1.3782539,1.3860629,1.2298868,1.0737107,0.9136301,0.75745404,0.60127795,0.48024148,0.359205,0.23816854,0.12103647,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.031235218,0.05075723,0.07418364,0.093705654,0.113227665,0.14446288,0.1756981,0.21083772,0.24207294,0.27330816,0.23426414,0.19131571,0.14836729,0.10541886,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.078088045,0.15617609,0.23426414,0.30844778,0.38653582,0.7340276,1.077615,1.4212024,1.7686942,2.1122816,2.463678,2.8111696,3.1625657,3.513962,3.8614538,3.8965936,3.9278288,3.959064,3.9942036,4.025439,4.388548,4.755562,5.1186714,5.4856853,5.8487945,6.250948,6.649197,7.0513506,7.4495993,7.8517528,7.7385254,7.6252975,7.5120697,7.3988423,7.2856145,7.7307167,8.171914,8.6131115,9.058213,9.499411,9.878138,10.260769,10.639496,11.018223,11.400854,10.986988,10.573121,10.163159,9.749292,9.339331,10.042123,10.748819,11.4516115,12.158309,12.861101,12.041177,11.221252,10.401327,9.581403,8.761478,8.226576,7.6916723,7.1567693,6.621866,6.086963,6.044015,5.997162,5.9542136,5.9073606,5.8644123,6.114294,6.36808,6.621866,6.871748,7.125534,6.133816,5.1460023,4.154284,3.1664703,2.174752,2.0615244,1.9443923,1.8311646,1.7140326,1.6008049,1.5383345,1.475864,1.4133936,1.3509232,1.2884527,0.18741131,0.22645533,0.26159495,0.30063897,0.3357786,0.37482262,0.46071947,0.5505207,0.63641757,0.7262188,0.81211567,0.6871748,0.5622339,0.43729305,0.31235218,0.18741131,0.21083772,0.23816854,0.26159495,0.28892577,0.31235218,0.48805028,0.6637484,0.8394465,1.0112402,1.1869383,1.0737107,0.96438736,0.8511597,0.737932,0.62470436,0.5388075,0.44900626,0.3631094,0.27330816,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.3631094,0.41386664,0.46071947,0.5114767,0.5622339,0.76135844,0.96438736,1.1635119,1.3626363,1.5617609,1.2767396,0.9878138,0.698888,0.41386664,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.37482262,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,0.30063897,0.3513962,0.39824903,0.44900626,0.4997635,0.41386664,0.3240654,0.23816854,0.14836729,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.22645533,0.26159495,0.30063897,0.3357786,0.37482262,0.44900626,0.5231899,0.60127795,0.6754616,0.74964523,0.8745861,0.999527,1.1244678,1.2494087,1.3743496,1.4992905,1.6242313,1.7491722,1.8741131,1.999054,1.9639144,1.9248703,1.8858263,1.8506867,1.8116426,1.7765031,1.737459,1.698415,1.6632754,1.6242313,1.7999294,1.9756275,2.1513257,2.3231194,2.4988174,3.1235218,3.7482262,4.376835,5.001539,5.6262436,5.337318,5.0483923,4.7633705,4.474445,4.1894236,4.0605783,3.9356375,3.8106966,3.6857557,3.5608149,3.4514916,3.338264,3.2250361,3.1118085,2.998581,3.1000953,3.2016098,3.2992198,3.4007344,3.4983444,3.5373883,3.5764325,3.611572,3.6506162,3.6857557,3.9746814,4.263607,4.548629,4.8375545,5.12648,4.825841,4.5252023,4.224563,3.9239242,3.6232853,4.349504,5.0757227,5.801942,6.524256,7.250475,7.3129454,7.375416,7.437886,7.5003567,7.562827,7.336372,7.113821,6.8873653,6.66091,6.4383593,8.164105,9.885946,11.611692,13.337439,15.063184,14.586847,14.114414,13.638077,13.16174,12.689307,12.763491,12.837675,12.911859,12.986042,13.06413,14.649317,16.238409,17.823597,19.412687,21.00178,17.425346,13.848915,10.276386,6.699954,3.1235218,2.4988174,1.8741131,1.2494087,0.62470436,0.0,0.0,0.0,0.0,0.0,0.0,0.46071947,0.92534333,1.3860629,1.8506867,2.3114061,1.8506867,1.3860629,0.92534333,0.46071947,0.0,0.62470436,1.2494087,1.8741131,2.4988174,3.1235218,2.639376,2.1513257,1.6632754,1.175225,0.6871748,0.5505207,0.41386664,0.27330816,0.13665408,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5388075,1.0737107,1.6125181,2.1513257,2.6862288,3.0259118,3.3616903,3.7013733,4.037152,4.376835,3.7989833,3.2250361,2.6510892,2.0732377,1.4992905,6.098676,10.698062,15.3013525,19.900738,24.500124,20.775324,17.050524,13.325725,9.600925,5.8761253,5.9620223,6.0518236,6.13772,6.223617,6.3134184,6.364176,6.4110284,6.461786,6.5125427,6.5633,6.001066,5.4388323,4.8765984,4.3143644,3.7482262,3.7638438,3.775557,3.78727,3.7989833,3.8106966,4.037152,4.263607,4.4861584,4.7126136,4.939069,4.8765984,4.814128,4.7516575,4.689187,4.6267166,4.6110992,4.5993857,4.5876727,4.575959,4.564246,4.337791,4.1113358,3.8887846,3.6623292,3.435874,3.174279,2.912684,2.6510892,2.3855898,2.1239948,2.174752,2.2255092,2.2762666,2.3231194,2.3738766,2.1981785,2.0263848,1.8506867,1.6749885,1.4992905,1.475864,1.4485333,1.4251068,1.4016805,1.3743496,1.3001659,1.2259823,1.1517987,1.0737107,0.999527,0.97610056,0.94876975,0.92534333,0.9019169,0.8745861,0.76135844,0.6481308,0.5388075,0.42557985,0.31235218,0.37482262,0.43729305,0.4997635,0.5622339,0.62470436,0.6481308,0.6754616,0.698888,0.7262188,0.74964523,0.6871748,0.62470436,0.5622339,0.4997635,0.43729305,0.7262188,1.0112402,1.3001659,1.5890918,1.8741131,1.5500476,1.2259823,0.9019169,0.57394713,0.24988174,0.3513962,0.44900626,0.5505207,0.6481308,0.74964523,0.80040246,0.8511597,0.9019169,0.94876975,0.999527,1.5734742,2.1513257,2.7252727,3.2992198,3.873167,3.1000953,2.3231194,1.5500476,0.77307165,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.57394713,1.0268579,1.475864,1.9248703,2.3738766,2.8385005,3.2992198,3.7638438,4.224563,4.689187,5.001539,5.3138914,5.6262436,5.938596,6.250948,5.4388323,4.6267166,3.8106966,2.998581,2.1864653,3.4514916,4.7126136,5.9737353,7.238762,8.499884,8.773191,9.050405,9.323712,9.600925,9.874233,8.862993,7.8517528,6.8366084,5.825368,4.814128,5.138193,5.462259,5.786324,6.114294,6.4383593,5.786324,5.138193,4.4861584,3.8380275,3.1859922,3.1391394,3.0883822,3.0376248,2.9868677,2.9361105,2.8111696,2.6862288,2.5612879,2.436347,2.3114061,1.8506867,1.3860629,0.92534333,0.46071947,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.1639849,0.19912452,0.23816854,0.27330816,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.6481308,0.9878138,1.3235924,1.6632754,1.999054,2.35045,2.7018464,3.049338,3.4007344,3.7482262,3.6623292,3.5764325,3.4866312,3.4007344,3.310933,3.873167,4.4393053,5.001539,5.563773,6.126007,6.5008297,6.8756523,7.250475,7.6252975,8.00012,7.9259367,7.8517528,7.773665,7.699481,7.6252975,8.125061,8.624825,9.124588,9.6243515,10.124115,10.573121,11.0260315,11.475039,11.924045,12.373051,11.763964,11.150972,10.537982,9.924991,9.311999,10.299813,11.287627,12.27544,13.263254,14.251068,13.036799,11.826434,10.612165,9.4018,8.187531,7.6643414,7.137247,6.6140575,6.086963,5.563773,5.473972,5.388075,5.298274,5.212377,5.12648,5.5130157,5.899552,6.2860875,6.676528,7.0630636,6.012779,4.9624953,3.912211,2.8619268,1.8116426,1.5890918,1.3626363,1.1361811,0.9136301,0.6871748,0.737932,0.78868926,0.8394465,0.8862993,0.93705654,0.26159495,0.28111696,0.30063897,0.3240654,0.3435874,0.3631094,0.42948425,0.4958591,0.5661383,0.63251317,0.698888,0.59737355,0.4958591,0.39434463,0.28892577,0.18741131,0.21474212,0.24207294,0.26940376,0.29673457,0.3240654,0.46462387,0.60518235,0.74574083,0.8862993,1.0268579,0.92924774,0.8355421,0.7418364,0.6442264,0.5505207,0.4997635,0.44900626,0.39824903,0.3513962,0.30063897,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.113227665,0.1756981,0.23816854,0.30063897,0.3631094,0.42557985,0.49195468,0.5583295,0.62079996,0.6871748,0.81211567,0.93705654,1.0619974,1.1869383,1.3118792,1.0854238,0.8589685,0.62860876,0.40215343,0.1756981,0.1835069,0.19522011,0.20693332,0.21474212,0.22645533,0.21474212,0.20693332,0.19522011,0.1835069,0.1756981,0.15227169,0.12884527,0.10932326,0.08589685,0.062470436,0.113227665,0.1639849,0.21083772,0.26159495,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.08589685,0.10932326,0.12884527,0.15227169,0.1756981,0.1756981,0.1756981,0.1756981,0.1756981,0.1756981,0.20693332,0.23426414,0.26549935,0.29673457,0.3240654,0.359205,0.39434463,0.42948425,0.46462387,0.4997635,0.40996224,0.32016098,0.23035973,0.14055848,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.08980125,0.093705654,0.093705654,0.09761006,0.10151446,0.10932326,0.12103647,0.12884527,0.14055848,0.14836729,0.18741131,0.22645533,0.26159495,0.30063897,0.3357786,0.44510186,0.5544251,0.659844,0.76916724,0.8745861,0.97219616,1.0698062,1.1674163,1.2650263,1.3626363,1.475864,1.5890918,1.698415,1.8116426,1.9248703,1.901444,1.8819219,1.8584955,1.8350691,1.8116426,1.7882162,1.7686942,1.7452679,1.7218413,1.698415,1.9092526,2.1161861,2.3231194,2.5300527,2.736986,3.2836022,3.8341231,4.380739,4.927356,5.473972,5.2006636,4.93126,4.657952,4.3846436,4.1113358,3.9902992,3.8692627,3.7443218,3.6232853,3.4983444,3.39683,3.2953155,3.193801,3.0883822,2.9868677,3.06886,3.1469483,3.2289407,3.3070288,3.3890212,3.5959544,3.8067923,4.01763,4.2284675,4.4393053,4.5447245,4.6540475,4.759466,4.8687897,4.9742084,4.7126136,4.4510183,4.1894236,3.9239242,3.6623292,4.661856,5.661383,6.66091,7.6643414,8.663869,8.296855,7.9337454,7.5667315,7.2036223,6.8366084,6.8951745,6.9537406,7.008402,7.066968,7.125534,8.921559,10.721489,12.517513,14.313539,16.113468,15.418485,14.727406,14.036326,13.341343,12.650263,12.892336,13.134409,13.376482,13.618555,13.860628,14.989,16.113468,17.237936,18.362404,19.486872,16.238409,12.993851,9.745388,6.4969254,3.2484627,2.6003318,1.9482968,1.3001659,0.6481308,0.0,0.0,0.0,0.0,0.0,0.0,0.6520352,1.3040704,1.9561055,2.6081407,3.2640803,2.9868677,2.7135596,2.436347,2.1630387,1.8858263,2.1396124,2.3933985,2.6432803,2.8970666,3.1508527,2.697942,2.2450314,1.7921207,1.33921,0.8862993,0.7106012,0.5309987,0.3553006,0.1756981,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.42948425,0.8589685,1.2884527,1.7218413,2.1513257,2.77603,3.4007344,4.025439,4.650143,5.2748475,4.630621,3.9902992,3.3460727,2.7057507,2.0615244,5.610626,9.155824,12.704925,16.254026,19.799223,16.909966,14.020708,11.131451,8.238289,5.349031,5.4505453,5.548156,5.64967,5.7511845,5.8487945,5.840986,5.833177,5.8292727,5.8214636,5.813655,5.3724575,4.93126,4.493967,4.0527697,3.611572,3.6701381,3.7287042,3.7833657,3.8419318,3.900498,4.0137253,4.1308575,4.2440853,4.3612175,4.474445,4.365122,4.2557983,4.1464753,4.0332475,3.9239242,3.9434462,3.959064,3.978586,3.9942036,4.0137253,3.951255,3.8887846,3.8263142,3.7638438,3.7013733,3.4514916,3.2016098,2.951728,2.7018464,2.4480603,2.463678,2.475391,2.4871042,2.4988174,2.514435,2.4285383,2.3426414,2.2567444,2.1708477,2.0888553,1.9639144,1.8389735,1.7140326,1.5890918,1.4641509,1.4212024,1.3782539,1.3353056,1.2923572,1.2494087,1.1713207,1.0932326,1.0190489,0.94096094,0.8628729,0.8160201,0.76916724,0.71841,0.6715572,0.62470436,0.6559396,0.6910792,0.7223144,0.75354964,0.78868926,0.78088045,0.77307165,0.76526284,0.75745404,0.74964523,0.7418364,0.7301232,0.71841,0.7106012,0.698888,0.92534333,1.1517987,1.3743496,1.6008049,1.8233559,1.6125181,1.4016805,1.1869383,0.97610056,0.76135844,0.76916724,0.77307165,0.77697605,0.78088045,0.78868926,0.96048295,1.1322767,1.3040704,1.475864,1.6515622,1.999054,2.3465457,2.6940374,3.0415294,3.3890212,2.87364,2.358259,1.8428779,1.3274968,0.81211567,0.679366,0.5466163,0.41386664,0.28111696,0.14836729,0.4997635,0.8511597,1.1986516,1.5500476,1.901444,2.3933985,2.8892577,3.3851168,3.8809757,4.376835,4.6228123,4.8687897,5.1186714,5.364649,5.610626,5.0132523,4.415879,3.8185053,3.2211318,2.6237583,3.7716527,4.9156423,6.0596323,7.2036223,8.351517,8.632633,8.913751,9.198771,9.479889,9.761005,8.976221,8.187531,7.3988423,6.6140575,5.825368,5.813655,5.801942,5.786324,5.774611,5.7628975,5.2045684,4.646239,4.0918136,3.533484,2.9751544,2.9673457,2.959537,2.951728,2.9439192,2.9361105,2.8463092,2.7565079,2.6667068,2.5769055,2.4871042,1.9912452,1.4914817,0.9956226,0.4958591,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,0.32016098,0.23816854,0.16008049,0.078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.23816854,0.29283017,0.3435874,0.39824903,0.44900626,0.42557985,0.40605783,0.38263142,0.359205,0.3357786,0.27721256,0.21864653,0.15617609,0.09761006,0.039044023,0.078088045,0.12103647,0.1639849,0.20693332,0.24988174,0.5309987,0.8160201,1.097137,1.3782539,1.6632754,1.9756275,2.2879796,2.6003318,2.912684,3.2250361,3.2211318,3.213323,3.2094188,3.2055142,3.2016098,3.619381,4.0332475,4.4510183,4.8687897,5.2865605,5.716045,6.141625,6.571109,6.996689,7.426173,7.3597984,7.2934237,7.230953,7.164578,7.098203,7.5862536,8.070399,8.554545,9.0386915,9.526741,10.073358,10.619974,11.166591,11.713207,12.263727,11.639023,11.014318,10.38571,9.761005,9.136301,10.073358,11.00651,11.943566,12.8767185,13.813775,12.619028,11.428185,10.2334385,9.042596,7.8517528,7.355894,6.860035,6.364176,5.8683167,5.376362,5.22409,5.0757227,4.9234514,4.775084,4.6267166,4.911738,5.2006636,5.4856853,5.774611,6.0635366,5.138193,4.2167544,3.2953155,2.3738766,1.4485333,1.2689307,1.0893283,0.9097257,0.7301232,0.5505207,0.6481308,0.74574083,0.8433509,0.94096094,1.038571,0.3357786,0.339683,0.3435874,0.3435874,0.3474918,0.3513962,0.39824903,0.44510186,0.49195468,0.5388075,0.58566034,0.5075723,0.42557985,0.3474918,0.26940376,0.18741131,0.21864653,0.24597734,0.27721256,0.30844778,0.3357786,0.44119745,0.5466163,0.6520352,0.75745404,0.8628729,0.78478485,0.7066968,0.62860876,0.5544251,0.47633708,0.46071947,0.44900626,0.43729305,0.42557985,0.41386664,0.3513962,0.28892577,0.22645533,0.1639849,0.10151446,0.1639849,0.22645533,0.28892577,0.3513962,0.41386664,0.49195468,0.57394713,0.6520352,0.7340276,0.81211567,0.8628729,0.9136301,0.96438736,1.0112402,1.0619974,0.8941081,0.7262188,0.5583295,0.39434463,0.22645533,0.25769055,0.28892577,0.3240654,0.3553006,0.38653582,0.37872702,0.3709182,0.3631094,0.359205,0.3513962,0.29283017,0.23426414,0.1756981,0.12103647,0.062470436,0.10151446,0.13665408,0.1756981,0.21083772,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,0.08199245,0.10151446,0.12103647,0.14055848,0.1639849,0.1639849,0.1639849,0.1639849,0.1639849,0.1639849,0.21083772,0.25769055,0.30454338,0.3513962,0.39824903,0.42167544,0.44119745,0.46071947,0.48024148,0.4997635,0.40605783,0.31625658,0.22255093,0.12884527,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.10541886,0.09761006,0.08980125,0.08199245,0.07418364,0.08199245,0.08980125,0.09761006,0.10541886,0.113227665,0.14836729,0.18741131,0.22645533,0.26159495,0.30063897,0.44119745,0.58175594,0.71841,0.8589685,0.999527,1.0698062,1.1400855,1.2103647,1.2806439,1.3509232,1.4485333,1.5500476,1.6515622,1.7491722,1.8506867,1.8428779,1.8350691,1.8272603,1.8194515,1.8116426,1.8038338,1.796025,1.7882162,1.7843118,1.7765031,2.0146716,2.2567444,2.494913,2.7330816,2.9751544,3.4436827,3.9161155,4.3846436,4.853172,5.3256044,5.067914,4.8102236,4.552533,4.2948427,4.037152,3.9161155,3.7989833,3.677947,3.5569105,3.435874,3.3460727,3.252367,3.1586614,3.06886,2.9751544,3.0337205,3.096191,3.154757,3.213323,3.2757936,3.6584249,4.041056,4.423688,4.806319,5.1889505,5.114767,5.040583,4.970304,4.8961205,4.825841,4.5993857,4.376835,4.1503797,3.9239242,3.7013733,4.9742084,6.250948,7.523783,8.800523,10.073358,9.280765,8.488171,7.6955767,6.9068875,6.114294,6.453977,6.79366,7.1333427,7.473026,7.812709,9.682918,11.553126,13.423335,15.293544,17.163752,16.254026,15.344301,14.430671,13.520945,12.611219,13.021181,13.431144,13.841106,14.251068,14.661031,15.324779,15.988527,16.64837,17.31212,17.975868,15.055375,12.134882,9.21439,6.2938967,3.3734035,2.7018464,2.0263848,1.3509232,0.6754616,0.0,0.0,0.0,0.0,0.0,0.0,0.8433509,1.6867018,2.5261483,3.3694992,4.21285,4.126953,4.037152,3.951255,3.8614538,3.775557,3.6545205,3.533484,3.416352,3.2953155,3.174279,2.7565079,2.338737,1.9209659,1.5031948,1.0893283,0.8706817,0.6520352,0.43338865,0.21864653,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3240654,0.6442264,0.96829176,1.2884527,1.6125181,2.5261483,3.435874,4.349504,5.263134,6.1767645,5.466163,4.755562,4.044961,3.3343596,2.6237583,5.1186714,7.6135845,10.108498,12.603411,15.098324,13.044608,10.990892,8.933272,6.8795567,4.825841,4.939069,5.0483923,5.1616197,5.2748475,5.388075,5.3217,5.2592297,5.192855,5.12648,5.0640097,4.743849,4.4275923,4.1113358,3.7911747,3.474918,3.5764325,3.6818514,3.7833657,3.8848803,3.9863946,3.9942036,3.998108,4.0020123,4.0059166,4.0137253,3.853645,3.697469,3.541293,3.3812122,3.2250361,3.2718892,3.3187418,3.3655949,3.416352,3.4632049,3.5608149,3.6623292,3.7638438,3.8614538,3.9629683,3.7247996,3.4866312,3.2484627,3.0141985,2.77603,2.7486992,2.7252727,2.7018464,2.6745155,2.6510892,2.6549935,2.6588979,2.6667068,2.6706111,2.6745155,2.4480603,2.2255092,1.999054,1.7765031,1.5500476,1.5383345,1.5305257,1.5188124,1.5110037,1.4992905,1.3704453,1.2415999,1.1088502,0.98000497,0.8511597,0.8667773,0.8862993,0.9019169,0.92143893,0.93705654,0.94096094,0.94096094,0.94486535,0.94876975,0.94876975,0.9097257,0.8706817,0.8316377,0.78868926,0.74964523,0.79259366,0.8355421,0.8784905,0.92143893,0.96438736,1.1244678,1.2884527,1.4485333,1.6125181,1.7765031,1.6749885,1.5734742,1.475864,1.3743496,1.2767396,1.1869383,1.0932326,1.0034313,0.9136301,0.8238289,1.1205635,1.4133936,1.7101282,2.0068626,2.2996929,2.4207294,2.541766,2.6588979,2.7799344,2.900971,2.6432803,2.3894942,2.135708,1.8819219,1.6242313,1.3353056,1.0463798,0.75354964,0.46462387,0.1756981,0.42557985,0.6754616,0.92534333,1.175225,1.4251068,1.9522011,2.4792955,3.0063896,3.533484,4.0605783,4.2440853,4.4275923,4.6110992,4.7907014,4.9742084,4.591577,4.2089458,3.8263142,3.4436827,3.0610514,4.0918136,5.1186714,6.1455293,7.172387,8.1992445,8.488171,8.781001,9.069926,9.358852,9.651682,9.085544,8.52331,7.9610763,7.3988423,6.8366084,6.4891167,6.13772,5.786324,5.4388323,5.087436,4.6228123,4.1581883,3.6935644,3.2289407,2.7643168,2.795552,2.8306916,2.8658314,2.900971,2.9361105,2.8814487,2.8267872,2.7721257,2.717464,2.6628022,2.1318035,1.5969005,1.0659018,0.5309987,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.31625658,0.38653582,0.45291066,0.5192855,0.58566034,0.59346914,0.59737355,0.60127795,0.60908675,0.61299115,0.5036679,0.39824903,0.28892577,0.1835069,0.07418364,0.09761006,0.12103647,0.14055848,0.1639849,0.18741131,0.41386664,0.6442264,0.8706817,1.097137,1.3235924,1.6008049,1.8741131,2.1513257,2.4246337,2.7018464,2.77603,2.854118,2.9322062,3.0102942,3.0883822,3.3616903,3.631094,3.9044023,4.1777105,4.4510183,4.93126,5.4115014,5.891743,6.36808,6.8483214,6.79366,6.7389984,6.6843367,6.629675,6.575013,7.043542,7.5159745,7.984503,8.453031,8.925464,9.56969,10.213917,10.858143,11.506273,12.150499,11.514082,10.87376,10.237343,9.600925,8.960603,9.846903,10.729298,11.611692,12.494087,13.376482,12.201257,11.029937,9.858616,8.683391,7.5120697,7.0474463,6.5828223,6.1181984,5.6535745,5.1889505,4.9742084,4.7633705,4.548629,4.337791,4.123049,4.3143644,4.5017757,4.689187,4.8765984,5.0640097,4.267512,3.4710135,2.67842,1.8819219,1.0893283,0.95267415,0.8160201,0.6832704,0.5466163,0.41386664,0.5583295,0.7027924,0.8472553,0.9917182,1.1361811,0.41386664,0.39824903,0.38263142,0.3670138,0.3513962,0.3357786,0.3631094,0.39434463,0.42167544,0.44900626,0.47633708,0.41777104,0.359205,0.30063897,0.24597734,0.18741131,0.21864653,0.25378615,0.28502136,0.31625658,0.3513962,0.42167544,0.48805028,0.5583295,0.62860876,0.698888,0.64032197,0.58175594,0.5192855,0.46071947,0.39824903,0.42557985,0.44900626,0.47633708,0.4997635,0.5231899,0.44900626,0.37482262,0.30063897,0.22645533,0.14836729,0.21083772,0.27330816,0.3357786,0.39824903,0.46071947,0.5583295,0.6520352,0.74574083,0.8433509,0.93705654,0.9136301,0.8862993,0.8628729,0.8394465,0.81211567,0.7066968,0.59737355,0.48805028,0.38263142,0.27330816,0.3318742,0.38653582,0.44119745,0.4958591,0.5505207,0.5466163,0.5388075,0.5349031,0.5309987,0.5231899,0.43338865,0.339683,0.24597734,0.15617609,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.078088045,0.09761006,0.113227665,0.13274968,0.14836729,0.14836729,0.14836729,0.14836729,0.14836729,0.14836729,0.21474212,0.28111696,0.3435874,0.40996224,0.47633708,0.48024148,0.48414588,0.48805028,0.4958591,0.4997635,0.40605783,0.30844778,0.21474212,0.12103647,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.12103647,0.10151446,0.08589685,0.06637484,0.05075723,0.05466163,0.058566034,0.06637484,0.07027924,0.07418364,0.113227665,0.14836729,0.18741131,0.22645533,0.26159495,0.43338865,0.60908675,0.78088045,0.95267415,1.1244678,1.1674163,1.2103647,1.2533131,1.2962615,1.33921,1.4251068,1.5110037,1.6008049,1.6867018,1.7765031,1.7843118,1.7882162,1.796025,1.8038338,1.8116426,1.8194515,1.8272603,1.8350691,1.8428779,1.8506867,2.1239948,2.3933985,2.6667068,2.9400148,3.213323,3.6037633,3.998108,4.388548,4.7828927,5.173333,4.93126,4.689187,4.447114,4.2050414,3.9629683,3.8458362,3.7287042,3.611572,3.49444,3.3734035,3.2914112,3.2094188,3.1274261,3.0454338,2.9634414,3.0024853,3.0415294,3.0805733,3.1235218,3.1625657,3.716991,4.271416,4.825841,5.3841705,5.938596,5.6848097,5.4310236,5.181142,4.927356,4.6735697,4.4861584,4.298747,4.1113358,3.9239242,3.736513,5.2865605,6.8366084,8.386656,9.936704,11.486752,10.268578,9.0465,7.8283267,6.606249,5.388075,6.008875,6.6335793,7.2543793,7.8790836,8.499884,10.444276,12.384764,14.329156,16.269644,18.214037,17.085665,15.957292,14.828919,13.700547,12.576079,13.153932,13.731783,14.30573,14.883581,15.461433,15.660558,15.863586,16.062712,16.261835,16.46096,13.868437,11.275913,8.683391,6.0908675,3.4983444,2.7994564,2.1005683,1.4016805,0.698888,0.0,0.0,0.0,0.0,0.0,0.0,1.0307622,2.0654287,3.096191,4.1308575,5.1616197,5.263134,5.3607445,5.462259,5.563773,5.661383,5.169429,4.677474,4.185519,3.6935644,3.2016098,2.8189783,2.436347,2.0537157,1.6710842,1.2884527,1.0307622,0.77307165,0.5153811,0.25769055,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21474212,0.42948425,0.6442264,0.8589685,1.0737107,2.2762666,3.474918,4.6735697,5.8761253,7.0747766,6.297801,5.520825,4.743849,3.9668727,3.1859922,4.630621,6.0713453,7.5159745,8.956698,10.401327,9.17925,7.9610763,6.7389984,5.520825,4.298747,4.423688,4.548629,4.6735697,4.7985106,4.9234514,4.802415,4.6813784,4.5564375,4.435401,4.3143644,4.1191444,3.9239242,3.7287042,3.533484,3.338264,3.4866312,3.631094,3.7794614,3.9278288,4.0761957,3.970777,3.8653584,3.7599394,3.6545205,3.5491016,3.3460727,3.1391394,2.9361105,2.7291772,2.5261483,2.6042364,2.67842,2.7565079,2.8345962,2.912684,3.174279,3.435874,3.7013733,3.9629683,4.224563,3.998108,3.775557,3.5491016,3.3265507,3.1000953,3.0376248,2.9751544,2.912684,2.8502135,2.787743,2.8814487,2.979059,3.0727646,3.1664703,3.2640803,2.9361105,2.612045,2.2879796,1.9639144,1.6359446,1.6593709,1.6827974,1.7062237,1.7257458,1.7491722,1.5656652,1.3860629,1.2025559,1.0190489,0.8394465,0.92143893,1.0034313,1.0854238,1.1674163,1.2494087,1.2220778,1.1947471,1.1674163,1.1400855,1.1127546,1.038571,0.96829176,0.8941081,0.8238289,0.74964523,0.8433509,0.94096094,1.0346665,1.1283722,1.2259823,1.3235924,1.4251068,1.5266213,1.6242313,1.7257458,1.737459,1.7491722,1.7608855,1.7765031,1.7882162,1.6008049,1.4172981,1.2337911,1.0463798,0.8628729,1.2806439,1.698415,2.1161861,2.533957,2.951728,2.8424048,2.7330816,2.6276627,2.5183394,2.4129205,2.416825,2.4207294,2.4285383,2.4324427,2.436347,1.9912452,1.542239,1.0932326,0.6481308,0.19912452,0.3513962,0.4997635,0.6481308,0.80040246,0.94876975,1.5110037,2.069333,2.631567,3.1898966,3.7482262,3.8692627,3.9863946,4.1035266,4.220659,4.337791,4.169902,4.0020123,3.8341231,3.6662338,3.4983444,4.4119744,5.3217,6.2314262,7.141152,8.050878,8.347612,8.644346,8.941081,9.24172,9.538455,9.198771,8.862993,8.52331,8.187531,7.8517528,7.1606736,6.473499,5.786324,5.099149,4.4119744,4.041056,3.6662338,3.2953155,2.9243972,2.5495746,2.6276627,2.7057507,2.7838387,2.8619268,2.9361105,2.9165885,2.8970666,2.8775444,2.8580225,2.8385005,2.2684577,1.7023194,1.1361811,0.5661383,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.39434463,0.47633708,0.5583295,0.6442264,0.7262188,0.75745404,0.78868926,0.8238289,0.8550641,0.8862993,0.7340276,0.57785153,0.42167544,0.26940376,0.113227665,0.113227665,0.11713207,0.12103647,0.12103647,0.12494087,0.29673457,0.46852827,0.6442264,0.8160201,0.9878138,1.2259823,1.4641509,1.698415,1.9365835,2.174752,2.3348327,2.494913,2.6549935,2.815074,2.9751544,3.1039999,3.2289407,3.357786,3.4866312,3.611572,4.1464753,4.677474,5.2084727,5.743376,6.2743745,6.2314262,6.184573,6.141625,6.094772,6.0518236,6.504734,6.9615493,7.4144597,7.871275,8.324185,9.066022,9.811763,10.553599,11.295436,12.037272,11.389141,10.737106,10.088976,9.43694,8.78881,9.616543,10.44818,11.275913,12.107552,12.939189,11.783486,10.631687,9.479889,8.32809,7.1762915,6.7389984,6.3056097,5.8683167,5.434928,5.001539,4.7243266,4.4510183,4.173806,3.900498,3.6232853,3.7130866,3.7989833,3.8887846,3.9746814,4.0605783,3.39683,2.7291772,2.0615244,1.3938715,0.7262188,0.63641757,0.5466163,0.45681506,0.3631094,0.27330816,0.46852827,0.659844,0.8511597,1.0463798,1.2376955,0.48805028,0.45681506,0.42167544,0.39044023,0.359205,0.3240654,0.3318742,0.339683,0.3474918,0.3553006,0.3631094,0.3279698,0.29283017,0.25769055,0.22255093,0.18741131,0.22255093,0.25769055,0.29283017,0.3279698,0.3631094,0.39824903,0.43338865,0.46852827,0.5036679,0.5388075,0.4958591,0.45291066,0.40996224,0.3670138,0.3240654,0.38653582,0.44900626,0.5114767,0.57394713,0.63641757,0.5505207,0.46071947,0.37482262,0.28892577,0.19912452,0.26159495,0.3240654,0.38653582,0.44900626,0.5114767,0.62079996,0.7340276,0.8433509,0.95267415,1.0619974,0.96438736,0.8628729,0.76135844,0.6637484,0.5622339,0.5153811,0.46852827,0.42167544,0.3709182,0.3240654,0.40215343,0.48024148,0.5583295,0.63641757,0.7106012,0.7106012,0.7066968,0.7066968,0.7027924,0.698888,0.57394713,0.44510186,0.31625658,0.19131571,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.078088045,0.093705654,0.10932326,0.12103647,0.13665408,0.13665408,0.13665408,0.13665408,0.13665408,0.13665408,0.21864653,0.30063897,0.38653582,0.46852827,0.5505207,0.5388075,0.5309987,0.5192855,0.5114767,0.4997635,0.40215343,0.30454338,0.20693332,0.10932326,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.031235218,0.06637484,0.09761006,0.12884527,0.1639849,0.13665408,0.10932326,0.078088045,0.05075723,0.023426414,0.027330816,0.031235218,0.031235218,0.03513962,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.22645533,0.42948425,0.63641757,0.8394465,1.0463798,1.2494087,1.2650263,1.2806439,1.2962615,1.3118792,1.3235924,1.4016805,1.475864,1.5500476,1.6242313,1.698415,1.7218413,1.7452679,1.7686942,1.7882162,1.8116426,1.8350691,1.8584955,1.8819219,1.901444,1.9248703,2.2294137,2.533957,2.8385005,3.1469483,3.4514916,3.7638438,4.0801005,4.396357,4.7087092,5.024966,4.7985106,4.5681505,4.3416953,4.11524,3.8887846,3.7716527,3.6584249,3.541293,3.4280653,3.310933,3.240654,3.1664703,3.096191,3.0220075,2.951728,2.97125,2.9907722,3.0102942,3.0298162,3.049338,3.775557,4.50568,5.2318993,5.958118,6.688241,6.2548523,5.8214636,5.388075,4.958591,4.5252023,4.376835,4.224563,4.0761957,3.9239242,3.775557,5.5989127,7.426173,9.249529,11.076789,12.900145,11.252487,9.60483,7.957172,6.309514,4.661856,5.5676775,6.473499,7.37932,8.281238,9.187058,11.20173,13.216402,15.231073,17.245745,19.26432,17.917301,16.574188,15.227169,13.884054,12.537036,13.282777,14.028518,14.774258,15.516094,16.261835,16.00024,15.738646,15.473146,15.211552,14.949956,12.685403,10.42085,8.156297,5.891743,3.6232853,2.900971,2.174752,1.4485333,0.7262188,0.0,0.0,0.0,0.0,0.0,0.0,1.2220778,2.4441557,3.6662338,4.8883114,6.114294,6.3993154,6.688241,6.9732623,7.262188,7.551114,6.6843367,5.8214636,4.9546866,4.0918136,3.2250361,2.8775444,2.5300527,2.182561,1.8350691,1.4875772,1.1908426,0.8941081,0.59346914,0.29673457,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10932326,0.21474212,0.3240654,0.42948425,0.5388075,2.0263848,3.513962,5.001539,6.4891167,7.9766936,7.1294384,6.2860875,5.4388323,4.5954814,3.7482262,4.138666,4.5291066,4.919547,5.309987,5.700427,5.3138914,4.93126,4.5447245,4.1581883,3.775557,3.912211,4.0488653,4.1894236,4.3260775,4.462732,4.283129,4.1035266,3.9239242,3.7443218,3.5608149,3.4905357,3.416352,3.3460727,3.2718892,3.2016098,3.3929255,3.5842414,3.775557,3.970777,4.1620927,3.9473507,3.7326086,3.5178664,3.3031244,3.0883822,2.8345962,2.5808098,2.330928,2.077142,1.8233559,1.9326792,2.0380979,2.1474214,2.2567444,2.3621633,2.787743,3.213323,3.638903,4.0605783,4.4861584,4.2753205,4.0605783,3.8497405,3.638903,3.4241607,3.3265507,3.2250361,3.1235218,3.0259118,2.9243972,3.1118085,3.2953155,3.4788225,3.6662338,3.8497405,3.4241607,2.998581,2.5769055,2.1513257,1.7257458,1.7804074,1.8350691,1.8897307,1.9443923,1.999054,1.7647898,1.5305257,1.2962615,1.0580931,0.8238289,0.97219616,1.1205635,1.2689307,1.4133936,1.5617609,1.5031948,1.4485333,1.3899672,1.3314011,1.2767396,1.1713207,1.0659018,0.96048295,0.8550641,0.74964523,0.8980125,1.0463798,1.1908426,1.33921,1.4875772,1.5266213,1.5617609,1.6008049,1.6359446,1.6749885,1.7999294,1.9248703,2.0498111,2.174752,2.2996929,2.018576,1.7413634,1.4602464,1.1791295,0.9019169,1.4407244,1.979532,2.5183394,3.0610514,3.5998588,3.2640803,2.9283018,2.5964274,2.260649,1.9248703,2.1903696,2.455869,2.7213683,2.9868677,3.2484627,2.6432803,2.0380979,1.43682,0.8316377,0.22645533,0.27330816,0.3240654,0.37482262,0.42557985,0.47633708,1.0659018,1.6593709,2.25284,2.8463092,3.435874,3.4905357,3.541293,3.5959544,3.6467118,3.7013733,3.7482262,3.795079,3.8419318,3.8887846,3.9356375,4.728231,5.520825,6.3134184,7.1060123,7.898606,8.203149,8.511597,8.81614,9.120684,9.425227,9.311999,9.198771,9.085544,8.976221,8.862993,7.8361354,6.813182,5.786324,4.7633705,3.736513,3.4593005,3.1781836,2.8970666,2.6159496,2.338737,2.455869,2.5769055,2.697942,2.8189783,2.9361105,2.951728,2.9673457,2.9829633,2.998581,3.0141985,2.4090161,1.8077383,1.2064602,0.60127795,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.47243267,0.5700427,0.6676528,0.76526284,0.8628729,0.92143893,0.98390937,1.0424755,1.1010414,1.1635119,0.96048295,0.75745404,0.5544251,0.3513962,0.14836729,0.13274968,0.113227665,0.09761006,0.078088045,0.062470436,0.1796025,0.29673457,0.41386664,0.5309987,0.6481308,0.8511597,1.0502841,1.2494087,1.4485333,1.6515622,1.893635,2.135708,2.377781,2.619854,2.8619268,2.8463092,2.8267872,2.8111696,2.7916477,2.77603,3.3616903,3.9434462,4.5291066,5.114767,5.700427,5.6652875,5.630148,5.5950084,5.559869,5.5247293,5.9659266,6.4032197,6.844417,7.2856145,7.726812,8.566258,9.405705,10.2451515,11.084598,11.924045,11.2642,10.600452,9.936704,9.276859,8.6131115,9.390087,10.167064,10.944039,11.721016,12.501896,11.365715,10.2334385,9.101162,7.968885,6.8366084,6.4305506,6.028397,5.6223392,5.2162814,4.814128,4.474445,4.138666,3.7989833,3.4632049,3.1235218,3.1118085,3.1000953,3.0883822,3.076669,3.0610514,2.522244,1.9834363,1.4407244,0.9019169,0.3631094,0.31625658,0.27330816,0.22645533,0.1835069,0.13665408,0.37872702,0.61689556,0.8589685,1.097137,1.33921,0.5622339,0.5114767,0.46071947,0.41386664,0.3631094,0.31235218,0.30063897,0.28892577,0.27330816,0.26159495,0.24988174,0.23816854,0.22645533,0.21083772,0.19912452,0.18741131,0.22645533,0.26159495,0.30063897,0.3357786,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.3513962,0.3240654,0.30063897,0.27330816,0.24988174,0.3513962,0.44900626,0.5505207,0.6481308,0.74964523,0.6481308,0.5505207,0.44900626,0.3513962,0.24988174,0.31235218,0.37482262,0.43729305,0.4997635,0.5622339,0.6871748,0.81211567,0.93705654,1.0619974,1.1869383,1.0112402,0.8394465,0.6637484,0.48805028,0.31235218,0.3240654,0.3357786,0.3513962,0.3631094,0.37482262,0.47633708,0.57394713,0.6754616,0.77307165,0.8745861,0.8745861,0.8745861,0.8745861,0.8745861,0.8745861,0.7106012,0.5505207,0.38653582,0.22645533,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.22645533,0.3240654,0.42557985,0.5231899,0.62470436,0.60127795,0.57394713,0.5505207,0.5231899,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.42557985,0.6637484,0.9019169,1.1361811,1.3743496,1.3626363,1.3509232,1.33921,1.3235924,1.3118792,1.3743496,1.43682,1.4992905,1.5617609,1.6242313,1.6632754,1.698415,1.737459,1.7765031,1.8116426,1.8506867,1.8858263,1.9248703,1.9639144,1.999054,2.338737,2.6745155,3.0141985,3.349977,3.6857557,3.9239242,4.1620927,4.4002614,4.6384296,4.8765984,4.661856,4.4510183,4.2362766,4.025439,3.8106966,3.7013733,3.5881457,3.474918,3.3616903,3.2484627,3.1859922,3.1235218,3.0610514,2.998581,2.9361105,2.9361105,2.9361105,2.9361105,2.9361105,2.9361105,3.8380275,4.73604,5.6379566,6.5359693,7.437886,6.824895,6.211904,5.5989127,4.985922,4.376835,4.263607,4.1503797,4.037152,3.9239242,3.8106966,5.911265,8.011833,10.112402,12.212971,14.313539,12.236397,10.163159,8.086017,6.012779,3.9356375,5.12648,6.3134184,7.5003567,8.687295,9.874233,11.963089,14.048039,16.136894,18.22575,20.310701,18.74894,17.18718,15.625418,14.063657,12.501896,13.411622,14.325252,15.238882,16.148607,17.062239,16.33602,15.613705,14.8874855,14.161267,13.438952,11.498465,9.561881,7.6252975,5.688714,3.7482262,2.998581,2.2489357,1.4992905,0.74964523,0.0,0.0,0.0,0.0,0.0,0.0,1.4133936,2.8267872,4.2362766,5.64967,7.0630636,7.5394006,8.011833,8.488171,8.960603,9.43694,8.1992445,6.9615493,5.7238536,4.4861584,3.2484627,2.9361105,2.6237583,2.3114061,1.999054,1.6867018,1.3509232,1.0112402,0.6754616,0.3357786,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.7765031,3.5491016,5.3256044,7.098203,8.874706,7.9610763,7.0513506,6.13772,5.22409,4.3143644,3.6506162,2.9868677,2.3231194,1.6632754,0.999527,1.4485333,1.901444,2.35045,2.7994564,3.2484627,3.4007344,3.5491016,3.7013733,3.8497405,3.998108,3.7638438,3.5256753,3.2875066,3.049338,2.8111696,2.8619268,2.912684,2.9634414,3.0141985,3.0610514,3.2992198,3.5373883,3.775557,4.0137253,4.251894,3.9239242,3.5998588,3.2757936,2.951728,2.6237583,2.3231194,2.0263848,1.7257458,1.4251068,1.1244678,1.261122,1.4016805,1.5383345,1.6749885,1.8116426,2.4012074,2.9868677,3.5764325,4.1620927,4.7516575,4.548629,4.349504,4.1503797,3.951255,3.7482262,3.611572,3.474918,3.338264,3.2016098,3.0610514,3.338264,3.611572,3.8887846,4.1620927,4.4393053,3.912211,3.3890212,2.8619268,2.338737,1.8116426,1.901444,1.9873407,2.0732377,2.1630387,2.2489357,1.9639144,1.6749885,1.3860629,1.1010414,0.81211567,1.0268579,1.2376955,1.4485333,1.6632754,1.8741131,1.7882162,1.698415,1.6125181,1.5266213,1.43682,1.3001659,1.1635119,1.0268579,0.8862993,0.74964523,0.94876975,1.1517987,1.3509232,1.5500476,1.7491722,1.7257458,1.698415,1.6749885,1.6515622,1.6242313,1.8623998,2.1005683,2.338737,2.5769055,2.8111696,2.436347,2.0615244,1.6867018,1.3118792,0.93705654,1.6008049,2.260649,2.9243972,3.5881457,4.251894,3.6857557,3.1235218,2.5612879,1.999054,1.43682,1.9639144,2.4871042,3.0141985,3.5373883,4.0605783,3.2992198,2.5378613,1.7765031,1.0112402,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.62470436,1.2494087,1.8741131,2.4988174,3.1235218,3.1118085,3.1000953,3.0883822,3.076669,3.0610514,3.3265507,3.5881457,3.8497405,4.1113358,4.376835,5.0483923,5.7238536,6.3993154,7.0747766,7.7502384,8.062591,8.374943,8.687295,8.999647,9.311999,9.425227,9.538455,9.651682,9.761005,9.874233,8.511597,7.1489606,5.786324,4.423688,3.0610514,2.87364,2.6862288,2.4988174,2.3114061,2.1239948,2.2879796,2.4480603,2.612045,2.77603,2.9361105,2.9868677,3.0376248,3.0883822,3.1391394,3.1859922,2.5495746,1.9131571,1.2767396,0.63641757,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.5505207,0.6637484,0.77307165,0.8862993,0.999527,1.0893283,1.175225,1.261122,1.3509232,1.43682,1.1869383,0.93705654,0.6871748,0.43729305,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.47633708,0.63641757,0.80040246,0.96438736,1.1244678,1.4485333,1.7765031,2.1005683,2.4246337,2.7486992,2.5886188,2.4246337,2.260649,2.1005683,1.9365835,2.5769055,3.213323,3.8497405,4.4861584,5.12648,5.099149,5.0757227,5.0483923,5.024966,5.001539,5.423215,5.8487945,6.2743745,6.699954,7.125534,8.062591,8.999647,9.936704,10.87376,11.810817,11.139259,10.4637985,9.788337,9.112875,8.437413,9.163632,9.885946,10.612165,11.338385,12.0606985,10.951848,9.839094,8.726339,7.6135845,6.5008297,6.126007,5.7511845,5.376362,5.001539,4.6267166,4.224563,3.8263142,3.4241607,3.0259118,2.6237583,2.514435,2.4012074,2.2879796,2.174752,2.0615244,1.6515622,1.2376955,0.8238289,0.41386664,0.0,0.0,0.0,0.0,0.0,0.0,0.28892577,0.57394713,0.8628729,1.1517987,1.43682,0.5231899,0.5036679,0.48024148,0.45681506,0.43338865,0.41386664,0.39434463,0.37872702,0.359205,0.3435874,0.3240654,0.31625658,0.30454338,0.29673457,0.28502136,0.27330816,0.30844778,0.3435874,0.37872702,0.41386664,0.44900626,0.43338865,0.42167544,0.40605783,0.39044023,0.37482262,0.3631094,0.3513962,0.3357786,0.3240654,0.31235218,0.39044023,0.46852827,0.5466163,0.62079996,0.698888,0.62470436,0.5505207,0.47633708,0.39824903,0.3240654,0.3709182,0.41386664,0.46071947,0.5036679,0.5505207,0.6871748,0.8238289,0.96438736,1.1010414,1.2376955,1.0580931,0.8784905,0.698888,0.5192855,0.3357786,0.3709182,0.40605783,0.44119745,0.47633708,0.5114767,0.58566034,0.6637484,0.737932,0.81211567,0.8862993,0.9058213,0.92143893,0.94096094,0.95657855,0.97610056,0.79259366,0.60908675,0.42557985,0.24597734,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.07027924,0.078088045,0.08589685,0.093705654,0.10151446,0.10151446,0.10541886,0.10932326,0.10932326,0.113227665,1.33921,2.5612879,3.78727,5.0132523,6.239235,5.1616197,4.084005,3.0063896,1.9287747,0.8511597,0.679366,0.5114767,0.339683,0.1717937,0.0,0.078088045,0.15617609,0.23426414,0.30844778,0.38653582,0.30844778,0.23426414,0.15617609,0.078088045,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.18741131,0.22645533,0.26159495,0.30063897,0.3357786,0.39824903,0.45681506,0.5192855,0.57785153,0.63641757,0.679366,0.71841,0.75745404,0.79649806,0.8394465,0.8941081,0.95267415,1.0112402,1.0659018,1.1244678,1.1322767,1.1400855,1.1478943,1.1557031,1.1635119,1.2455044,1.3274968,1.4094892,1.4914817,1.5734742,1.6086137,1.639849,1.6710842,1.7062237,1.737459,1.7725986,1.8077383,1.8428779,1.8780174,1.9131571,2.2137961,2.514435,2.8111696,3.1118085,3.4124475,3.5959544,3.7833657,3.9668727,4.154284,4.337791,4.3612175,4.388548,4.4119744,4.4393053,4.462732,4.2089458,3.959064,3.7052777,3.4514916,3.2016098,3.1586614,3.1196175,3.0805733,3.0415294,2.998581,2.951728,2.9048753,2.8580225,2.8111696,2.7643168,3.7013733,4.6423345,5.5832953,6.524256,7.461313,6.910792,6.356367,5.805846,5.251421,4.7009,4.689187,4.6735697,4.661856,4.650143,4.6384296,6.4969254,8.359325,10.217821,12.076316,13.938716,11.943566,9.952321,7.9610763,5.9659266,3.9746814,5.4154058,6.8561306,8.296855,9.733675,11.174399,12.583888,13.989473,15.398962,16.804546,18.214037,17.323833,16.43363,15.543426,14.653222,13.763018,14.750832,15.74255,16.734268,17.722082,18.7138,17.483913,16.254026,15.024139,13.794253,12.564366,10.77615,8.987934,7.1997175,5.4115014,3.6232853,2.9283018,2.233318,1.5383345,0.8433509,0.14836729,0.12884527,0.10932326,0.08980125,0.07027924,0.05075723,1.5461433,3.0415294,4.5369153,6.028397,7.523783,7.7697606,8.015738,8.261715,8.503788,8.749765,7.918128,7.0903945,6.2587566,5.4310236,4.5993857,4.0332475,3.4632049,2.8970666,2.330928,1.7608855,1.620327,1.475864,1.3353056,1.1908426,1.0502841,1.1713207,1.2884527,1.4094892,1.5305257,1.6515622,1.5539521,1.456342,1.358732,1.261122,1.1635119,1.0698062,0.97610056,0.8862993,0.79259366,0.698888,0.5583295,0.42167544,0.28111696,0.14055848,0.0,0.0,0.0,0.0,0.0,0.0,1.4290112,2.854118,4.283129,5.708236,7.137247,6.4891167,5.8370814,5.1889505,4.5369153,3.8887846,3.2718892,2.6510892,2.0341935,1.4172981,0.80040246,1.1596074,1.5188124,1.8819219,2.241127,2.6003318,2.736986,2.87364,3.0141985,3.1508527,3.2875066,3.1586614,3.0337205,2.9048753,2.77603,2.6510892,2.67842,2.7057507,2.7330816,2.7604125,2.787743,2.97125,3.1586614,3.3421683,3.5256753,3.7130866,3.5256753,3.3421683,3.1586614,2.97125,2.787743,2.5183394,2.25284,1.9834363,1.717937,1.4485333,1.5305257,1.6086137,1.6906061,1.7686942,1.8506867,2.3075018,2.7643168,3.2211318,3.6818514,4.138666,3.9942036,3.8458362,3.7013733,3.5569105,3.4124475,3.3343596,3.2562714,3.1781836,3.1039999,3.0259118,3.2679846,3.5100577,3.7521305,3.9942036,4.2362766,3.8106966,3.3812122,2.9556324,2.5261483,2.1005683,2.1708477,2.2450314,2.3192148,2.3894942,2.463678,2.1591344,1.8584955,1.5539521,1.2533131,0.94876975,1.1517987,1.3548276,1.5578566,1.7608855,1.9639144,1.8584955,1.7530766,1.6476578,1.542239,1.43682,1.2884527,1.1361811,0.9878138,0.8394465,0.6871748,0.95657855,1.2220778,1.4914817,1.756981,2.0263848,1.9834363,1.9404879,1.8975395,1.8545911,1.8116426,1.9639144,2.1161861,2.2684577,2.4207294,2.5769055,2.4051118,2.233318,2.0654287,1.893635,1.7257458,2.1083772,2.494913,2.8814487,3.2640803,3.6506162,3.2836022,2.9165885,2.5456703,2.1786566,1.8116426,2.2684577,2.7213683,3.1781836,3.631094,4.087909,3.4827268,2.8775444,2.2723622,1.6671798,1.0619974,0.8667773,0.6676528,0.46852827,0.27330816,0.07418364,0.5583295,1.0463798,1.5305257,2.0146716,2.4988174,2.4910088,2.4792955,2.4714866,2.4597735,2.4480603,2.795552,3.1391394,3.4866312,3.8302186,4.173806,4.5993857,5.024966,5.4505453,5.8761253,6.3017054,6.5437784,6.7897553,7.0357327,7.28171,7.523783,7.601871,7.676055,7.7502384,7.824422,7.898606,6.8287997,5.755089,4.6813784,3.611572,2.5378613,2.3699722,2.2020829,2.0341935,1.8663043,1.698415,1.8311646,1.9600099,2.0888553,2.2216048,2.35045,2.3894942,2.4285383,2.4714866,2.5105307,2.5495746,2.0380979,1.5305257,1.0190489,0.5114767,0.0,0.45291066,0.9058213,1.358732,1.8116426,2.260649,1.893635,1.5227169,1.1517987,0.78088045,0.41386664,0.3318742,0.24597734,0.1639849,0.08199245,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.10151446,0.1796025,0.25769055,0.3357786,0.41386664,0.5388075,0.6637484,0.78868926,0.9136301,1.038571,0.9956226,0.95267415,0.9097257,0.8667773,0.8238289,0.92924774,1.0346665,1.1400855,1.2455044,1.3509232,1.4329157,1.5149081,1.5969005,1.678893,1.7608855,1.8116426,1.8584955,1.9053483,1.9522011,1.999054,2.0537157,2.1083772,2.1669433,2.2216048,2.2762666,2.194274,2.1161861,2.0341935,1.9561055,1.8741131,2.0537157,2.2294137,2.4090161,2.5847144,2.7643168,2.6042364,2.4480603,2.2918842,2.1318035,1.9756275,2.494913,3.0141985,3.533484,4.056674,4.575959,4.646239,4.7204223,4.7907014,4.8648853,4.939069,5.3256044,5.7121406,6.098676,6.4891167,6.8756523,7.621393,8.36323,9.108971,9.854712,10.600452,10.0265045,9.448653,8.874706,8.300759,7.726812,8.253906,8.784905,9.315904,9.846903,10.373997,9.589212,8.804427,8.019642,7.2348576,6.4500723,6.133816,5.813655,5.4973984,5.181142,4.860981,4.493967,4.126953,3.7599394,3.3929255,3.0259118,2.900971,2.7799344,2.6588979,2.533957,2.4129205,1.9678187,1.5227169,1.077615,0.63251317,0.18741131,0.20302892,0.21864653,0.23426414,0.24597734,0.26159495,0.5075723,0.75354964,0.9956226,1.2415999,1.4875772,0.48805028,0.49195468,0.4958591,0.5036679,0.5075723,0.5114767,0.48805028,0.46852827,0.44510186,0.42167544,0.39824903,0.39434463,0.38653582,0.37872702,0.3709182,0.3631094,0.39434463,0.42557985,0.46071947,0.49195468,0.5231899,0.4958591,0.46462387,0.43338865,0.40605783,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.42948425,0.48414588,0.5388075,0.59346914,0.6481308,0.60127795,0.5505207,0.4997635,0.44900626,0.39824903,0.42557985,0.45681506,0.48414588,0.5114767,0.5388075,0.6871748,0.8394465,0.9878138,1.1361811,1.2884527,1.1010414,0.91753453,0.7340276,0.5466163,0.3631094,0.42167544,0.47633708,0.5349031,0.59346914,0.6481308,0.698888,0.74964523,0.80040246,0.8511597,0.9019169,0.93315214,0.96829176,1.0034313,1.038571,1.0737107,0.8706817,0.6715572,0.46852827,0.26549935,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.06637484,0.06637484,0.07027924,0.07418364,0.07418364,0.078088045,0.08589685,0.08980125,0.093705654,0.10151446,2.4480603,4.7985106,7.1489606,9.499411,11.849861,9.721962,7.590158,5.4583545,3.330455,1.1986516,0.96048295,0.71841,0.48024148,0.23816854,0.0,0.15617609,0.30844778,0.46462387,0.62079996,0.77307165,0.62079996,0.46462387,0.30844778,0.15617609,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.22645533,0.3357786,0.44900626,0.5622339,0.6754616,0.79649806,0.9136301,1.0346665,1.1557031,1.2767396,1.3157835,1.358732,1.4016805,1.4446288,1.4875772,1.3665408,1.2415999,1.1205635,0.9956226,0.8745861,0.9019169,0.92924774,0.95657855,0.98390937,1.0112402,1.116659,1.2181735,1.319688,1.4212024,1.5266213,1.5539521,1.5812829,1.6086137,1.6359446,1.6632754,1.6945106,1.7257458,1.7608855,1.7921207,1.8233559,2.0888553,2.35045,2.612045,2.87364,3.1391394,3.2718892,3.4007344,3.533484,3.6662338,3.7989833,4.0605783,4.3260775,4.5876727,4.8492675,5.1108627,4.7204223,4.3260775,3.9356375,3.541293,3.1508527,3.1313305,3.1157131,3.096191,3.0805733,3.0610514,2.9673457,2.87364,2.77603,2.6823244,2.5886188,3.5686235,4.548629,5.5286336,6.5086384,7.4886436,6.996689,6.5008297,6.008875,5.5169206,5.024966,5.1108627,5.2006636,5.2865605,5.376362,5.462259,7.082586,8.702912,10.323239,11.943566,13.563893,11.650736,9.741484,7.832231,5.9229784,4.0137253,5.704332,7.3988423,9.089449,10.783959,12.4745655,13.200784,13.930907,14.657126,15.383345,16.113468,15.894821,15.676175,15.461433,15.242786,15.024139,16.093946,17.159847,18.22575,19.295555,20.361458,18.627903,16.894348,15.15689,13.423335,11.685876,10.049932,8.413987,6.774138,5.138193,3.4983444,2.8619268,2.2216048,1.5812829,0.94096094,0.30063897,0.26159495,0.21864653,0.1796025,0.14055848,0.10151446,1.678893,3.2562714,4.83365,6.4110284,7.988407,8.0040245,8.015738,8.031356,8.046973,8.062591,7.6409154,7.2192397,6.79366,6.3719845,5.950309,5.12648,4.3065557,3.4827268,2.6588979,1.8389735,1.8897307,1.9443923,1.9951496,2.0459068,2.1005683,2.2762666,2.455869,2.631567,2.8111696,2.9868677,2.854118,2.7213683,2.5886188,2.455869,2.3231194,2.1396124,1.9561055,1.7686942,1.5851873,1.4016805,1.1205635,0.8394465,0.5583295,0.28111696,0.0,0.0,0.0,0.0,0.0,0.0,1.0815194,2.1591344,3.240654,4.318269,5.3997884,5.0132523,4.6267166,4.2362766,3.8497405,3.4632049,2.8892577,2.3192148,1.7452679,1.1713207,0.60127795,0.8706817,1.1400855,1.4094892,1.678893,1.9482968,2.0732377,2.1981785,2.3231194,2.4480603,2.5769055,2.5573835,2.541766,2.522244,2.5066261,2.4871042,2.4910088,2.4988174,2.5027218,2.5066261,2.514435,2.6432803,2.77603,2.9087796,3.0415294,3.174279,3.1313305,3.084478,3.0415294,2.9946766,2.951728,2.7135596,2.4792955,2.2450314,2.0107672,1.7765031,1.796025,1.8194515,1.8428779,1.8663043,1.8858263,2.2137961,2.541766,2.8697357,3.1977055,3.5256753,3.435874,3.3460727,3.2562714,3.1664703,3.076669,3.057147,3.0415294,3.0220075,3.0063896,2.9868677,3.1977055,3.408543,3.619381,3.8263142,4.037152,3.7091823,3.377308,3.049338,2.717464,2.3855898,2.4441557,2.5027218,2.5612879,2.6159496,2.6745155,2.358259,2.0380979,1.7218413,1.4055848,1.0893283,1.2806439,1.4719596,1.6632754,1.8584955,2.0498111,1.9287747,1.8038338,1.6827974,1.5617609,1.43682,1.2767396,1.1127546,0.94876975,0.78868926,0.62470436,0.96048295,1.2962615,1.6281357,1.9639144,2.2996929,2.241127,2.1786566,2.1200905,2.0615244,1.999054,2.069333,2.135708,2.2020829,2.2684577,2.338737,2.3738766,2.4090161,2.4441557,2.4792955,2.514435,2.619854,2.7291772,2.8345962,2.9439192,3.049338,2.8775444,2.7057507,2.533957,2.358259,2.1864653,2.5730011,2.9556324,3.3421683,3.7287042,4.1113358,3.6662338,3.2172275,2.7682211,2.3231194,1.8741131,1.5305257,1.1869383,0.8394465,0.4958591,0.14836729,0.4958591,0.8394465,1.1869383,1.5305257,1.8741131,1.8663043,1.8584955,1.8506867,1.8467822,1.8389735,2.2645533,2.6940374,3.1196175,3.5491016,3.9746814,4.1503797,4.3260775,4.5017757,4.6735697,4.8492675,5.02887,5.2045684,5.3841705,5.559869,5.735567,5.774611,5.813655,5.8487945,5.8878384,5.9268827,5.142098,4.3612175,3.5764325,2.795552,2.0107672,1.8663043,1.717937,1.5695697,1.4212024,1.2767396,1.3743496,1.4680552,1.5656652,1.6632754,1.7608855,1.7921207,1.8233559,1.8506867,1.8819219,1.9131571,1.5305257,1.1478943,0.76526284,0.38263142,0.0,0.9058213,1.8116426,2.7135596,3.619381,4.5252023,3.7833657,3.0454338,2.3035975,1.5656652,0.8238289,0.659844,0.4958591,0.3318742,0.1639849,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.20693332,0.359205,0.5153811,0.6715572,0.8238289,0.9878138,1.1517987,1.3118792,1.475864,1.6359446,1.4407244,1.2415999,1.0463798,0.8472553,0.6481308,0.77307165,0.8941081,1.0190489,1.1400855,1.261122,1.678893,2.0927596,2.5066261,2.9243972,3.338264,3.4710135,3.6037633,3.736513,3.8692627,3.998108,4.0488653,4.095718,4.142571,4.1894236,4.2362766,3.9161155,3.59205,3.2718892,2.9478238,2.6237583,2.6549935,2.6862288,2.7135596,2.7447948,2.77603,2.6237583,2.4714866,2.3192148,2.1669433,2.0107672,2.416825,2.8189783,3.2211318,3.6232853,4.025439,4.193328,4.365122,4.5369153,4.704805,4.8765984,5.22409,5.575486,5.9268827,6.2743745,6.6257706,7.1762915,7.7307167,8.281238,8.835662,9.386183,8.913751,8.437413,7.9610763,7.4886436,7.012306,7.348085,7.6838636,8.015738,8.351517,8.687295,8.23048,7.773665,7.3168497,6.8561306,6.3993154,6.141625,5.8800297,5.618435,5.3607445,5.099149,4.7633705,4.4314966,4.095718,3.7599394,3.4241607,3.2914112,3.1586614,3.0259118,2.893162,2.7643168,2.2840753,1.8077383,1.3314011,0.8511597,0.37482262,0.40605783,0.43338865,0.46462387,0.4958591,0.5231899,0.7262188,0.92924774,1.1322767,1.3353056,1.5383345,0.44900626,0.48414588,0.5153811,0.5466163,0.58175594,0.61299115,0.58566034,0.5583295,0.5309987,0.5036679,0.47633708,0.46852827,0.46462387,0.46071947,0.45681506,0.44900626,0.48024148,0.5114767,0.5388075,0.5700427,0.60127795,0.5544251,0.5114767,0.46462387,0.42167544,0.37482262,0.38653582,0.39824903,0.41386664,0.42557985,0.43729305,0.46852827,0.5036679,0.5349031,0.5661383,0.60127795,0.57394713,0.5505207,0.5231899,0.4997635,0.47633708,0.48414588,0.4958591,0.5036679,0.5153811,0.5231899,0.6871748,0.8511597,1.0112402,1.175225,1.33921,1.1478943,0.95657855,0.76916724,0.57785153,0.38653582,0.46852827,0.5466163,0.62860876,0.7066968,0.78868926,0.81211567,0.8394465,0.8628729,0.8862993,0.9136301,0.96438736,1.0190489,1.0698062,1.1205635,1.175225,0.95267415,0.7301232,0.5075723,0.28502136,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.058566034,0.058566034,0.05466163,0.05075723,0.05075723,0.058566034,0.06637484,0.07418364,0.078088045,0.08589685,3.5608149,7.0357327,10.510651,13.985569,17.464392,14.278399,11.096312,7.914223,4.732136,1.5500476,1.2415999,0.92924774,0.62079996,0.30844778,0.0,0.23426414,0.46462387,0.698888,0.92924774,1.1635119,0.92924774,0.698888,0.46462387,0.23426414,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.26159495,0.44900626,0.63641757,0.8238289,1.0112402,1.1908426,1.3743496,1.5539521,1.7335546,1.9131571,1.9561055,2.0029583,2.0459068,2.0927596,2.135708,1.8350691,1.53443,1.2298868,0.92924774,0.62470436,0.6715572,0.71841,0.76916724,0.8160201,0.8628729,0.98390937,1.1088502,1.2298868,1.3509232,1.475864,1.4992905,1.5188124,1.542239,1.5656652,1.5890918,1.6164225,1.6476578,1.678893,1.7062237,1.737459,1.9639144,2.1864653,2.4129205,2.639376,2.8619268,2.9439192,3.0220075,3.1039999,3.182088,3.2640803,3.7638438,4.263607,4.7633705,5.263134,5.7628975,5.2318993,4.6969957,4.165997,3.631094,3.1000953,3.1039999,3.1118085,3.1157131,3.1196175,3.1235218,2.9829633,2.8385005,2.697942,2.5534792,2.4129205,3.4319696,4.4510183,5.473972,6.493021,7.5120697,7.0786815,6.649197,6.2158084,5.7824197,5.349031,5.5364423,5.7238536,5.911265,6.098676,6.2860875,7.6682463,9.0465,10.4286585,11.806912,13.189071,11.361811,9.530646,7.703386,5.8761253,4.0488653,5.9932575,7.941554,9.885946,11.8303385,13.774731,13.821584,13.868437,13.919194,13.966047,14.012899,14.465811,14.922626,15.37944,15.832351,16.289165,17.433157,18.577147,19.721136,20.86903,22.01302,19.771893,17.530766,15.293544,13.052417,10.81129,9.323712,7.8361354,6.348558,4.860981,3.3734035,2.7916477,2.2059872,1.620327,1.0346665,0.44900626,0.39044023,0.3318742,0.26940376,0.21083772,0.14836729,1.8116426,3.4710135,5.1303844,6.7897553,8.449126,8.234385,8.019642,7.8049,7.590158,7.375416,7.3597984,7.3441806,7.328563,7.3168497,7.3012323,6.223617,5.1460023,4.068387,2.9907722,1.9131571,2.1591344,2.4090161,2.6549935,2.900971,3.1508527,3.3851168,3.619381,3.853645,4.0918136,4.3260775,4.1581883,3.9902992,3.8224099,3.6545205,3.4866312,3.2094188,2.9322062,2.6549935,2.377781,2.1005683,1.678893,1.261122,0.8394465,0.42167544,0.0,0.0,0.0,0.0,0.0,0.0,0.7340276,1.4641509,2.1981785,2.9283018,3.6623292,3.5373883,3.4124475,3.2875066,3.1625657,3.0376248,2.5105307,1.9834363,1.456342,0.92924774,0.39824903,0.58175594,0.76135844,0.94096094,1.1205635,1.3001659,1.4133936,1.5266213,1.6359446,1.7491722,1.8623998,1.9561055,2.0459068,2.1396124,2.233318,2.3231194,2.3075018,2.2918842,2.2723622,2.2567444,2.2372224,2.3192148,2.397303,2.4792955,2.5573835,2.639376,2.7330816,2.8267872,2.9243972,3.018103,3.1118085,2.9087796,2.7057507,2.5066261,2.3035975,2.1005683,2.0654287,2.0302892,1.9951496,1.9600099,1.9248703,2.1239948,2.3192148,2.5183394,2.7135596,2.912684,2.8775444,2.8424048,2.8072653,2.7721257,2.736986,2.7799344,2.822883,2.8658314,2.9087796,2.951728,3.1274261,3.3031244,3.4827268,3.6584249,3.8380275,3.6037633,3.3734035,3.1391394,2.9087796,2.6745155,2.717464,2.7604125,2.803361,2.8463092,2.8892577,2.5534792,2.2216048,1.8897307,1.5578566,1.2259823,1.4055848,1.5890918,1.7725986,1.9561055,2.135708,1.999054,1.8584955,1.717937,1.5773785,1.43682,1.261122,1.0893283,0.9136301,0.737932,0.5622339,0.96438736,1.3665408,1.7686942,2.1708477,2.5769055,2.4988174,2.4207294,2.3426414,2.2645533,2.1864653,2.1708477,2.1513257,2.135708,2.1161861,2.1005683,2.338737,2.5808098,2.8189783,3.0610514,3.2992198,3.1313305,2.959537,2.7916477,2.619854,2.4480603,2.4714866,2.494913,2.5183394,2.541766,2.5612879,2.8775444,3.193801,3.506153,3.8224099,4.138666,3.8458362,3.5569105,3.2679846,2.979059,2.6862288,2.194274,1.7023194,1.2103647,0.71841,0.22645533,0.42948425,0.63641757,0.8394465,1.0463798,1.2494087,1.2455044,1.2415999,1.2337911,1.2298868,1.2259823,1.7335546,2.2450314,2.7565079,3.2640803,3.775557,3.7013733,3.6232853,3.5491016,3.474918,3.4007344,3.5100577,3.619381,3.7287042,3.8419318,3.951255,3.951255,3.951255,3.951255,3.951255,3.951255,3.4593005,2.9634414,2.4714866,1.979532,1.4875772,1.358732,1.2337911,1.1049459,0.97610056,0.8511597,0.9136301,0.98000497,1.0463798,1.1088502,1.175225,1.1947471,1.2142692,1.2337911,1.2533131,1.2767396,1.0190489,0.76526284,0.5114767,0.25378615,0.0,1.358732,2.7135596,4.0722914,5.4310236,6.785851,5.677001,4.5681505,3.4593005,2.3465457,1.2376955,0.9917182,0.7418364,0.4958591,0.24597734,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.30844778,0.5388075,0.77307165,1.0034313,1.2376955,1.43682,1.6359446,1.8389735,2.0380979,2.2372224,1.8858263,1.53443,1.1791295,0.8277333,0.47633708,0.61689556,0.75354964,0.8941081,1.0346665,1.175225,1.9209659,2.6706111,3.416352,4.165997,4.911738,5.1303844,5.349031,5.563773,5.7824197,6.001066,6.04011,6.0791545,6.1181984,6.1611466,6.2001905,5.6340523,5.0718184,4.50568,3.9395418,3.3734035,3.2562714,3.1391394,3.0220075,2.9048753,2.787743,2.639376,2.4910088,2.3465457,2.1981785,2.0498111,2.3348327,2.619854,2.9048753,3.1898966,3.474918,3.7443218,4.009821,4.279225,4.5447245,4.814128,5.12648,5.4388323,5.7511845,6.0635366,6.375889,6.735094,7.094299,7.453504,7.816613,8.175818,7.800996,7.426173,7.0513506,6.676528,6.3017054,6.4383593,6.578918,6.719476,6.860035,7.000593,6.871748,6.7389984,6.610153,6.481308,6.348558,6.1494336,5.9464045,5.743376,5.5403466,5.337318,5.036679,4.732136,4.4314966,4.126953,3.8263142,3.6818514,3.541293,3.39683,3.2562714,3.1118085,2.6042364,2.0927596,1.5812829,1.0737107,0.5622339,0.60908675,0.6520352,0.698888,0.7418364,0.78868926,0.94876975,1.1088502,1.2689307,1.4290112,1.5890918,0.41386664,0.47243267,0.5309987,0.59346914,0.6520352,0.7106012,0.679366,0.6481308,0.61689556,0.58175594,0.5505207,0.5466163,0.5466163,0.5427119,0.5388075,0.5388075,0.5661383,0.59346914,0.62079996,0.6481308,0.6754616,0.61689556,0.5544251,0.4958591,0.43338865,0.37482262,0.39824903,0.42557985,0.44900626,0.47633708,0.4997635,0.5114767,0.5192855,0.5309987,0.5388075,0.5505207,0.5505207,0.5505207,0.5505207,0.5505207,0.5505207,0.5427119,0.5349031,0.5270943,0.5192855,0.5114767,0.6871748,0.8628729,1.038571,1.2142692,1.3860629,1.1908426,0.9956226,0.80430686,0.60908675,0.41386664,0.5153811,0.61689556,0.71841,0.8238289,0.92534333,0.92534333,0.92534333,0.92534333,0.92534333,0.92534333,0.9956226,1.0659018,1.1361811,1.2064602,1.2767396,1.0307622,0.78868926,0.5466163,0.30454338,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05466163,0.046852827,0.039044023,0.031235218,0.023426414,0.03513962,0.046852827,0.05466163,0.06637484,0.07418364,4.6735697,9.272955,13.8762455,18.475632,23.075018,18.838741,14.606369,10.370092,6.133816,1.901444,1.5188124,1.1400855,0.76135844,0.37872702,0.0,0.30844778,0.62079996,0.92924774,1.2415999,1.5500476,1.2415999,0.92924774,0.62079996,0.30844778,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.30063897,0.5622339,0.8238289,1.0893283,1.3509232,1.5890918,1.8311646,2.069333,2.3114061,2.5495746,2.5964274,2.6432803,2.6940374,2.7408905,2.787743,2.3035975,1.8233559,1.33921,0.8589685,0.37482262,0.44119745,0.5114767,0.57785153,0.6442264,0.7106012,0.8550641,0.9956226,1.1400855,1.2806439,1.4251068,1.4407244,1.4602464,1.475864,1.4953861,1.5110037,1.5383345,1.5656652,1.5969005,1.6242313,1.6515622,1.8389735,2.0263848,2.2137961,2.4012074,2.5886188,2.6159496,2.6432803,2.6706111,2.697942,2.7252727,3.4632049,4.2011366,4.939069,5.6730967,6.4110284,5.7394714,5.067914,4.396357,3.7208953,3.049338,3.076669,3.1039999,3.1313305,3.1586614,3.1859922,2.998581,2.8072653,2.6159496,2.4285383,2.2372224,3.2992198,4.357313,5.4193106,6.477403,7.5394006,7.164578,6.79366,6.4188375,6.0479193,5.6730967,5.9620223,6.250948,6.5359693,6.824895,7.113821,8.253906,9.393991,10.534078,11.674163,12.814248,11.06898,9.323712,7.578445,5.833177,4.087909,6.2860875,8.484266,10.67854,12.8767185,15.074897,14.442384,13.809871,13.177358,12.544845,11.912332,13.040704,14.169076,15.293544,16.421915,17.550287,18.772366,19.994444,21.216522,22.4386,23.660677,20.915882,18.171087,15.426293,12.681499,9.936704,8.601398,7.262188,5.9268827,4.5876727,3.2484627,2.7213683,2.1903696,1.6593709,1.1283722,0.60127795,0.5192855,0.44119745,0.359205,0.28111696,0.19912452,1.9443923,3.6857557,5.4271193,7.168483,8.913751,8.468649,8.023546,7.578445,7.1333427,6.688241,7.0786815,7.473026,7.8634663,8.257811,8.648251,7.3168497,5.985449,4.6540475,3.3187418,1.9873407,2.4285383,2.87364,3.3148375,3.7560349,4.2011366,4.493967,4.786797,5.0757227,5.368553,5.661383,5.4583545,5.2592297,5.056201,4.853172,4.650143,4.279225,3.9083066,3.541293,3.1703746,2.7994564,2.241127,1.678893,1.1205635,0.5583295,0.0,0.0,0.0,0.0,0.0,0.0,0.38653582,0.76916724,1.1557031,1.5383345,1.9248703,2.0615244,2.1981785,2.338737,2.475391,2.612045,2.1318035,1.6476578,1.1635119,0.6832704,0.19912452,0.28892577,0.37872702,0.46852827,0.5583295,0.6481308,0.74964523,0.8511597,0.94876975,1.0502841,1.1517987,1.3509232,1.5539521,1.756981,1.9600099,2.1630387,2.1239948,2.0810463,2.0420024,2.0029583,1.9639144,1.9912452,2.018576,2.0459068,2.0732377,2.1005683,2.3348327,2.5690966,2.803361,3.0415294,3.2757936,3.1039999,2.9361105,2.7643168,2.5964274,2.4246337,2.330928,2.241127,2.1474214,2.0537157,1.9639144,2.0302892,2.096664,2.1669433,2.233318,2.2996929,2.3192148,2.338737,2.358259,2.3816853,2.4012074,2.5027218,2.6042364,2.7057507,2.8111696,2.912684,3.057147,3.2016098,3.3460727,3.49444,3.638903,3.5022488,3.3655949,3.232845,3.096191,2.9634414,2.9907722,3.018103,3.0454338,3.0727646,3.1000953,2.7526035,2.4051118,2.05762,1.7101282,1.3626363,1.53443,1.7062237,1.8819219,2.0537157,2.2255092,2.069333,1.9092526,1.7530766,1.5969005,1.43682,1.2494087,1.0619974,0.8745861,0.6871748,0.4997635,0.96829176,1.4407244,1.9092526,2.3816853,2.8502135,2.7565079,2.6588979,2.5651922,2.4714866,2.3738766,2.2723622,2.1708477,2.069333,1.9639144,1.8623998,2.3075018,2.7526035,3.1977055,3.6428072,4.087909,3.638903,3.193801,2.7447948,2.2957885,1.8506867,2.069333,2.2840753,2.5027218,2.7213683,2.9361105,3.182088,3.4280653,3.6740425,3.9161155,4.1620927,4.029343,3.8965936,3.7638438,3.631094,3.4983444,2.8580225,2.2216048,1.5812829,0.94096094,0.30063897,0.3631094,0.42948425,0.4958591,0.5583295,0.62470436,0.62079996,0.62079996,0.61689556,0.61689556,0.61299115,1.2064602,1.796025,2.3894942,2.9829633,3.5764325,3.2484627,2.9243972,2.6003318,2.2762666,1.9482968,1.9912452,2.0341935,2.077142,2.1200905,2.1630387,2.1239948,2.0888553,2.0498111,2.0107672,1.9756275,1.7725986,1.5695697,1.3665408,1.1635119,0.96438736,0.8550641,0.74574083,0.64032197,0.5309987,0.42557985,0.45681506,0.48805028,0.5231899,0.5544251,0.58566034,0.59737355,0.60908675,0.61689556,0.62860876,0.63641757,0.5114767,0.38263142,0.25378615,0.12884527,0.0,1.8116426,3.619381,5.4310236,7.238762,9.050405,7.570636,6.0908675,4.6110992,3.1313305,1.6515622,1.319688,0.9917182,0.659844,0.3318742,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.40996224,0.71841,1.0307622,1.33921,1.6515622,1.8858263,2.1239948,2.3621633,2.6003318,2.8385005,2.330928,1.8233559,1.3157835,0.80821127,0.30063897,0.45681506,0.61689556,0.77307165,0.92924774,1.0893283,2.1669433,3.2484627,4.3260775,5.407597,6.4891167,6.7897553,7.094299,7.394938,7.6955767,8.00012,8.031356,8.066495,8.097731,8.128965,8.164105,7.355894,6.547683,5.7394714,4.93126,4.123049,3.8614538,3.5959544,3.330455,3.0649557,2.7994564,2.6588979,2.514435,2.3738766,2.2294137,2.0888553,2.2567444,2.4207294,2.5886188,2.7565079,2.9243972,3.2914112,3.6545205,4.0215344,4.3846436,4.7516575,5.024966,5.298274,5.575486,5.8487945,6.126007,6.2938967,6.461786,6.6257706,6.79366,6.9615493,6.688241,6.4110284,6.13772,5.8644123,5.5871997,5.532538,5.477876,5.423215,5.368553,5.3138914,5.5091114,5.708236,5.903456,6.1025805,6.3017054,6.153338,6.008875,5.8644123,5.7199492,5.575486,5.3060827,5.036679,4.7633705,4.493967,4.224563,4.0722914,3.9200199,3.767748,3.6154766,3.4632049,2.920493,2.377781,1.8350691,1.2923572,0.74964523,0.80821127,0.8706817,0.92924774,0.9917182,1.0502841,1.1674163,1.2845483,1.4016805,1.5188124,1.6359446,0.37482262,0.46071947,0.5505207,0.63641757,0.7262188,0.81211567,0.77307165,0.737932,0.698888,0.6637484,0.62470436,0.62470436,0.62470436,0.62470436,0.62470436,0.62470436,0.6481308,0.6754616,0.698888,0.7262188,0.74964523,0.6754616,0.60127795,0.5231899,0.44900626,0.37482262,0.41386664,0.44900626,0.48805028,0.5231899,0.5622339,0.5505207,0.5388075,0.5231899,0.5114767,0.4997635,0.5231899,0.5505207,0.57394713,0.60127795,0.62470436,0.60127795,0.57394713,0.5505207,0.5231899,0.4997635,0.6871748,0.8745861,1.0619974,1.2494087,1.43682,1.2376955,1.038571,0.8355421,0.63641757,0.43729305,0.5622339,0.6871748,0.81211567,0.93705654,1.0619974,1.038571,1.0112402,0.9878138,0.96438736,0.93705654,1.0268579,1.1127546,1.1986516,1.2884527,1.3743496,1.1127546,0.8511597,0.58566034,0.3240654,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,5.786324,11.514082,17.237936,22.96179,28.685644,23.399082,18.112522,12.825961,7.535496,2.2489357,1.7999294,1.3509232,0.9019169,0.44900626,0.0,0.38653582,0.77307165,1.1635119,1.5500476,1.9365835,1.5500476,1.1635119,0.77307165,0.38653582,0.0,0.0,0.0,0.0,0.0,0.0,0.3357786,0.6754616,1.0112402,1.3509232,1.6867018,1.9873407,2.2879796,2.5886188,2.8892577,3.1859922,3.2367494,3.2875066,3.338264,3.3890212,3.435874,2.77603,2.1122816,1.4485333,0.78868926,0.12494087,0.21083772,0.30063897,0.38653582,0.47633708,0.5622339,0.7262188,0.8862993,1.0502841,1.2142692,1.3743496,1.3860629,1.4016805,1.4133936,1.4251068,1.43682,1.4641509,1.4875772,1.5110037,1.5383345,1.5617609,1.7140326,1.8623998,2.0107672,2.1630387,2.3114061,2.2879796,2.260649,2.2372224,2.2137961,2.1864653,3.1625657,4.138666,5.1108627,6.086963,7.0630636,6.250948,5.4388323,4.6267166,3.8106966,2.998581,3.049338,3.1000953,3.1508527,3.2016098,3.2484627,3.0141985,2.77603,2.5378613,2.2996929,2.0615244,3.1625657,4.263607,5.3607445,6.461786,7.562827,7.250475,6.9381227,6.6257706,6.3134184,6.001066,6.387602,6.774138,7.1606736,7.551114,7.9376497,8.835662,9.737579,10.6355915,11.537509,12.439425,10.77615,9.112875,7.4495993,5.786324,4.123049,6.575013,9.023073,11.475039,13.923099,16.375063,15.063184,13.751305,12.435521,11.123642,9.811763,11.611692,13.411622,15.211552,17.01148,18.81141,20.111576,21.411741,22.711908,24.012074,25.31224,22.063778,18.81141,15.562947,12.31058,9.062118,7.8751793,6.688241,5.5013027,4.3143644,3.1235218,2.6510892,2.174752,1.698415,1.2259823,0.74964523,0.6481308,0.5505207,0.44900626,0.3513962,0.24988174,2.0732377,3.900498,5.7238536,7.551114,9.37447,8.699008,8.023546,7.348085,6.676528,6.001066,6.801469,7.601871,8.398369,9.198771,9.999174,8.413987,6.824895,5.2358036,3.6506162,2.0615244,2.7018464,3.338264,3.9746814,4.6110992,5.251421,5.5989127,5.950309,6.3017054,6.649197,7.000593,6.7624245,6.524256,6.2860875,6.0518236,5.813655,5.349031,4.8883114,4.423688,3.9629683,3.4983444,2.7994564,2.1005683,1.4016805,0.698888,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.58566034,0.9878138,1.3860629,1.7882162,2.1864653,1.7491722,1.3118792,0.8745861,0.43729305,0.0,0.0,0.0,0.0,0.0,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.74964523,1.0619974,1.3743496,1.6867018,1.999054,1.9365835,1.8741131,1.8116426,1.7491722,1.6867018,1.6632754,1.6359446,1.6125181,1.5890918,1.5617609,1.9365835,2.3114061,2.6862288,3.0610514,3.435874,3.2992198,3.1625657,3.0259118,2.8892577,2.7486992,2.6003318,2.4480603,2.2996929,2.1513257,1.999054,1.9365835,1.8741131,1.8116426,1.7491722,1.6867018,1.7608855,1.8389735,1.9131571,1.9873407,2.0615244,2.2255092,2.3855898,2.5495746,2.7135596,2.87364,2.9868677,3.1000953,3.213323,3.3265507,3.435874,3.4007344,3.3616903,3.3265507,3.2875066,3.2484627,3.2640803,3.2757936,3.2875066,3.2992198,3.310933,2.951728,2.5886188,2.2255092,1.8623998,1.4992905,1.6632754,1.8233559,1.9873407,2.1513257,2.3114061,2.135708,1.9639144,1.7882162,1.6125181,1.43682,1.2376955,1.038571,0.8355421,0.63641757,0.43729305,0.97610056,1.5110037,2.0498111,2.5886188,3.1235218,3.0141985,2.900971,2.787743,2.6745155,2.5612879,2.3738766,2.1864653,1.999054,1.8116426,1.6242313,2.2762666,2.9243972,3.5764325,4.224563,4.8765984,4.1503797,3.4241607,2.7018464,1.9756275,1.2494087,1.6632754,2.0732377,2.4871042,2.900971,3.310933,3.4866312,3.6623292,3.8380275,4.0137253,4.1894236,4.21285,4.2362766,4.263607,4.2870336,4.3143644,3.5256753,2.736986,1.9482968,1.1635119,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.6754616,1.3509232,2.0263848,2.7018464,3.3734035,2.7994564,2.2255092,1.6515622,1.0737107,0.4997635,0.47633708,0.44900626,0.42557985,0.39824903,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.3513962,0.26159495,0.1756981,0.08589685,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.2645533,4.5252023,6.785851,9.050405,11.311053,9.464272,7.6135845,5.7628975,3.912211,2.0615244,1.6515622,1.2376955,0.8238289,0.41386664,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.5114767,0.9019169,1.2884527,1.6749885,2.0615244,2.338737,2.612045,2.8892577,3.1625657,3.435874,2.77603,2.1122816,1.4485333,0.78868926,0.12494087,0.30063897,0.47633708,0.6481308,0.8238289,0.999527,2.4129205,3.8263142,5.2358036,6.649197,8.062591,8.449126,8.835662,9.226103,9.612638,9.999174,10.0265045,10.049932,10.073358,10.100689,10.124115,9.073831,8.023546,6.9732623,5.9268827,4.8765984,4.462732,4.0488653,3.638903,3.2250361,2.8111696,2.6745155,2.5378613,2.4012074,2.260649,2.1239948,2.174752,2.2255092,2.2762666,2.3231194,2.3738766,2.8385005,3.2992198,3.7638438,4.224563,4.689187,4.9234514,5.1616197,5.3997884,5.6379566,5.8761253,5.8487945,5.825368,5.801942,5.774611,5.7511845,5.575486,5.3997884,5.22409,5.0483923,4.8765984,4.6267166,4.376835,4.123049,3.873167,3.6232853,4.1503797,4.6735697,5.2006636,5.7238536,6.250948,6.1611466,6.0752497,5.989353,5.899552,5.813655,5.575486,5.337318,5.099149,4.860981,4.6267166,4.462732,4.298747,4.138666,3.9746814,3.8106966,3.2367494,2.6628022,2.0888553,1.5110037,0.93705654,1.0112402,1.0893283,1.1635119,1.2376955,1.3118792,1.3860629,1.4641509,1.5383345,1.6125181,1.6867018,0.3513962,0.42167544,0.48805028,0.5583295,0.62860876,0.698888,0.6715572,0.64032197,0.60908675,0.58175594,0.5505207,0.5544251,0.5583295,0.5661383,0.5700427,0.57394713,0.59737355,0.62079996,0.6442264,0.6637484,0.6871748,0.62079996,0.5544251,0.48414588,0.41777104,0.3513962,0.38653582,0.42167544,0.45681506,0.48805028,0.5231899,0.5153811,0.5036679,0.4958591,0.48414588,0.47633708,0.5192855,0.5583295,0.60127795,0.6442264,0.6871748,0.6676528,0.6481308,0.62860876,0.60908675,0.58566034,0.7223144,0.8589685,0.9917182,1.1283722,1.261122,1.097137,0.93315214,0.76916724,0.60127795,0.43729305,0.5583295,0.679366,0.79649806,0.91753453,1.038571,0.9956226,0.95657855,0.91753453,0.8784905,0.8394465,0.8902037,0.94096094,0.9956226,1.0463798,1.1010414,0.8941081,0.6910792,0.48414588,0.28111696,0.07418364,0.07027924,0.06637484,0.058566034,0.05466163,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,5.7824197,11.2642,16.745981,22.231667,27.713448,22.657246,17.601046,12.548749,7.492548,2.436347,2.5261483,2.612045,2.7018464,2.787743,2.87364,2.8385005,2.7994564,2.7643168,2.7252727,2.6862288,2.1981785,1.7062237,1.2181735,0.7262188,0.23816854,0.21474212,0.19131571,0.1717937,0.14836729,0.12494087,0.48805028,0.8511597,1.2142692,1.5734742,1.9365835,2.2840753,2.6276627,2.97125,3.3187418,3.6623292,3.6935644,3.7208953,3.7521305,3.7833657,3.8106966,3.213323,2.6159496,2.018576,1.4212024,0.8238289,0.81211567,0.80040246,0.78868926,0.77307165,0.76135844,0.8472553,0.93315214,1.0190489,1.1010414,1.1869383,1.2220778,1.2572175,1.2923572,1.3274968,1.3626363,1.4016805,1.4407244,1.4836729,1.5227169,1.5617609,1.7140326,1.8623998,2.0107672,2.1630387,2.3114061,2.2762666,2.2372224,2.1981785,2.1630387,2.1239948,3.2484627,4.369026,5.493494,6.6140575,7.7385254,6.7702336,5.801942,4.83365,3.8692627,2.900971,2.920493,2.9400148,2.959537,2.979059,2.998581,2.912684,2.8267872,2.736986,2.6510892,2.5612879,3.6232853,4.6813784,5.743376,6.801469,7.8634663,7.558923,7.2582836,6.9537406,6.6531014,6.348558,6.6335793,6.914696,7.195813,7.480835,7.7619514,8.617016,9.47208,10.327144,11.182208,12.037272,10.58093,9.120684,7.6643414,6.2079997,4.7516575,6.8756523,9.0035515,11.131451,13.25935,15.387249,14.2901125,13.192975,12.095839,10.998701,9.901564,11.291532,12.685403,14.079274,15.469242,16.863113,17.565907,18.268698,18.97149,19.674282,20.37317,17.866545,15.359919,12.853292,10.346666,7.8361354,6.832704,5.8292727,4.8219366,3.8185053,2.8111696,2.4792955,2.1474214,1.815547,1.4836729,1.1517987,0.98000497,0.80821127,0.64032197,0.46852827,0.30063897,1.8545911,3.408543,4.9663997,6.520352,8.074304,8.905942,9.733675,10.565312,11.39695,12.224684,11.810817,11.400854,10.986988,10.573121,10.163159,8.804427,7.4417906,6.083059,4.7243266,3.3616903,3.716991,4.0722914,4.4275923,4.7828927,5.138193,5.493494,5.8487945,6.2040954,6.559396,6.910792,6.89127,6.871748,6.852226,6.832704,6.813182,6.6921453,6.571109,6.453977,6.3329406,6.211904,5.0132523,3.8185053,2.619854,1.4212024,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.62470436,1.1010414,1.5734742,2.0498111,2.5261483,2.0888553,1.6515622,1.2142692,0.77307165,0.3357786,0.3474918,0.359205,0.3670138,0.37872702,0.38653582,0.39434463,0.40215343,0.40996224,0.41777104,0.42557985,0.75354964,1.0854238,1.4133936,1.7452679,2.0732377,2.0341935,1.9951496,1.9561055,1.9131571,1.8741131,1.8584955,1.8389735,1.8233559,1.8038338,1.7882162,2.1630387,2.5378613,2.912684,3.2875066,3.6623292,3.5256753,3.3929255,3.2562714,3.1235218,2.9868677,2.7994564,2.612045,2.4246337,2.2372224,2.0498111,1.9873407,1.9248703,1.8623998,1.7999294,1.737459,1.8389735,1.9365835,2.0380979,2.135708,2.2372224,2.3933985,2.5534792,2.7096553,2.8658314,3.0259118,3.049338,3.06886,3.0922866,3.1157131,3.1391394,3.0805733,3.0220075,2.9634414,2.9087796,2.8502135,2.8658314,2.8853533,2.900971,2.920493,2.9361105,2.67842,2.416825,2.1591344,1.8975395,1.6359446,1.7491722,1.8584955,1.9678187,2.077142,2.1864653,2.0302892,1.8741131,1.7140326,1.5578566,1.4016805,1.1908426,0.98000497,0.76916724,0.5583295,0.3513962,0.8667773,1.3860629,1.901444,2.4207294,2.9361105,2.8463092,2.7526035,2.6588979,2.5690966,2.475391,2.3855898,2.2996929,2.2137961,2.1239948,2.0380979,2.533957,3.0337205,3.5295796,4.029343,4.5252023,3.8380275,3.1508527,2.463678,1.7765031,1.0893283,1.475864,1.8663043,2.2567444,2.6471848,3.0376248,3.260176,3.4827268,3.7052777,3.9278288,4.1503797,4.0605783,3.970777,3.8809757,3.7911747,3.7013733,3.0610514,2.4246337,1.7882162,1.1517987,0.5114767,0.40996224,0.30844778,0.20693332,0.10151446,0.0,0.0,0.0,0.0,0.0,0.0,0.5388075,1.0815194,1.620327,2.1591344,2.7018464,2.241127,1.7804074,1.319688,0.8589685,0.39824903,0.37872702,0.359205,0.339683,0.32016098,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.07027924,0.14055848,0.21083772,0.28111696,0.3513962,0.28111696,0.21083772,0.14055848,0.07027924,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.10932326,0.08199245,0.05466163,0.027330816,0.0,0.0,0.0,0.0,0.0,0.0,1.8116426,3.619381,5.4310236,7.238762,9.050405,7.5979667,6.1494336,4.7009,3.2484627,1.7999294,1.4407244,1.0815194,0.71841,0.359205,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10541886,0.15617609,0.21083772,0.26159495,0.26549935,0.26940376,0.26940376,0.27330816,0.27330816,0.22645533,0.1756981,0.12494087,0.07418364,0.023426414,0.13665408,0.24597734,0.3553006,0.46462387,0.57394713,0.9058213,1.2415999,1.5734742,1.9053483,2.2372224,2.416825,2.592523,2.7682211,2.9478238,3.1235218,2.631567,2.1396124,1.6476578,1.1557031,0.6637484,0.94486535,1.2259823,1.5110037,1.7921207,2.0732377,3.1469483,4.2167544,5.2865605,6.356367,7.426173,7.800996,8.175818,8.550641,8.925464,9.300286,9.807858,10.315431,10.823003,11.330575,11.838148,10.799577,9.761005,8.726339,7.687768,6.649197,6.2353306,5.8214636,5.4036927,4.989826,4.575959,4.165997,3.7599394,3.3538816,2.9439192,2.5378613,2.631567,2.7291772,2.822883,2.9165885,3.0141985,3.2992198,3.5881457,3.873167,4.1620927,4.4510183,4.806319,5.1616197,5.5169206,5.8683167,6.223617,6.1064854,5.989353,5.872221,5.755089,5.6379566,5.395884,5.153811,4.911738,4.6657605,4.423688,4.181615,3.9395418,3.697469,3.455396,3.213323,3.6428072,4.0722914,4.5017757,4.93126,5.3607445,5.4036927,5.4427366,5.481781,5.520825,5.563773,5.3021784,5.040583,4.7828927,4.521298,4.263607,4.142571,4.0215344,3.9044023,3.7833657,3.6623292,3.1664703,2.6706111,2.1786566,1.6827974,1.1869383,1.2298868,1.2728351,1.3157835,1.358732,1.4016805,1.43682,1.475864,1.5110037,1.5500476,1.5890918,0.3240654,0.37872702,0.42948425,0.48414588,0.5349031,0.58566034,0.5661383,0.5427119,0.5192855,0.4958591,0.47633708,0.48414588,0.4958591,0.5036679,0.5153811,0.5231899,0.5466163,0.5661383,0.58566034,0.60518235,0.62470436,0.5661383,0.5036679,0.44510186,0.38653582,0.3240654,0.359205,0.39044023,0.42167544,0.45681506,0.48805028,0.48024148,0.47243267,0.46462387,0.45681506,0.44900626,0.5114767,0.5700427,0.62860876,0.6910792,0.74964523,0.7340276,0.71841,0.7066968,0.6910792,0.6754616,0.75745404,0.8394465,0.92143893,1.0034313,1.0893283,0.95657855,0.8277333,0.698888,0.5661383,0.43729305,0.5544251,0.6676528,0.78088045,0.8980125,1.0112402,0.95657855,0.9019169,0.8472553,0.79259366,0.737932,0.75354964,0.77307165,0.78868926,0.80821127,0.8238289,0.679366,0.5309987,0.38263142,0.23426414,0.08589685,0.078088045,0.06637484,0.058566034,0.046852827,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.10932326,0.21474212,0.3240654,0.42948425,0.5388075,5.7785153,11.018223,16.25793,21.497639,26.737347,21.91541,17.093473,12.271536,7.445695,2.6237583,3.2484627,3.873167,4.5017757,5.12648,5.7511845,5.2865605,4.825841,4.3612175,3.900498,3.435874,2.8463092,2.25284,1.6593709,1.0659018,0.47633708,0.42948425,0.38653582,0.339683,0.29673457,0.24988174,0.63641757,1.0268579,1.4133936,1.7999294,2.1864653,2.5769055,2.9673457,3.357786,3.7482262,4.138666,4.1464753,4.1581883,4.165997,4.1777105,4.1894236,3.6545205,3.1235218,2.5886188,2.05762,1.5266213,1.4133936,1.3001659,1.1869383,1.0737107,0.96438736,0.96829176,0.97610056,0.98390937,0.9917182,0.999527,1.0580931,1.116659,1.1713207,1.2298868,1.2884527,1.3431144,1.397776,1.4524376,1.5070993,1.5617609,1.7140326,1.8623998,2.0107672,2.1630387,2.3114061,2.260649,2.2137961,2.1630387,2.1122816,2.0615244,3.3343596,4.60329,5.872221,7.141152,8.413987,7.289519,6.168956,5.044488,3.9239242,2.7994564,2.7916477,2.7799344,2.7682211,2.7604125,2.7486992,2.8111696,2.87364,2.9361105,2.998581,3.0610514,4.084005,5.1030536,6.1221027,7.141152,8.164105,7.871275,7.578445,7.2856145,6.9927845,6.699954,6.8756523,7.055255,7.230953,7.4105554,7.5862536,8.398369,9.20658,10.018696,10.826907,11.639023,10.38571,9.132397,7.8790836,6.6257706,5.376362,7.180196,8.98403,10.791768,12.595602,14.399435,13.51704,12.634645,11.752251,10.869856,9.987461,10.971371,11.959184,12.943093,13.927003,14.9109125,15.016331,15.12175,15.227169,15.332587,15.438006,13.673217,11.908427,10.143637,8.378847,6.6140575,5.7902284,4.9663997,4.1464753,3.3226464,2.4988174,2.3114061,2.1200905,1.9287747,1.7413634,1.5500476,1.3118792,1.0698062,0.8316377,0.58956474,0.3513962,1.6359446,2.920493,4.2050414,5.4895897,6.774138,9.108971,11.443803,13.778636,16.113468,18.448301,16.82407,15.199838,13.575606,11.951375,10.323239,9.190963,8.058686,6.9264097,5.794133,4.661856,4.73604,4.806319,4.8805027,4.950782,5.024966,5.3841705,5.743376,6.1064854,6.46569,6.824895,7.0240197,7.2192397,7.4183645,7.6135845,7.812709,8.03526,8.257811,8.480362,8.702912,8.925464,7.230953,5.5364423,3.8380275,2.1435168,0.44900626,0.359205,0.26940376,0.1796025,0.08980125,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.6637484,1.2142692,1.7608855,2.3114061,2.8619268,2.4246337,1.9873407,1.5500476,1.1127546,0.6754616,0.6949836,0.7145056,0.7340276,0.75354964,0.77307165,0.7027924,0.62860876,0.5583295,0.48414588,0.41386664,0.76135844,1.1088502,1.456342,1.8038338,2.1513257,2.1318035,2.1161861,2.096664,2.0810463,2.0615244,2.0537157,2.0420024,2.0341935,2.0224805,2.0107672,2.3855898,2.7643168,3.1391394,3.513962,3.8887846,3.7560349,3.6232853,3.4905357,3.357786,3.2250361,2.998581,2.77603,2.5495746,2.3231194,2.1005683,2.0380979,1.9756275,1.9131571,1.8506867,1.7882162,1.9131571,2.0380979,2.1630387,2.2879796,2.4129205,2.5651922,2.717464,2.8697357,3.0220075,3.174279,3.1079042,3.0415294,2.97125,2.9048753,2.8385005,2.7604125,2.6823244,2.6042364,2.5261483,2.4480603,2.4714866,2.494913,2.5183394,2.541766,2.5612879,2.4051118,2.2489357,2.0888553,1.9326792,1.7765031,1.8311646,1.8897307,1.9482968,2.0068626,2.0615244,1.9209659,1.7843118,1.6437533,1.5031948,1.3626363,1.1439898,0.92143893,0.7027924,0.48414588,0.26159495,0.76135844,1.2572175,1.7530766,2.25284,2.7486992,2.67842,2.6042364,2.533957,2.4597735,2.3855898,2.4012074,2.4129205,2.4246337,2.436347,2.4480603,2.795552,3.1391394,3.4866312,3.8302186,4.173806,3.5256753,2.87364,2.2255092,1.5734742,0.92534333,1.2923572,1.6593709,2.0263848,2.3933985,2.7643168,3.0337205,3.3031244,3.5725281,3.8419318,4.1113358,3.9083066,3.7013733,3.4983444,3.2914112,3.0883822,2.6003318,2.1122816,1.6242313,1.1361811,0.6481308,0.5192855,0.39044023,0.26159495,0.12884527,0.0,0.0,0.0,0.0,0.0,0.0,0.40605783,0.80821127,1.2142692,1.620327,2.0263848,1.678893,1.3353056,0.9917182,0.6442264,0.30063897,0.28502136,0.26940376,0.25378615,0.23816854,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.05075723,0.10541886,0.15617609,0.21083772,0.26159495,0.21083772,0.15617609,0.10541886,0.05075723,0.0,0.05466163,0.10932326,0.1639849,0.21864653,0.27330816,0.21864653,0.1639849,0.10932326,0.05466163,0.0,0.0,0.0,0.0,0.0,0.0,1.358732,2.7135596,4.0722914,5.4310236,6.785851,5.735567,4.689187,3.638903,2.5886188,1.5383345,1.2298868,0.92143893,0.61689556,0.30844778,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10541886,0.21083772,0.31625658,0.42167544,0.5231899,0.5309987,0.5349031,0.5388075,0.5466163,0.5505207,0.44900626,0.3513962,0.24988174,0.14836729,0.05075723,0.24597734,0.44119745,0.63641757,0.8316377,1.0268579,1.3040704,1.5812829,1.8584955,2.135708,2.4129205,2.4910088,2.5730011,2.6510892,2.7330816,2.8111696,2.4910088,2.1669433,1.8467822,1.5227169,1.1986516,1.5890918,1.979532,2.3699722,2.7604125,3.1508527,3.8770714,4.60329,5.3334136,6.0596323,6.785851,7.1489606,7.5120697,7.8751793,8.238289,8.601398,9.589212,10.58093,11.568744,12.560462,13.548276,12.525322,11.498465,10.475512,9.448653,8.4257,8.007929,7.590158,7.172387,6.754616,6.336845,5.661383,4.9820175,4.3065557,3.6271896,2.951728,3.0883822,3.2289407,3.3694992,3.5100577,3.6506162,3.7638438,3.873167,3.9863946,4.0996222,4.21285,4.6852827,5.1577153,5.630148,6.1025805,6.575013,6.364176,6.153338,5.9464045,5.735567,5.5247293,5.2162814,4.903929,4.5954814,4.283129,3.9746814,3.7404175,3.506153,3.2718892,3.0337205,2.7994564,3.135235,3.4710135,3.8067923,4.138666,4.474445,4.6423345,4.8102236,4.9781127,5.1460023,5.3138914,5.02887,4.747753,4.466636,4.181615,3.900498,3.8224099,3.7443218,3.6662338,3.5881457,3.513962,3.096191,2.6823244,2.2684577,1.8506867,1.43682,1.4485333,1.456342,1.4680552,1.475864,1.4875772,1.4875772,1.4875772,1.4875772,1.4875772,1.4875772,0.30063897,0.3357786,0.3709182,0.40605783,0.44119745,0.47633708,0.46071947,0.44510186,0.42948425,0.41386664,0.39824903,0.41386664,0.42948425,0.44510186,0.46071947,0.47633708,0.49195468,0.5114767,0.5270943,0.5466163,0.5622339,0.5114767,0.45681506,0.40605783,0.3513962,0.30063897,0.3318742,0.359205,0.39044023,0.42167544,0.44900626,0.44510186,0.44119745,0.43338865,0.42948425,0.42557985,0.5036679,0.58175594,0.6559396,0.7340276,0.81211567,0.80430686,0.79259366,0.78088045,0.77307165,0.76135844,0.79259366,0.8238289,0.8511597,0.8823949,0.9136301,0.8160201,0.7223144,0.62860876,0.5309987,0.43729305,0.5466163,0.6559396,0.76916724,0.8784905,0.9878138,0.91753453,0.8472553,0.77697605,0.7066968,0.63641757,0.62079996,0.60127795,0.58566034,0.5661383,0.5505207,0.46071947,0.3709182,0.28111696,0.19131571,0.10151446,0.08589685,0.07027924,0.05466163,0.039044023,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.15617609,0.30844778,0.46462387,0.62079996,0.77307165,5.7707067,10.768341,15.765976,20.76361,25.761246,21.173573,16.581997,11.990419,7.4027467,2.8111696,3.9746814,5.138193,6.3017054,7.461313,8.624825,7.7385254,6.8483214,5.9620223,5.0757227,4.1894236,3.49444,2.7994564,2.1005683,1.4055848,0.7106012,0.6442264,0.57785153,0.5114767,0.44119745,0.37482262,0.78868926,1.1986516,1.6125181,2.0263848,2.436347,2.87364,3.3070288,3.7443218,4.1777105,4.6110992,4.60329,4.591577,4.5837684,4.572055,4.564246,4.095718,3.6271896,3.1586614,2.6940374,2.2255092,2.0107672,1.7999294,1.5890918,1.3743496,1.1635119,1.0932326,1.0229534,0.95267415,0.8823949,0.81211567,0.8941081,0.97219616,1.0541886,1.1322767,1.2142692,1.2806439,1.3509232,1.4212024,1.4914817,1.5617609,1.7140326,1.8623998,2.0107672,2.1630387,2.3114061,2.2489357,2.1864653,2.1239948,2.0615244,1.999054,3.416352,4.83365,6.250948,7.6682463,9.085544,7.8088045,6.532065,5.2553253,3.978586,2.7018464,2.6588979,2.619854,2.5808098,2.541766,2.4988174,2.7135596,2.9243972,3.1391394,3.349977,3.5608149,4.5408196,5.520825,6.5008297,7.480835,8.460839,8.179723,7.898606,7.6135845,7.3324676,7.0513506,7.1216297,7.195813,7.266093,7.3402762,7.4105554,8.175818,8.941081,9.706344,10.471607,11.23687,10.19049,9.14411,8.093826,7.0474463,6.001066,7.480835,8.964508,10.44818,11.931853,13.411622,12.743969,12.076316,11.408664,10.741011,10.073358,10.651209,11.229061,11.806912,12.384764,12.962616,12.470661,11.978706,11.486752,10.990892,10.498938,9.475985,8.456935,7.433982,6.4110284,5.388075,4.747753,4.1074314,3.4671092,2.8267872,2.1864653,2.1396124,2.0927596,2.0459068,1.999054,1.9482968,1.639849,1.3314011,1.0190489,0.7106012,0.39824903,1.4133936,2.4285383,3.4436827,4.4588275,5.473972,9.315904,13.153932,16.995863,20.83389,24.675823,21.837322,18.998821,16.164225,13.325725,10.487225,9.581403,8.675582,7.773665,6.8678436,5.9620223,5.7511845,5.5442514,5.3334136,5.1225758,4.911738,5.278752,5.6418614,6.008875,6.3719845,6.7389984,7.152865,7.5667315,7.9805984,8.398369,8.812236,9.378374,9.940608,10.506746,11.072885,11.639023,9.444749,7.2543793,5.0601053,2.8658314,0.6754616,0.5388075,0.40605783,0.26940376,0.13665408,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.698888,1.3235924,1.9482968,2.5769055,3.2016098,2.7643168,2.3231194,1.8858263,1.4485333,1.0112402,1.0424755,1.0737107,1.1010414,1.1322767,1.1635119,1.0112402,0.8589685,0.7066968,0.5544251,0.39824903,0.76526284,1.1283722,1.4953861,1.8584955,2.2255092,2.2294137,2.233318,2.241127,2.2450314,2.2489357,2.2489357,2.2450314,2.241127,2.241127,2.2372224,2.612045,2.9868677,3.3616903,3.736513,4.1113358,3.9824903,3.853645,3.7208953,3.59205,3.4632049,3.2016098,2.9361105,2.6745155,2.4129205,2.1513257,2.0888553,2.0263848,1.9639144,1.901444,1.8389735,1.9873407,2.135708,2.2879796,2.436347,2.5886188,2.7330816,2.8814487,3.0298162,3.1781836,3.3265507,3.1664703,3.0102942,2.854118,2.6940374,2.5378613,2.4402514,2.3426414,2.2450314,2.1474214,2.0498111,2.077142,2.1044729,2.1318035,2.1591344,2.1864653,2.1318035,2.077142,2.0224805,1.9678187,1.9131571,1.9170616,1.9209659,1.9287747,1.9326792,1.9365835,1.815547,1.6906061,1.5695697,1.4485333,1.3235924,1.0932326,0.8667773,0.63641757,0.40605783,0.1756981,0.6520352,1.1283722,1.6086137,2.084951,2.5612879,2.5105307,2.455869,2.4051118,2.3543546,2.2996929,2.4129205,2.5261483,2.639376,2.7486992,2.8619268,3.0532427,3.2484627,3.4397783,3.631094,3.8263142,3.213323,2.6003318,1.9873407,1.3743496,0.76135844,1.1088502,1.4524376,1.796025,2.1435168,2.4871042,2.803361,3.1235218,3.4397783,3.7560349,4.0761957,3.7560349,3.435874,3.1157131,2.795552,2.475391,2.135708,1.7999294,1.4641509,1.1244678,0.78868926,0.62860876,0.47243267,0.31625658,0.15617609,0.0,0.0,0.0,0.0,0.0,0.0,0.26940376,0.5388075,0.80821127,1.0815194,1.3509232,1.1205635,0.8902037,0.659844,0.42948425,0.19912452,0.19131571,0.1796025,0.1717937,0.16008049,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.08199245,0.1639849,0.24597734,0.3318742,0.41386664,0.3318742,0.24597734,0.1639849,0.08199245,0.0,0.0,0.0,0.0,0.0,0.0,0.9058213,1.8116426,2.7135596,3.619381,4.5252023,3.873167,3.2250361,2.5769055,1.9248703,1.2767396,1.0190489,0.76526284,0.5114767,0.25378615,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15617609,0.31625658,0.47243267,0.62860876,0.78868926,0.79649806,0.80430686,0.80821127,0.8160201,0.8238289,0.6754616,0.5231899,0.37482262,0.22645533,0.07418364,0.3553006,0.63641757,0.9136301,1.1947471,1.475864,1.698415,1.9209659,2.1435168,2.366068,2.5886188,2.5690966,2.5534792,2.533957,2.5183394,2.4988174,2.3465457,2.194274,2.0420024,1.8897307,1.737459,2.233318,2.7330816,3.2289407,3.7287042,4.224563,4.6110992,4.9937305,5.380266,5.7668023,6.1494336,6.5008297,6.8483214,7.1997175,7.551114,7.898606,9.37447,10.84643,12.318389,13.790349,15.262308,14.251068,13.235924,12.224684,11.213444,10.198298,9.780528,9.358852,8.941081,8.519405,8.101635,7.152865,6.2040954,5.2592297,4.31046,3.3616903,3.5491016,3.7326086,3.9161155,4.1035266,4.2870336,4.224563,4.1620927,4.0996222,4.037152,3.9746814,4.564246,5.153811,5.743376,6.336845,6.9264097,6.621866,6.321227,6.016684,5.716045,5.4115014,5.036679,4.657952,4.279225,3.9044023,3.5256753,3.2992198,3.06886,2.8424048,2.6159496,2.3855898,2.6276627,2.8658314,3.1079042,3.3460727,3.5881457,3.8809757,4.1777105,4.474445,4.7672753,5.0640097,4.755562,4.4510183,4.1464753,3.8419318,3.5373883,3.5022488,3.4671092,3.4319696,3.39683,3.3616903,3.0259118,2.6940374,2.358259,2.0224805,1.6867018,1.6632754,1.6437533,1.620327,1.5969005,1.5734742,1.5383345,1.4992905,1.4641509,1.4251068,1.3860629,0.27330816,0.29283017,0.30844778,0.3279698,0.3435874,0.3631094,0.3553006,0.3474918,0.339683,0.3318742,0.3240654,0.3435874,0.3631094,0.38653582,0.40605783,0.42557985,0.44119745,0.45681506,0.46852827,0.48414588,0.4997635,0.45681506,0.40996224,0.3631094,0.32016098,0.27330816,0.30063897,0.3318742,0.359205,0.38653582,0.41386664,0.40996224,0.40605783,0.40605783,0.40215343,0.39824903,0.4958591,0.58956474,0.6832704,0.78088045,0.8745861,0.8706817,0.8667773,0.8589685,0.8550641,0.8511597,0.8277333,0.80430686,0.78088045,0.76135844,0.737932,0.679366,0.61689556,0.5583295,0.4958591,0.43729305,0.5427119,0.6481308,0.75354964,0.8589685,0.96438736,0.8784905,0.79259366,0.7066968,0.62079996,0.5388075,0.48414588,0.43338865,0.37872702,0.3279698,0.27330816,0.24207294,0.21083772,0.1756981,0.14446288,0.113227665,0.093705654,0.07418364,0.05075723,0.031235218,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.20302892,0.40605783,0.60908675,0.80821127,1.0112402,5.7668023,10.522364,15.277926,20.033487,24.78905,20.431738,16.074425,11.713207,7.355894,2.998581,4.7009,6.3993154,8.101635,9.80005,11.498465,10.186585,8.874706,7.562827,6.250948,4.939069,4.138666,3.3421683,2.5456703,1.7491722,0.94876975,0.8589685,0.76916724,0.679366,0.58956474,0.4997635,0.93705654,1.3743496,1.8116426,2.2489357,2.6862288,3.1664703,3.6467118,4.126953,4.607195,5.087436,5.056201,5.02887,4.997635,4.9663997,4.939069,4.5369153,4.1308575,3.7287042,3.3265507,2.9243972,2.612045,2.2996929,1.9873407,1.6749885,1.3626363,1.2142692,1.0659018,0.92143893,0.77307165,0.62470436,0.7262188,0.8316377,0.93315214,1.0346665,1.1361811,1.2220778,1.3079748,1.3938715,1.475864,1.5617609,1.7140326,1.8623998,2.0107672,2.1630387,2.3114061,2.2372224,2.1630387,2.0888553,2.0107672,1.9365835,3.5022488,5.067914,6.6335793,8.1992445,9.761005,8.32809,6.899079,5.466163,4.0332475,2.6003318,2.5300527,2.4597735,2.3894942,2.3192148,2.2489357,2.612045,2.9751544,3.338264,3.7013733,4.0605783,5.001539,5.9425,6.883461,7.824422,8.761478,8.488171,8.218767,7.9454584,7.6721506,7.3988423,7.367607,7.336372,7.3012323,7.269997,7.238762,7.957172,8.675582,9.397896,10.116306,10.838621,9.99527,9.151918,8.308568,7.4691215,6.6257706,7.785378,8.944985,10.104593,11.2642,12.423808,11.970898,11.521891,11.06898,10.61607,10.163159,10.331048,10.502842,10.670732,10.8425255,11.014318,9.921086,8.831758,7.7424297,6.6531014,5.563773,5.282656,5.001539,4.7243266,4.4432096,4.1620927,3.7052777,3.2484627,2.7916477,2.330928,1.8741131,1.9717231,2.0654287,2.1591344,2.2567444,2.35045,1.9717231,1.5890918,1.2103647,0.8316377,0.44900626,1.1947471,1.9404879,2.6862288,3.4280653,4.173806,9.518932,14.864059,20.209187,25.554314,30.899439,26.850574,22.801708,18.74894,14.700074,10.651209,9.971844,9.296382,8.617016,7.941554,7.262188,6.7702336,6.278279,5.786324,5.2943697,4.7985106,5.169429,5.5403466,5.911265,6.278279,6.649197,7.28171,7.914223,8.546737,9.17925,9.811763,10.721489,11.62731,12.533132,13.442857,14.348679,11.6585455,8.968412,6.278279,3.5881457,0.9019169,0.71841,0.5388075,0.359205,0.1796025,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.737932,1.43682,2.135708,2.8385005,3.5373883,3.1000953,2.6628022,2.2255092,1.7882162,1.3509232,1.3899672,1.4290112,1.4680552,1.5110037,1.5500476,1.3157835,1.0854238,0.8511597,0.62079996,0.38653582,0.76916724,1.1517987,1.53443,1.9170616,2.2996929,2.3270237,2.3543546,2.3816853,2.4090161,2.436347,2.4441557,2.4480603,2.4519646,2.455869,2.463678,2.8385005,3.213323,3.5881457,3.9629683,4.337791,4.2089458,4.084005,3.9551594,3.8263142,3.7013733,3.4007344,3.1000953,2.7994564,2.4988174,2.1981785,2.135708,2.0732377,2.0107672,1.9482968,1.8858263,2.0615244,2.2372224,2.4129205,2.5886188,2.7643168,2.9048753,3.049338,3.1898966,3.3343596,3.474918,3.2289407,2.979059,2.7330816,2.4831998,2.2372224,2.1200905,2.0029583,1.8858263,1.7686942,1.6515622,1.6827974,1.7140326,1.7491722,1.7804074,1.8116426,1.8584955,1.9092526,1.9561055,2.0029583,2.0498111,2.0029583,1.9561055,1.9092526,1.8584955,1.8116426,1.7062237,1.6008049,1.4992905,1.3938715,1.2884527,1.0463798,0.80821127,0.5661383,0.3279698,0.08589685,0.5466163,1.0034313,1.4602464,1.9170616,2.3738766,2.3426414,2.3114061,2.2762666,2.2450314,2.2137961,2.4246337,2.639376,2.8502135,3.0610514,3.2757936,3.3148375,3.3538816,3.39683,3.435874,3.474918,2.900971,2.3231194,1.7491722,1.175225,0.60127795,0.92143893,1.2455044,1.5656652,1.8897307,2.2137961,2.5769055,2.9439192,3.3070288,3.6740425,4.037152,3.6037633,3.1664703,2.7330816,2.2957885,1.8623998,1.6749885,1.4875772,1.3001659,1.1127546,0.92534333,0.7418364,0.5544251,0.3709182,0.1835069,0.0,0.0,0.0,0.0,0.0,0.0,0.13665408,0.26940376,0.40605783,0.5388075,0.6754616,0.5583295,0.44510186,0.3318742,0.21474212,0.10151446,0.093705654,0.08980125,0.08589685,0.078088045,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.10932326,0.21864653,0.3318742,0.44119745,0.5505207,0.44119745,0.3318742,0.21864653,0.10932326,0.0,0.0,0.0,0.0,0.0,0.0,0.45291066,0.9058213,1.358732,1.8116426,2.260649,2.0107672,1.7608855,1.5110037,1.261122,1.0112402,0.80821127,0.60908675,0.40605783,0.20302892,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21083772,0.42167544,0.62860876,0.8394465,1.0502841,1.0580931,1.0698062,1.0815194,1.0893283,1.1010414,0.9019169,0.698888,0.4997635,0.30063897,0.10151446,0.46462387,0.8316377,1.1947471,1.5617609,1.9248703,2.0927596,2.260649,2.4285383,2.5964274,2.7643168,2.6471848,2.533957,2.416825,2.3035975,2.1864653,2.2059872,2.2216048,2.241127,2.2567444,2.2762666,2.8814487,3.4866312,4.0918136,4.6930914,5.298274,5.3412223,5.3841705,5.4271193,5.4700675,5.5130157,5.8487945,6.1884775,6.524256,6.8639393,7.1997175,9.155824,11.108025,13.06413,15.020235,16.976341,15.976814,14.973383,13.973856,12.974329,11.974802,11.553126,11.131451,10.705871,10.284196,9.86252,8.644346,7.426173,6.211904,4.9937305,3.775557,4.0059166,4.2362766,4.466636,4.6930914,4.9234514,4.689187,4.4510183,4.21285,3.9746814,3.736513,4.4432096,5.153811,5.860508,6.5672045,7.2739015,6.8795567,6.4852123,6.0908675,5.6965227,5.298274,4.853172,4.40807,3.9668727,3.521771,3.076669,2.854118,2.6354716,2.416825,2.194274,1.9756275,2.1200905,2.2645533,2.4090161,2.5534792,2.7018464,3.1235218,3.5451972,3.9668727,4.388548,4.814128,4.4861584,4.1581883,3.8302186,3.5022488,3.174279,3.182088,3.1898966,3.1977055,3.2055142,3.213323,2.9556324,2.7018464,2.4480603,2.194274,1.9365835,1.8819219,1.8272603,1.7725986,1.717937,1.6632754,1.5890918,1.5110037,1.43682,1.3626363,1.2884527,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.27330816,0.30063897,0.3240654,0.3513962,0.37482262,0.38653582,0.39824903,0.41386664,0.42557985,0.43729305,0.39824903,0.3631094,0.3240654,0.28892577,0.24988174,0.27330816,0.30063897,0.3240654,0.3513962,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.48805028,0.60127795,0.7106012,0.8238289,0.93705654,0.93705654,0.93705654,0.93705654,0.93705654,0.93705654,0.8628729,0.78868926,0.7106012,0.63641757,0.5622339,0.5388075,0.5114767,0.48805028,0.46071947,0.43729305,0.5388075,0.63641757,0.737932,0.8394465,0.93705654,0.8394465,0.737932,0.63641757,0.5388075,0.43729305,0.3513962,0.26159495,0.1756981,0.08589685,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24988174,0.4997635,0.74964523,0.999527,1.2494087,5.7628975,10.276386,14.785972,19.29946,23.81295,19.685997,15.562947,11.435994,7.3129454,3.1859922,5.423215,7.6643414,9.901564,12.138786,14.376009,12.63855,10.901091,9.163632,7.426173,5.688714,4.786797,3.8887846,2.9868677,2.0888553,1.1869383,1.0737107,0.96438736,0.8511597,0.737932,0.62470436,1.0893283,1.5500476,2.0107672,2.475391,2.9361105,3.4632049,3.9863946,4.513489,5.036679,5.563773,5.5130157,5.462259,5.4115014,5.3607445,5.3138914,4.9742084,4.6384296,4.298747,3.9629683,3.6232853,3.213323,2.7994564,2.3855898,1.9756275,1.5617609,1.33921,1.1127546,0.8862993,0.6637484,0.43729305,0.5622339,0.6871748,0.81211567,0.93705654,1.0619974,1.1635119,1.261122,1.3626363,1.4641509,1.5617609,1.7140326,1.8623998,2.0107672,2.1630387,2.3114061,2.2255092,2.135708,2.0498111,1.9639144,1.8741131,3.5881457,5.298274,7.012306,8.726339,10.436467,8.85128,7.262188,5.6730967,4.087909,2.4988174,2.4012074,2.2996929,2.1981785,2.1005683,1.999054,2.514435,3.0259118,3.5373883,4.0488653,4.564246,5.462259,6.364176,7.262188,8.164105,9.062118,8.800523,8.538928,8.273428,8.011833,7.7502384,7.6135845,7.47693,7.336372,7.1997175,7.0630636,7.7385254,8.413987,9.089449,9.761005,10.436467,9.80005,9.163632,8.52331,7.8868923,7.250475,8.086017,8.925464,9.761005,10.600452,11.435994,11.20173,10.963562,10.725393,10.487225,10.249056,10.010887,9.776623,9.538455,9.300286,9.062118,7.375416,5.688714,3.998108,2.3114061,0.62470436,1.0893283,1.5500476,2.0107672,2.475391,2.9361105,2.6628022,2.3855898,2.1122816,1.8389735,1.5617609,1.7999294,2.0380979,2.2762666,2.514435,2.7486992,2.2996929,1.8506867,1.4016805,0.94876975,0.4997635,0.97610056,1.4485333,1.9248703,2.4012074,2.87364,9.725866,16.574188,23.426414,30.274734,37.12306,31.863827,26.600693,21.337559,16.074425,10.81129,10.362284,9.913278,9.464272,9.01136,8.562354,7.7892823,7.012306,6.239235,5.462259,4.689187,5.0640097,5.4388323,5.813655,6.1884775,6.5633,7.4105554,8.261715,9.112875,9.964035,10.81129,12.0606985,13.314012,14.56342,15.812829,17.062239,13.8762455,10.686349,7.5003567,4.3143644,1.1244678,0.9019169,0.6754616,0.44900626,0.22645533,0.0,0.0,0.0,0.0,0.0,0.0,0.77307165,1.5500476,2.3231194,3.1000953,3.873167,3.435874,2.998581,2.5612879,2.1239948,1.6867018,1.737459,1.7882162,1.8389735,1.8858263,1.9365835,1.6242313,1.3118792,0.999527,0.6871748,0.37482262,0.77697605,1.175225,1.5734742,1.9756275,2.3738766,2.4246337,2.475391,2.5261483,2.5769055,2.6237583,2.639376,2.6510892,2.6628022,2.6745155,2.6862288,3.0610514,3.435874,3.8106966,4.1894236,4.564246,4.4393053,4.3143644,4.1894236,4.0605783,3.9356375,3.5998588,3.2640803,2.9243972,2.5886188,2.2489357,2.1864653,2.1239948,2.0615244,1.999054,1.9365835,2.135708,2.338737,2.5378613,2.736986,2.9361105,3.076669,3.213323,3.349977,3.4866312,3.6232853,3.2875066,2.951728,2.612045,2.2762666,1.9365835,1.7999294,1.6632754,1.5266213,1.3860629,1.2494087,1.2884527,1.3235924,1.3626363,1.4016805,1.43682,1.5890918,1.737459,1.8858263,2.0380979,2.1864653,2.0888553,1.9873407,1.8858263,1.7882162,1.6867018,1.6008049,1.5110037,1.4251068,1.33921,1.2494087,0.999527,0.74964523,0.4997635,0.24988174,0.0,0.43729305,0.8745861,1.3118792,1.7491722,2.1864653,2.174752,2.1630387,2.1513257,2.135708,2.1239948,2.436347,2.7486992,3.0610514,3.3734035,3.6857557,3.5764325,3.4632049,3.349977,3.2367494,3.1235218,2.5886188,2.0498111,1.5110037,0.97610056,0.43729305,0.737932,1.038571,1.33921,1.6359446,1.9365835,2.35045,2.7643168,3.174279,3.5881457,3.998108,3.4514916,2.900971,2.35045,1.7999294,1.2494087,1.2142692,1.175225,1.1361811,1.1010414,1.0619974,0.8511597,0.63641757,0.42557985,0.21083772,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13665408,0.27330816,0.41386664,0.5505207,0.6871748,0.5505207,0.41386664,0.27330816,0.13665408,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14836729,0.30063897,0.44900626,0.60127795,0.74964523,0.60127795,0.44900626,0.30063897,0.14836729,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26159495,0.5231899,0.78868926,1.0502841,1.3118792,1.3235924,1.33921,1.3509232,1.3626363,1.3743496,1.1244678,0.8745861,0.62470436,0.37482262,0.12494087,0.57394713,1.0268579,1.475864,1.9248703,2.3738766,2.4871042,2.6003318,2.7135596,2.8267872,2.9361105,2.7252727,2.514435,2.2996929,2.0888553,1.8741131,2.0615244,2.2489357,2.436347,2.6237583,2.8111696,3.5256753,4.2362766,4.950782,5.661383,6.375889,6.0752497,5.774611,5.473972,5.173333,4.8765984,5.2006636,5.5247293,5.8487945,6.1767645,6.5008297,8.937177,11.373524,13.813775,16.250122,18.68647,17.698656,16.710842,15.723028,14.739119,13.751305,13.325725,12.900145,12.4745655,12.0489855,11.623405,10.135828,8.648251,7.1606736,5.677001,4.1894236,4.462732,4.73604,5.0132523,5.2865605,5.563773,5.1499066,4.73604,4.3260775,3.912211,3.4983444,4.3260775,5.1499066,5.9737353,6.801469,7.6252975,7.137247,6.649197,6.1611466,5.6730967,5.1889505,4.6735697,4.1620927,3.6506162,3.1391394,2.6237583,2.4129205,2.1981785,1.9873407,1.7765031,1.5617609,1.6125181,1.6632754,1.7140326,1.7608855,1.8116426,2.3621633,2.912684,3.4632049,4.0137253,4.564246,4.21285,3.8614538,3.513962,3.1625657,2.8111696,2.8619268,2.912684,2.9634414,3.0141985,3.0610514,2.8892577,2.7135596,2.5378613,2.3621633,2.1864653,2.1005683,2.0107672,1.9248703,1.8389735,1.7491722,1.6359446,1.5266213,1.4133936,1.3001659,1.1869383,0.30063897,0.29673457,0.29673457,0.29283017,0.28892577,0.28892577,0.28111696,0.27721256,0.27330816,0.26940376,0.26159495,0.28111696,0.30063897,0.3240654,0.3435874,0.3631094,0.37482262,0.38653582,0.39824903,0.41386664,0.42557985,0.39434463,0.359205,0.3279698,0.29673457,0.26159495,0.28502136,0.30844778,0.3318742,0.3513962,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.46852827,0.5661383,0.659844,0.75354964,0.8511597,0.8433509,0.8355421,0.8277333,0.8199245,0.81211567,0.78478485,0.75745404,0.7301232,0.7027924,0.6754616,0.6871748,0.698888,0.7106012,0.7262188,0.737932,0.80430686,0.8706817,0.94096094,1.0073358,1.0737107,0.96438736,0.8511597,0.737932,0.62470436,0.5114767,0.45681506,0.40215343,0.3474918,0.29283017,0.23816854,0.21083772,0.1835069,0.15617609,0.12884527,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.41386664,0.8238289,1.2376955,1.6515622,2.0615244,5.6809053,9.296382,12.915763,16.531239,20.15062,16.675701,13.204688,9.733675,6.2587566,2.787743,4.5291066,6.2743745,8.015738,9.757101,11.498465,10.131924,8.765383,7.3988423,6.028397,4.661856,3.9200199,3.1781836,2.436347,1.6906061,0.94876975,0.93315214,0.92143893,0.9058213,0.8902037,0.8745861,1.2845483,1.6945106,2.1044729,2.514435,2.9243972,3.3655949,3.8106966,4.251894,4.6930914,5.138193,5.1303844,5.1225758,5.114767,5.1069584,5.099149,4.845363,4.591577,4.3338866,4.0801005,3.8263142,3.541293,3.260176,2.979059,2.6940374,2.4129205,2.2098918,2.0068626,1.8038338,1.6008049,1.4016805,1.3548276,1.3118792,1.2650263,1.2181735,1.175225,1.2572175,1.33921,1.4212024,1.5031948,1.5890918,1.7413634,1.8975395,2.0537157,2.2059872,2.3621633,2.3231194,2.2879796,2.2489357,2.2137961,2.174752,3.7247996,5.2748475,6.824895,8.374943,9.924991,8.453031,6.9810715,5.5091114,4.0332475,2.5612879,2.5456703,2.5261483,2.5105307,2.4910088,2.475391,3.0883822,3.7052777,4.318269,4.9351645,5.548156,6.1299114,6.7116675,7.289519,7.871275,8.449126,8.191436,7.929841,7.6682463,7.4105554,7.1489606,7.113821,7.0786815,7.043542,7.008402,6.9732623,7.5159745,8.058686,8.601398,9.14411,9.686822,9.20658,8.726339,8.246098,7.7658563,7.2856145,8.0040245,8.718531,9.433036,10.147541,10.862047,10.741011,10.61607,10.495033,10.373997,10.249056,10.221725,10.194394,10.167064,10.139732,10.112402,8.535024,6.957645,5.380266,3.802888,2.2255092,2.6588979,3.0883822,3.521771,3.9551594,4.388548,3.9551594,3.521771,3.0883822,2.6588979,2.2255092,2.280171,2.3348327,2.3894942,2.4441557,2.4988174,2.1474214,1.796025,1.4407244,1.0893283,0.737932,1.1088502,1.4836729,1.8545911,2.2294137,2.6003318,8.784905,14.969479,21.15405,27.338625,33.523197,30.454338,27.381573,24.30881,21.236044,18.163279,16.796738,15.434102,14.067561,12.70102,11.338385,10.631687,9.921086,9.21439,8.507692,7.800996,8.382751,8.964508,9.546264,10.131924,10.71368,10.299813,9.885946,9.475985,9.062118,8.648251,9.651682,10.651209,11.650736,12.650263,13.64979,11.100216,8.550641,6.001066,3.4514916,0.9019169,0.80430686,0.7106012,0.61689556,0.5192855,0.42557985,0.37872702,0.3357786,0.28892577,0.24597734,0.19912452,0.9058213,1.6164225,2.3231194,3.0298162,3.736513,3.3616903,2.9829633,2.6042364,2.2294137,1.8506867,2.0810463,2.3153105,2.5456703,2.7799344,3.0141985,2.5808098,2.1474214,1.7140326,1.2806439,0.8511597,1.1439898,1.4407244,1.7335546,2.0302892,2.3231194,2.5183394,2.7096553,2.900971,3.096191,3.2875066,3.3031244,3.3187418,3.3343596,3.3460727,3.3616903,3.638903,3.912211,4.1894236,4.462732,4.73604,4.5837684,4.4314966,4.279225,4.126953,3.9746814,3.6271896,3.279698,2.9322062,2.5847144,2.2372224,2.1786566,2.1161861,2.05762,1.999054,1.9365835,2.0341935,2.1278992,2.2216048,2.3192148,2.4129205,2.5612879,2.7135596,2.8619268,3.0141985,3.1625657,2.854118,2.541766,2.233318,1.9209659,1.6125181,1.5812829,1.5539521,1.5227169,1.4914817,1.4641509,1.4719596,1.4836729,1.4914817,1.5031948,1.5110037,1.6359446,1.756981,1.8819219,2.0029583,2.1239948,2.1083772,2.096664,2.0810463,2.0654287,2.0498111,1.9443923,1.8350691,1.7257458,1.620327,1.5110037,1.2650263,1.0190489,0.76916724,0.5231899,0.27330816,0.6559396,1.038571,1.4212024,1.8038338,2.1864653,2.1435168,2.096664,2.0537157,2.0068626,1.9639144,2.2372224,2.514435,2.787743,3.0610514,3.338264,3.193801,3.0532427,2.9087796,2.7682211,2.6237583,2.1981785,1.7686942,1.3431144,0.9136301,0.48805028,0.77307165,1.0619974,1.3509232,1.6359446,1.9248703,2.397303,2.8697357,3.3421683,3.814601,4.2870336,3.7130866,3.1391394,2.5612879,1.9873407,1.4133936,1.3235924,1.2376955,1.1517987,1.0619974,0.97610056,0.8511597,0.7301232,0.60908675,0.48414588,0.3631094,0.339683,0.31625658,0.29673457,0.27330816,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.113227665,0.22645533,0.3357786,0.44900626,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.14055848,0.28111696,0.42167544,0.5583295,0.698888,0.5661383,0.42948425,0.29673457,0.16008049,0.023426414,0.15617609,0.28502136,0.41386664,0.5466163,0.6754616,0.5388075,0.40605783,0.26940376,0.13665408,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5700427,1.1400855,1.7101282,2.280171,2.8502135,2.822883,2.795552,2.7682211,2.7408905,2.7135596,2.3621633,2.0107672,1.6632754,1.3118792,0.96438736,1.3860629,1.8077383,2.2294137,2.6510892,3.076669,2.979059,2.8814487,2.7838387,2.6862288,2.5886188,2.7291772,2.87364,3.0141985,3.1586614,3.2992198,3.6506162,3.998108,4.349504,4.7009,5.0483923,5.4895897,5.930787,6.36808,6.8092775,7.250475,6.9810715,6.7116675,6.4383593,6.168956,5.899552,6.153338,6.4110284,6.6648145,6.918601,7.1762915,8.976221,10.780055,12.583888,14.383818,16.187653,15.441911,14.69617,13.954333,13.208592,12.4628525,12.236397,12.013845,11.787391,11.560935,11.338385,10.073358,8.812236,7.551114,6.2860875,5.024966,5.1186714,5.2162814,5.309987,5.4036927,5.5013027,5.0718184,4.6384296,4.2089458,3.7794614,3.349977,3.959064,4.5681505,5.181142,5.7902284,6.3993154,6.141625,5.883934,5.6262436,5.368553,5.1108627,4.552533,3.9942036,3.4319696,2.87364,2.3114061,2.2255092,2.135708,2.0498111,1.9639144,1.8741131,1.893635,1.9131571,1.9365835,1.9561055,1.9756275,2.3543546,2.736986,3.1157131,3.49444,3.873167,3.6662338,3.4593005,3.252367,3.0454338,2.8385005,2.9087796,2.979059,3.049338,3.1157131,3.1859922,3.0727646,2.9556324,2.8424048,2.7291772,2.612045,2.436347,2.260649,2.0888553,1.9131571,1.737459,1.6281357,1.5188124,1.4055848,1.2962615,1.1869383,0.3513962,0.3435874,0.339683,0.3357786,0.3318742,0.3240654,0.31625658,0.30454338,0.29673457,0.28502136,0.27330816,0.28892577,0.30454338,0.32016098,0.3357786,0.3513962,0.3631094,0.37482262,0.38653582,0.39824903,0.41386664,0.38653582,0.359205,0.3318742,0.30063897,0.27330816,0.29673457,0.31625658,0.3357786,0.3553006,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.45291066,0.5309987,0.60908675,0.6832704,0.76135844,0.74574083,0.7340276,0.71841,0.7027924,0.6871748,0.7066968,0.7262188,0.74574083,0.76916724,0.78868926,0.8394465,0.8862993,0.93705654,0.9878138,1.038571,1.0737107,1.1088502,1.1439898,1.1791295,1.2142692,1.0893283,0.96438736,0.8394465,0.7106012,0.58566034,0.5661383,0.5427119,0.5192855,0.4958591,0.47633708,0.39434463,0.31625658,0.23426414,0.15617609,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.57394713,1.1517987,1.7257458,2.2996929,2.87364,5.5989127,8.320281,11.04165,13.766922,16.48829,13.6693125,10.84643,8.027451,5.2084727,2.3855898,3.6349986,4.8805027,6.1299114,7.37932,8.624825,7.629202,6.629675,5.6340523,4.6345253,3.638903,3.0532427,2.4675822,1.8819219,1.2962615,0.7106012,0.79649806,0.8784905,0.96048295,1.0424755,1.1244678,1.4836729,1.8389735,2.1981785,2.5534792,2.912684,3.2718892,3.631094,3.9942036,4.3534083,4.7126136,4.747753,4.7828927,4.8180323,4.853172,4.8883114,4.716518,4.5408196,4.369026,4.1972322,4.025439,3.873167,3.7208953,3.5686235,3.416352,3.2640803,3.0805733,2.900971,2.7213683,2.541766,2.3621633,2.1474214,1.9326792,1.717937,1.5031948,1.2884527,1.3509232,1.4172981,1.4836729,1.5461433,1.6125181,1.7725986,1.9326792,2.0927596,2.25284,2.4129205,2.4246337,2.436347,2.4480603,2.463678,2.475391,3.8614538,5.251421,6.6374836,8.023546,9.413514,8.054782,6.6960497,5.3412223,3.9824903,2.6237583,2.690133,2.7565079,2.8189783,2.8853533,2.951728,3.6662338,4.3846436,5.1030536,5.8214636,6.5359693,6.7975645,7.0591593,7.3168497,7.578445,7.8361354,7.578445,7.320754,7.0630636,6.8092775,6.551587,6.617962,6.6843367,6.7507114,6.8209906,6.8873653,7.297328,7.70729,8.117252,8.527214,8.937177,8.6131115,8.292951,7.968885,7.648724,7.3246584,7.918128,8.511597,9.101162,9.694631,10.2881,10.280292,10.272482,10.264673,10.256865,10.249056,10.432563,10.61607,10.795672,10.979179,11.162686,9.694631,8.226576,6.75852,5.2943697,3.8263142,4.2284675,4.630621,5.0327744,5.434928,5.8370814,5.2475166,4.657952,4.068387,3.4788225,2.8892577,2.7604125,2.631567,2.5066261,2.377781,2.2489357,1.9951496,1.7413634,1.4836729,1.2298868,0.97610056,1.2455044,1.5149081,1.7843118,2.0537157,2.3231194,7.843944,13.364769,18.885593,24.406418,29.92334,29.040943,28.158548,27.276154,26.393759,25.511364,23.231194,20.951023,18.67085,16.39068,14.114414,13.4740925,12.83377,12.193448,11.553126,10.912805,11.701493,12.494087,13.282777,14.0714655,14.864059,13.189071,11.514082,9.839094,8.164105,6.4891167,7.238762,7.988407,8.738052,9.487698,10.237343,8.324185,6.4110284,4.5017757,2.5886188,0.6754616,0.7106012,0.74574083,0.78088045,0.8160201,0.8511597,0.76135844,0.6715572,0.58175594,0.48805028,0.39824903,1.038571,1.678893,2.3192148,2.959537,3.5998588,3.2836022,2.9634414,2.6471848,2.330928,2.0107672,2.4285383,2.8424048,3.2562714,3.6740425,4.087909,3.533484,2.9829633,2.4285383,1.8780174,1.3235924,1.5149081,1.7062237,1.893635,2.084951,2.2762666,2.6081407,2.9439192,3.279698,3.6154766,3.951255,3.9668727,3.9863946,4.0020123,4.0215344,4.037152,4.21285,4.388548,4.564246,4.73604,4.911738,4.732136,4.552533,4.3729305,4.193328,4.0137253,3.6545205,3.2992198,2.9400148,2.5808098,2.2255092,2.1669433,2.1083772,2.0537157,1.9951496,1.9365835,1.9287747,1.9170616,1.9092526,1.8975395,1.8858263,2.0498111,2.2137961,2.3738766,2.5378613,2.7018464,2.416825,2.135708,1.8506867,1.5695697,1.2884527,1.3665408,1.4407244,1.5188124,1.5969005,1.6749885,1.6593709,1.639849,1.6242313,1.6047094,1.5890918,1.6827974,1.7765031,1.8741131,1.9678187,2.0615244,2.1318035,2.2020829,2.2723622,2.3426414,2.4129205,2.2840753,2.1591344,2.0302892,1.901444,1.7765031,1.5305257,1.2845483,1.038571,0.79649806,0.5505207,0.8784905,1.2064602,1.53443,1.8584955,2.1864653,2.1083772,2.0341935,1.9561055,1.8780174,1.7999294,2.0380979,2.2762666,2.514435,2.7486992,2.9868677,2.815074,2.6432803,2.4714866,2.2957885,2.1239948,1.8077383,1.4914817,1.1713207,0.8550641,0.5388075,0.81211567,1.0893283,1.3626363,1.6359446,1.9131571,2.4441557,2.979059,3.5100577,4.041056,4.575959,3.9746814,3.3734035,2.77603,2.174752,1.5734742,1.43682,1.3001659,1.1635119,1.0268579,0.8862993,0.8550641,0.8238289,0.78868926,0.75745404,0.7262188,0.679366,0.63641757,0.58956474,0.5466163,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.3513962,0.26159495,0.1756981,0.08589685,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.12884527,0.26159495,0.39044023,0.5192855,0.6481308,0.5309987,0.40996224,0.28892577,0.1717937,0.05075723,0.29673457,0.5466163,0.79259366,1.038571,1.2884527,1.0307622,0.77307165,0.5153811,0.25769055,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.8784905,1.7530766,2.631567,3.5100577,4.388548,4.318269,4.251894,4.185519,4.1191444,4.0488653,3.5998588,3.1508527,2.7018464,2.2489357,1.7999294,2.194274,2.5886188,2.9868677,3.3812122,3.775557,3.4671092,3.1586614,2.854118,2.5456703,2.2372224,2.7330816,3.232845,3.7287042,4.2284675,4.7243266,5.2358036,5.7511845,6.262661,6.774138,7.2856145,7.453504,7.621393,7.7892823,7.957172,8.125061,7.8868923,7.6448197,7.406651,7.164578,6.9264097,7.1099167,7.2934237,7.480835,7.6643414,7.8517528,9.019169,10.186585,11.354002,12.521418,13.688834,13.185166,12.681499,12.181735,11.678067,11.174399,11.150972,11.123642,11.100216,11.076789,11.0494585,10.010887,8.976221,7.9376497,6.899079,5.8644123,5.7785153,5.6926184,5.606722,5.520825,5.4388323,4.989826,4.5408196,4.095718,3.6467118,3.2016098,3.5959544,3.9902992,4.3846436,4.7789884,5.173333,5.1460023,5.1186714,5.0913405,5.0640097,5.036679,4.4314966,3.8224099,3.213323,2.6081407,1.999054,2.0380979,2.0732377,2.1122816,2.1513257,2.1864653,2.1786566,2.1669433,2.1591344,2.1474214,2.135708,2.3465457,2.5573835,2.7682211,2.979059,3.1859922,3.1235218,3.057147,2.9907722,2.9283018,2.8619268,2.951728,3.0415294,3.1313305,3.2211318,3.310933,3.2562714,3.2016098,3.1469483,3.0922866,3.0376248,2.77603,2.5105307,2.2489357,1.9873407,1.7257458,1.6164225,1.5110037,1.4016805,1.2962615,1.1869383,0.39824903,0.39434463,0.38653582,0.37872702,0.3709182,0.3631094,0.3474918,0.3318742,0.31625658,0.30063897,0.28892577,0.29673457,0.30844778,0.31625658,0.3279698,0.3357786,0.3513962,0.3631094,0.37482262,0.38653582,0.39824903,0.37872702,0.3553006,0.3318742,0.30844778,0.28892577,0.30454338,0.3240654,0.339683,0.359205,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.43338865,0.4958591,0.5544251,0.61689556,0.6754616,0.6520352,0.62860876,0.60908675,0.58566034,0.5622339,0.62860876,0.698888,0.76526284,0.8316377,0.9019169,0.9878138,1.0737107,1.1635119,1.2494087,1.33921,1.33921,1.3431144,1.3431144,1.3470187,1.3509232,1.2142692,1.0737107,0.93705654,0.80040246,0.6637484,0.6715572,0.6832704,0.6910792,0.7027924,0.7106012,0.58175594,0.44900626,0.31625658,0.1835069,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.737932,1.475864,2.2137961,2.951728,3.6857557,5.5169206,7.3441806,9.171441,10.998701,12.825961,10.6590185,8.488171,6.321227,4.154284,1.9873407,2.7408905,3.4905357,4.2440853,4.997635,5.7511845,5.1225758,4.493967,3.8692627,3.240654,2.612045,2.1864653,1.756981,1.3314011,0.9019169,0.47633708,0.6559396,0.8355421,1.0151446,1.1947471,1.3743496,1.678893,1.9834363,2.2918842,2.5964274,2.900971,3.1781836,3.455396,3.7326086,4.009821,4.2870336,4.365122,4.4432096,4.521298,4.5993857,4.6735697,4.5837684,4.493967,4.4041657,4.3143644,4.224563,4.2011366,4.181615,4.1581883,4.134762,4.1113358,3.9551594,3.7989833,3.638903,3.4827268,3.3265507,2.9400148,2.5534792,2.1708477,1.7843118,1.4016805,1.4485333,1.4953861,1.542239,1.5890918,1.6359446,1.8038338,1.9678187,2.1318035,2.2957885,2.463678,2.5261483,2.5886188,2.6510892,2.7135596,2.77603,3.998108,5.22409,6.4500723,7.676055,8.898132,7.656533,6.4149327,5.173333,3.9317331,2.6862288,2.8345962,2.9829633,3.1313305,3.2757936,3.4241607,4.2440853,5.0640097,5.883934,6.703859,7.523783,7.465217,7.406651,7.3441806,7.2856145,7.223144,6.969358,6.715572,6.461786,6.2040954,5.950309,6.1181984,6.289992,6.461786,6.629675,6.801469,7.0786815,7.355894,7.633106,7.910319,8.187531,8.023546,7.8556576,7.6916723,7.5276875,7.363703,7.832231,8.300759,8.773191,9.24172,9.714153,9.8195715,9.928895,10.034314,10.143637,10.249056,10.6434,11.033841,11.428185,11.818625,12.212971,10.8542385,9.499411,8.140678,6.7819467,5.423215,5.7980375,6.168956,6.5437784,6.914696,7.2856145,6.5398736,5.794133,5.044488,4.298747,3.5491016,3.240654,2.9283018,2.619854,2.3114061,1.999054,1.8428779,1.6867018,1.5266213,1.3704453,1.2142692,1.3782539,1.5461433,1.7140326,1.8819219,2.0498111,6.902983,11.760059,16.613232,21.470308,26.32348,27.631454,28.93943,30.247404,31.55538,32.863354,29.665648,26.471848,23.278046,20.084246,16.88654,16.316498,15.74255,15.168603,14.59856,14.024612,15.024139,16.019762,17.019289,18.014912,19.010534,16.074425,13.138313,10.198298,7.262188,4.3260775,4.825841,5.3256044,5.825368,6.3251314,6.824895,5.548156,4.2753205,2.998581,1.7257458,0.44900626,0.61689556,0.78088045,0.94486535,1.1088502,1.2767396,1.1400855,1.0034313,0.8706817,0.7340276,0.60127795,1.1713207,1.7452679,2.3192148,2.8892577,3.4632049,3.2055142,2.9478238,2.690133,2.4324427,2.174752,2.7721257,3.3694992,3.9668727,4.564246,5.1616197,4.4900627,3.8185053,3.1430438,2.4714866,1.7999294,1.8858263,1.9717231,2.0537157,2.1396124,2.2255092,2.7018464,3.1781836,3.6584249,4.134762,4.6110992,4.630621,4.6540475,4.6735697,4.6930914,4.7126136,4.786797,4.860981,4.939069,5.0132523,5.087436,4.8805027,4.6735697,4.466636,4.2557983,4.0488653,3.6818514,3.3148375,2.9478238,2.5808098,2.2137961,2.1591344,2.1005683,2.0459068,1.9912452,1.9365835,1.8233559,1.7062237,1.5929961,1.475864,1.3626363,1.5383345,1.7140326,1.8858263,2.0615244,2.2372224,1.9834363,1.7257458,1.4719596,1.2181735,0.96438736,1.1478943,1.3314011,1.5188124,1.7023194,1.8858263,1.8428779,1.796025,1.7530766,1.7062237,1.6632754,1.7296503,1.796025,1.8663043,1.9326792,1.999054,2.15523,2.3114061,2.463678,2.619854,2.77603,2.6276627,2.4792955,2.330928,2.1864653,2.0380979,1.796025,1.5539521,1.3118792,1.0659018,0.8238289,1.097137,1.3704453,1.6437533,1.9131571,2.1864653,2.077142,1.9678187,1.8584955,1.7491722,1.6359446,1.8389735,2.0380979,2.2372224,2.436347,2.639376,2.436347,2.233318,2.0302892,1.8272603,1.6242313,1.4172981,1.2103647,1.0034313,0.79649806,0.58566034,0.8511597,1.1127546,1.3743496,1.6359446,1.901444,2.4910088,3.084478,3.677947,4.271416,4.860981,4.2362766,3.611572,2.9868677,2.3621633,1.737459,1.5500476,1.3626363,1.175225,0.9878138,0.80040246,0.8589685,0.9136301,0.97219616,1.0307622,1.0893283,1.0190489,0.95267415,0.8862993,0.8160201,0.74964523,0.60127795,0.44900626,0.30063897,0.14836729,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.12103647,0.23816854,0.359205,0.48024148,0.60127795,0.4958591,0.39044023,0.28502136,0.1796025,0.07418364,0.44119745,0.80430686,1.1713207,1.53443,1.901444,1.5188124,1.1400855,0.76135844,0.37872702,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1869383,2.3699722,3.5569105,4.7399445,5.9268827,5.8175592,5.708236,5.602817,5.493494,5.388075,4.8375545,4.2870336,3.736513,3.1859922,2.639376,3.0063896,3.3734035,3.7404175,4.1074314,4.474445,3.959064,3.4397783,2.9243972,2.4051118,1.8858263,2.7408905,3.59205,4.4432096,5.298274,6.1494336,6.824895,7.5003567,8.175818,8.85128,9.526741,9.421323,9.315904,9.2104845,9.105066,8.999647,8.78881,8.581876,8.371038,8.160201,7.9493628,8.066495,8.179723,8.296855,8.410083,8.52331,9.058213,9.589212,10.124115,10.655114,11.186112,10.928422,10.666827,10.409137,10.147541,9.885946,10.061645,10.237343,10.413041,10.588739,10.764437,9.948417,9.136301,8.324185,7.5120697,6.699954,6.434455,6.168956,5.903456,5.6418614,5.376362,4.911738,4.4432096,3.978586,3.513962,3.049338,3.2289407,3.408543,3.5881457,3.7716527,3.951255,4.154284,4.3534083,4.5564375,4.759466,4.9624953,4.3065557,3.6506162,2.998581,2.3426414,1.6867018,1.8506867,2.0107672,2.174752,2.338737,2.4988174,2.4597735,2.4207294,2.3816853,2.338737,2.2996929,2.338737,2.3816853,2.4207294,2.4597735,2.4988174,2.5769055,2.6549935,2.7330816,2.8111696,2.8892577,2.998581,3.1079042,3.2172275,3.3265507,3.435874,3.4436827,3.4475873,3.4514916,3.4593005,3.4632049,3.1118085,2.7643168,2.4129205,2.0615244,1.7140326,1.6086137,1.5031948,1.397776,1.2923572,1.1869383,0.44900626,0.44119745,0.42948425,0.42167544,0.40996224,0.39824903,0.37872702,0.359205,0.339683,0.32016098,0.30063897,0.30454338,0.30844778,0.31625658,0.32016098,0.3240654,0.3357786,0.3513962,0.3631094,0.37482262,0.38653582,0.3709182,0.3513962,0.3357786,0.31625658,0.30063897,0.31625658,0.3318742,0.3435874,0.359205,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.41777104,0.46071947,0.5036679,0.5466163,0.58566034,0.5583295,0.5270943,0.4958591,0.46852827,0.43729305,0.5544251,0.6676528,0.78088045,0.8980125,1.0112402,1.1361811,1.261122,1.3860629,1.5110037,1.6359446,1.6086137,1.5773785,1.5461433,1.5188124,1.4875772,1.33921,1.1869383,1.038571,0.8862993,0.737932,0.78088045,0.8238289,0.8667773,0.9058213,0.94876975,0.76526284,0.58175594,0.39434463,0.21083772,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.9019169,1.7999294,2.7018464,3.5998588,4.5017757,5.4310236,6.364176,7.297328,8.23048,9.163632,7.648724,6.133816,4.618908,3.1039999,1.5890918,1.8467822,2.1005683,2.358259,2.6159496,2.87364,2.6159496,2.358259,2.1005683,1.8467822,1.5890918,1.3157835,1.0463798,0.77697605,0.5075723,0.23816854,0.5153811,0.79259366,1.0698062,1.3470187,1.6242313,1.8780174,2.1318035,2.3816853,2.6354716,2.8892577,3.0805733,3.2757936,3.4710135,3.6662338,3.8614538,3.9824903,4.1035266,4.220659,4.3416953,4.462732,4.454923,4.447114,4.4393053,4.4314966,4.423688,4.533011,4.6384296,4.747753,4.853172,4.9624953,4.825841,4.6930914,4.5564375,4.423688,4.2870336,3.7326086,3.1781836,2.6237583,2.069333,1.5110037,1.542239,1.5734742,1.6008049,1.6320401,1.6632754,1.8311646,2.0029583,2.1708477,2.3426414,2.514435,2.6237583,2.736986,2.8502135,2.9634414,3.076669,4.138666,5.2006636,6.262661,7.3246584,8.386656,7.2582836,6.133816,5.0054436,3.8770714,2.7486992,2.979059,3.2094188,3.4397783,3.6701381,3.900498,4.8219366,5.743376,6.6687193,7.590158,8.511597,8.13287,7.7541428,7.3715115,6.9927845,6.6140575,6.3602715,6.1064854,5.8566036,5.602817,5.349031,5.6223392,5.8956475,6.168956,6.4383593,6.7116675,6.8561306,7.000593,7.1489606,7.2934237,7.437886,7.4300776,7.422269,7.4144597,7.406651,7.3988423,7.746334,8.093826,8.441318,8.78881,9.136301,9.358852,9.581403,9.803954,10.0265045,10.249056,10.8542385,11.455516,12.056794,12.658072,13.263254,12.013845,10.768341,9.518932,8.273428,7.0240197,7.367607,7.7111945,8.050878,8.3944645,8.738052,7.832231,6.9264097,6.0205884,5.1186714,4.21285,3.7208953,3.2289407,2.7330816,2.241127,1.7491722,1.6906061,1.6281357,1.5695697,1.5110037,1.4485333,1.5149081,1.5812829,1.6437533,1.7101282,1.7765031,5.9659266,10.155351,14.344774,18.534197,22.723621,26.221966,29.72031,33.218655,36.713093,40.211437,36.104008,31.992672,27.881336,23.773905,19.662569,19.158901,18.651329,18.147661,17.643993,17.136421,18.342882,19.549341,20.751898,21.958359,23.160913,18.963682,14.762545,10.561408,6.364176,2.1630387,2.4129205,2.6628022,2.912684,3.1625657,3.4124475,2.77603,2.135708,1.4992905,0.8628729,0.22645533,0.5192855,0.8160201,1.1088502,1.4055848,1.698415,1.5188124,1.33921,1.1596074,0.98000497,0.80040246,1.3040704,1.8116426,2.3153105,2.8189783,3.3265507,3.1274261,2.9283018,2.7330816,2.533957,2.338737,3.1157131,3.8965936,4.677474,5.4583545,6.239235,5.446641,4.6540475,3.8614538,3.06886,2.2762666,2.2567444,2.233318,2.2137961,2.194274,2.174752,2.795552,3.416352,4.0332475,4.6540475,5.2748475,5.298274,5.3217,5.3412223,5.364649,5.388075,5.3607445,5.337318,5.3138914,5.2865605,5.263134,5.02887,4.7907014,4.5564375,4.322173,4.087909,3.7091823,3.3343596,2.9556324,2.5769055,2.1981785,2.1474214,2.096664,2.0420024,1.9912452,1.9365835,1.717937,1.4992905,1.2767396,1.0580931,0.8394465,1.0268579,1.2142692,1.4016805,1.5890918,1.7765031,1.5461433,1.319688,1.0932326,0.8667773,0.63641757,0.92924774,1.2220778,1.5149081,1.8077383,2.1005683,2.0263848,1.9561055,1.8819219,1.8116426,1.737459,1.7765031,1.815547,1.8584955,1.8975395,1.9365835,2.1786566,2.416825,2.6588979,2.8970666,3.1391394,2.97125,2.803361,2.6354716,2.4675822,2.2996929,2.0615244,1.8194515,1.5812829,1.33921,1.1010414,1.3157835,1.53443,1.7530766,1.9717231,2.1864653,2.0459068,1.901444,1.7608855,1.6164225,1.475864,1.6359446,1.7999294,1.9639144,2.1239948,2.2879796,2.0537157,1.8233559,1.5890918,1.358732,1.1244678,1.0268579,0.92924774,0.8316377,0.7340276,0.63641757,0.8862993,1.1361811,1.3860629,1.6359446,1.8858263,2.541766,3.193801,3.8458362,4.4978714,5.1499066,4.5017757,3.8497405,3.2016098,2.5495746,1.901444,1.6632754,1.4251068,1.1869383,0.94876975,0.7106012,0.8589685,1.0073358,1.1557031,1.3040704,1.4485333,1.358732,1.2689307,1.1791295,1.0893283,0.999527,0.80040246,0.60127795,0.39824903,0.19912452,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.10932326,0.21864653,0.3318742,0.44119745,0.5505207,0.46071947,0.3709182,0.28111696,0.19131571,0.10151446,0.58175594,1.0659018,1.5461433,2.0302892,2.514435,2.0107672,1.5070993,1.0034313,0.5036679,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.4914817,2.9868677,4.478349,5.969831,7.461313,7.3168497,7.168483,7.0201154,6.871748,6.7233806,6.0752497,5.423215,4.775084,4.123049,3.474918,3.814601,4.154284,4.493967,4.83365,5.173333,4.447114,3.7208953,2.9907722,2.2645533,1.5383345,2.7447948,3.951255,5.1616197,6.36808,7.57454,8.413987,9.249529,10.088976,10.924518,11.763964,11.385237,11.00651,10.631687,10.25296,9.874233,9.694631,9.515028,9.335425,9.155824,8.976221,9.019169,9.066022,9.108971,9.155824,9.198771,9.097258,8.995743,8.894228,8.78881,8.687295,8.671678,8.652155,8.636538,8.617016,8.601398,8.976221,9.351044,9.725866,10.100689,10.475512,9.885946,9.300286,8.710721,8.125061,7.5394006,7.094299,6.649197,6.2040954,5.758993,5.3138914,4.829746,4.3455997,3.8653584,3.3812122,2.900971,2.8658314,2.8306916,2.795552,2.7604125,2.7252727,3.1586614,3.5881457,4.0215344,4.454923,4.8883114,4.185519,3.4827268,2.7799344,2.077142,1.3743496,1.6632754,1.9482968,2.2372224,2.5261483,2.8111696,2.7408905,2.6706111,2.6042364,2.533957,2.463678,2.330928,2.2020829,2.0732377,1.9443923,1.8116426,2.0341935,2.25284,2.4714866,2.6940374,2.912684,3.0415294,3.174279,3.3031244,3.4319696,3.5608149,3.6271896,3.6935644,3.7560349,3.8224099,3.8887846,3.4514916,3.0141985,2.5769055,2.135708,1.698415,1.5969005,1.4953861,1.3938715,1.2884527,1.1869383,0.4997635,0.48805028,0.47633708,0.46071947,0.44900626,0.43729305,0.41386664,0.38653582,0.3631094,0.3357786,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.3240654,0.3357786,0.3513962,0.3631094,0.37482262,0.3631094,0.3513962,0.3357786,0.3240654,0.31235218,0.3240654,0.3357786,0.3513962,0.3631094,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.39824903,0.42557985,0.44900626,0.47633708,0.4997635,0.46071947,0.42557985,0.38653582,0.3513962,0.31235218,0.47633708,0.63641757,0.80040246,0.96438736,1.1244678,1.2884527,1.4485333,1.6125181,1.7765031,1.9365835,1.8741131,1.8116426,1.7491722,1.6867018,1.6242313,1.4641509,1.3001659,1.1361811,0.97610056,0.81211567,0.8862993,0.96438736,1.038571,1.1127546,1.1869383,0.94876975,0.7106012,0.47633708,0.23816854,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0619974,2.1239948,3.1859922,4.251894,5.3138914,5.349031,5.388075,5.423215,5.462259,5.5013027,4.6384296,3.775557,2.912684,2.0498111,1.1869383,0.94876975,0.7106012,0.47633708,0.23816854,0.0,0.113227665,0.22645533,0.3357786,0.44900626,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.37482262,0.74964523,1.1244678,1.4992905,1.8741131,2.0732377,2.2762666,2.475391,2.6745155,2.87364,2.9868677,3.1000953,3.213323,3.3265507,3.435874,3.5998588,3.7638438,3.9239242,4.087909,4.251894,4.3260775,4.4002614,4.474445,4.548629,4.6267166,4.860981,5.099149,5.337318,5.575486,5.813655,5.700427,5.5871997,5.473972,5.3607445,5.251421,4.5252023,3.7989833,3.076669,2.35045,1.6242313,1.6359446,1.6515622,1.6632754,1.6749885,1.6867018,1.8623998,2.0380979,2.2137961,2.3855898,2.5612879,2.7252727,2.8892577,3.049338,3.213323,3.3734035,4.2753205,5.173333,6.0752497,6.9732623,7.8751793,6.8639393,5.8487945,4.8375545,3.8263142,2.8111696,3.1235218,3.435874,3.7482262,4.0605783,4.376835,5.3997884,6.426646,7.4495993,8.476458,9.499411,8.800523,8.101635,7.3988423,6.699954,6.001066,5.7511845,5.5013027,5.251421,5.001539,4.7516575,5.12648,5.5013027,5.8761253,6.250948,6.6257706,6.6374836,6.649197,6.66091,6.676528,6.688241,6.8366084,6.98888,7.137247,7.2856145,7.437886,7.6643414,7.8868923,8.113348,8.335898,8.562354,8.898132,9.237816,9.573594,9.913278,10.249056,11.061172,11.873287,12.689307,13.501423,14.313539,13.173453,12.037272,10.901091,9.761005,8.624825,8.937177,9.249529,9.561881,9.874233,10.186585,9.124588,8.062591,7.000593,5.938596,4.8765984,4.2011366,3.5256753,2.8502135,2.174752,1.4992905,1.5383345,1.5734742,1.6125181,1.6515622,1.6867018,1.6515622,1.6125181,1.5734742,1.5383345,1.4992905,5.024966,8.550641,12.076316,15.601992,19.123762,24.812477,30.50119,36.186,41.874714,47.563427,42.538464,37.513496,32.488533,27.463566,22.4386,22.001307,21.564014,21.12672,20.689428,20.24823,21.661623,23.075018,24.48841,25.901804,27.311295,21.849035,16.386776,10.924518,5.462259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.42557985,0.8511597,1.2767396,1.698415,2.1239948,1.901444,1.6749885,1.4485333,1.2259823,0.999527,1.43682,1.8741131,2.3114061,2.7486992,3.1859922,3.049338,2.912684,2.77603,2.639376,2.4988174,3.4632049,4.423688,5.388075,6.348558,7.3129454,6.3993154,5.4856853,4.575959,3.6623292,2.7486992,2.6237583,2.4988174,2.3738766,2.2489357,2.1239948,2.8892577,3.6506162,4.4119744,5.173333,5.938596,5.9620223,5.989353,6.012779,6.036206,6.0635366,5.938596,5.813655,5.688714,5.563773,5.4388323,5.173333,4.911738,4.650143,4.388548,4.123049,3.736513,3.349977,2.9634414,2.5769055,2.1864653,2.135708,2.0888553,2.0380979,1.9873407,1.9365835,1.6125181,1.2884527,0.96438736,0.63641757,0.31235218,0.5114767,0.7106012,0.9136301,1.1127546,1.3118792,1.1127546,0.9136301,0.7106012,0.5114767,0.31235218,0.7106012,1.1127546,1.5110037,1.9131571,2.3114061,2.2137961,2.1122816,2.0107672,1.9131571,1.8116426,1.8233559,1.8389735,1.8506867,1.8623998,1.8741131,2.1981785,2.5261483,2.8502135,3.174279,3.4983444,3.310933,3.1235218,2.9361105,2.7486992,2.5612879,2.3231194,2.0888553,1.8506867,1.6125181,1.3743496,1.5383345,1.698415,1.8623998,2.0263848,2.1864653,2.0107672,1.8389735,1.6632754,1.4875772,1.3118792,1.43682,1.5617609,1.6867018,1.8116426,1.9365835,1.6749885,1.4133936,1.1517987,0.8862993,0.62470436,0.63641757,0.6481308,0.6637484,0.6754616,0.6871748,0.92534333,1.1635119,1.4016805,1.6359446,1.8741131,2.5886188,3.2992198,4.0137253,4.7243266,5.4388323,4.7633705,4.087909,3.4124475,2.736986,2.0615244,1.7765031,1.4875772,1.1986516,0.9136301,0.62470436,0.8628729,1.1010414,1.33921,1.5734742,1.8116426,1.698415,1.5890918,1.475864,1.3626363,1.2494087,0.999527,0.74964523,0.4997635,0.24988174,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.42557985,0.3513962,0.27330816,0.19912452,0.12494087,0.7262188,1.3235924,1.9248703,2.5261483,3.1235218,2.4988174,1.8741131,1.2494087,0.62470436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.7999294,3.5998588,5.3997884,7.1997175,8.999647,8.812236,8.624825,8.437413,8.250002,8.062591,7.3129454,6.5633,5.813655,5.0640097,4.3143644,4.6267166,4.939069,5.251421,5.563773,5.8761253,4.939069,3.998108,3.0610514,2.1239948,1.1869383,2.7486992,4.3143644,5.8761253,7.437886,8.999647,9.999174,10.998701,11.998228,13.001659,14.001186,13.349152,12.70102,12.0489855,11.400854,10.748819,10.600452,10.44818,10.299813,10.151445,9.999174,9.975748,9.948417,9.924991,9.901564,9.874233,9.136301,8.398369,7.6643414,6.9264097,6.1884775,6.4110284,6.6374836,6.8639393,7.08649,7.3129454,7.8868923,8.460839,9.0386915,9.612638,10.186585,9.823476,9.464272,9.101162,8.738052,8.374943,7.7502384,7.125534,6.5008297,5.8761253,5.251421,4.7516575,4.2479897,3.7482262,3.2484627,2.7486992,2.4988174,2.2489357,1.999054,1.7491722,1.4992905,2.1630387,2.8267872,3.4866312,4.1503797,4.814128,4.0605783,3.310933,2.5612879,1.8116426,1.0619974,1.475864,1.8858263,2.2996929,2.7135596,3.1235218,3.0259118,2.9243972,2.8267872,2.7252727,2.6237583,2.3231194,2.0263848,1.7257458,1.4251068,1.1244678,1.4875772,1.8506867,2.2137961,2.5769055,2.9361105,3.0883822,3.2367494,3.3890212,3.5373883,3.6857557,3.8106966,3.9356375,4.0605783,4.1894236,4.3143644,3.78727,3.2640803,2.736986,2.2137961,1.6867018,1.5890918,1.4875772,1.3860629,1.2884527,1.1869383,0.5231899,0.5114767,0.4997635,0.48805028,0.47633708,0.46071947,0.44119745,0.41777104,0.39434463,0.3709182,0.3513962,0.3513962,0.3513962,0.3513962,0.3513962,0.3513962,0.359205,0.3631094,0.3709182,0.37872702,0.38653582,0.37872702,0.3670138,0.359205,0.3474918,0.3357786,0.3631094,0.38653582,0.41386664,0.43729305,0.46071947,0.46071947,0.45681506,0.45681506,0.45291066,0.44900626,0.47243267,0.4958591,0.5192855,0.5388075,0.5622339,0.5309987,0.4958591,0.46462387,0.43338865,0.39824903,0.5466163,0.6910792,0.8355421,0.98000497,1.1244678,1.3274968,1.5305257,1.7335546,1.9365835,2.135708,2.1239948,2.1083772,2.0927596,2.077142,2.0615244,1.8311646,1.6008049,1.3743496,1.1439898,0.9136301,0.95657855,1.0034313,1.0463798,1.0932326,1.1361811,0.9097257,0.6832704,0.45681506,0.22645533,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.92924774,1.8545911,2.7838387,3.7091823,4.6384296,4.591577,4.5408196,4.493967,4.447114,4.4002614,3.7091823,3.018103,2.330928,1.639849,0.94876975,0.76135844,0.5700427,0.37872702,0.19131571,0.0,0.093705654,0.19131571,0.28502136,0.37872702,0.47633708,0.48024148,0.48414588,0.48805028,0.4958591,0.4997635,0.75354964,1.0112402,1.2650263,1.5188124,1.7765031,1.9678187,2.1591344,2.3543546,2.5456703,2.736986,2.8189783,2.8970666,2.979059,3.057147,3.1391394,3.3694992,3.6037633,3.8341231,4.068387,4.298747,4.298747,4.298747,4.298747,4.298747,4.298747,4.548629,4.794606,5.040583,5.290465,5.5364423,5.466163,5.3919797,5.3217,5.2475166,5.173333,4.5369153,3.900498,3.2640803,2.6237583,1.9873407,2.1005683,2.2177005,2.330928,2.4480603,2.5612879,2.5300527,2.4988174,2.463678,2.4324427,2.4012074,2.5105307,2.619854,2.7291772,2.8385005,2.951728,3.7443218,4.5408196,5.3334136,6.1299114,6.9264097,6.0908675,5.2553253,4.4197836,3.5842414,2.7486992,2.9868677,3.2211318,3.455396,3.68966,3.9239242,4.825841,5.7316628,6.6335793,7.535496,8.437413,7.8634663,7.2856145,6.7116675,6.13772,5.563773,5.3607445,5.1616197,4.9624953,4.7633705,4.564246,4.841459,5.1186714,5.395884,5.6730967,5.950309,6.1025805,6.2548523,6.407124,6.559396,6.7116675,6.89127,7.066968,7.2465706,7.422269,7.601871,7.7619514,7.9259367,8.086017,8.250002,8.413987,8.710721,9.007456,9.304191,9.600925,9.901564,10.592644,11.283723,11.978706,12.6697855,13.360865,12.294963,11.229061,10.159255,9.093353,8.023546,8.371038,8.718531,9.066022,9.413514,9.761005,8.81614,7.871275,6.9264097,5.9815445,5.036679,4.3534083,3.6662338,2.9829633,2.2957885,1.6125181,1.6086137,1.6008049,1.5969005,1.5929961,1.5890918,1.5656652,1.5461433,1.5266213,1.5070993,1.4875772,4.3026514,7.1177254,9.932799,12.747873,15.562947,20.615244,25.66754,30.719837,35.772133,40.82443,37.673576,34.52663,31.375776,28.224924,25.074072,26.393759,27.713448,29.033134,30.356728,31.676416,29.938957,28.201498,26.464039,24.72658,22.98912,18.389734,13.794253,9.194867,4.5954814,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.39434463,0.78868926,1.1869383,1.5812829,1.9756275,1.7765031,1.5734742,1.3743496,1.175225,0.97610056,1.5656652,2.15523,2.7447948,3.3343596,3.9239242,3.9434462,3.9668727,3.9863946,4.0059166,4.025439,4.884407,5.743376,6.606249,7.465217,8.324185,8.226576,8.125061,8.023546,7.9259367,7.824422,7.336372,6.8483214,6.364176,5.8761253,5.388075,5.8800297,6.3719845,6.8639393,7.355894,7.8517528,7.5979667,7.3441806,7.094299,6.8405128,6.5867267,6.3719845,6.1572423,5.9425,5.727758,5.5130157,5.1186714,4.7243266,4.3260775,3.9317331,3.5373883,3.3070288,3.076669,2.8463092,2.6159496,2.3855898,2.3855898,2.3855898,2.3855898,2.3855898,2.3855898,2.260649,2.135708,2.0107672,1.8858263,1.7608855,1.698415,1.6359446,1.5734742,1.5110037,1.4485333,1.2572175,1.0659018,0.8706817,0.679366,0.48805028,0.98390937,1.4836729,1.979532,2.4792955,2.9751544,2.8072653,2.639376,2.4714866,2.3035975,2.135708,2.0380979,1.9443923,1.8467822,1.7491722,1.6515622,2.0146716,2.3816853,2.7447948,3.1118085,3.474918,3.2250361,2.9751544,2.7252727,2.475391,2.2255092,2.0380979,1.8545911,1.6710842,1.4836729,1.3001659,1.53443,1.7647898,1.999054,2.2294137,2.463678,2.1903696,1.9170616,1.6437533,1.3743496,1.1010414,1.358732,1.620327,1.8819219,2.1396124,2.4012074,2.1044729,1.8116426,1.5149081,1.2181735,0.92534333,0.9136301,0.9058213,0.8941081,0.8862993,0.8745861,1.1322767,1.3899672,1.6476578,1.9053483,2.1630387,2.7018464,3.240654,3.7833657,4.322173,4.860981,4.3455997,3.8263142,3.310933,2.7916477,2.2762666,1.9209659,1.5695697,1.2181735,0.8667773,0.5114767,0.7106012,0.9058213,1.1049459,1.3040704,1.4992905,1.475864,1.4485333,1.4251068,1.4016805,1.3743496,1.6125181,1.8506867,2.0888553,2.3231194,2.5612879,2.0498111,1.5383345,1.0268579,0.5114767,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.015617609,0.015617609,0.019522011,0.023426414,0.023426414,0.03513962,0.046852827,0.05466163,0.06637484,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,0.3631094,0.3318742,0.29673457,0.26159495,0.22645533,0.7145056,1.2064602,1.6945106,2.1864653,2.6745155,2.5456703,2.416825,2.2840753,2.15523,2.0263848,1.7491722,1.4719596,1.1908426,0.9136301,0.63641757,0.5192855,0.40215343,0.28502136,0.1678893,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.5149081,3.0298162,4.5447245,6.0596323,7.57454,7.590158,7.605776,7.621393,7.633106,7.648724,7.461313,7.2739015,7.08649,6.899079,6.7116675,6.9537406,7.195813,7.4417906,7.6838636,7.9259367,6.7663293,5.610626,4.4510183,3.2953155,2.135708,3.506153,4.8765984,6.2470436,7.617489,8.987934,10.069453,11.150972,12.236397,13.317916,14.399435,13.602938,12.806439,12.006037,11.209538,10.413041,10.034314,9.651682,9.272955,8.894228,8.511597,8.453031,8.39056,8.331994,8.273428,8.210958,7.617489,7.0240197,6.426646,5.833177,5.2358036,5.45445,5.6730967,5.891743,6.1064854,6.3251314,6.9068875,7.4886436,8.074304,8.65606,9.237816,8.761478,8.281238,7.8049,7.328563,6.8483214,6.46569,6.0791545,5.6965227,5.309987,4.9234514,4.5993857,4.2753205,3.951255,3.6232853,3.2992198,3.084478,2.8697357,2.6549935,2.4402514,2.2255092,2.736986,3.2484627,3.7638438,4.2753205,4.786797,4.1620927,3.5373883,2.912684,2.2879796,1.6632754,1.9482968,2.2372224,2.5261483,2.8111696,3.1000953,2.97125,2.8385005,2.7096553,2.5808098,2.4480603,2.2216048,1.9912452,1.7608855,1.5305257,1.3001659,1.6242313,1.9482968,2.2762666,2.6003318,2.9243972,3.096191,3.2640803,3.435874,3.6037633,3.775557,3.7794614,3.7833657,3.7911747,3.795079,3.7989833,3.3655949,2.9361105,2.5027218,2.069333,1.6359446,1.5969005,1.5539521,1.5110037,1.4680552,1.4251068,0.5505207,0.5388075,0.5231899,0.5114767,0.4997635,0.48805028,0.46852827,0.44900626,0.42557985,0.40605783,0.38653582,0.38653582,0.38653582,0.38653582,0.38653582,0.38653582,0.39044023,0.39434463,0.39434463,0.39824903,0.39824903,0.39434463,0.38653582,0.37872702,0.3709182,0.3631094,0.39824903,0.43729305,0.47633708,0.5114767,0.5505207,0.5466163,0.5388075,0.5349031,0.5309987,0.5231899,0.5466163,0.5661383,0.58566034,0.60518235,0.62470436,0.59737355,0.5700427,0.5427119,0.5153811,0.48805028,0.61689556,0.7418364,0.8706817,0.9956226,1.1244678,1.3665408,1.6086137,1.8506867,2.096664,2.338737,2.3699722,2.4012074,2.436347,2.4675822,2.4988174,2.2020829,1.9053483,1.6086137,1.3118792,1.0112402,1.0268579,1.0424755,1.0580931,1.0737107,1.0893283,0.8706817,0.6520352,0.43338865,0.21864653,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.79259366,1.5851873,2.377781,3.1703746,3.9629683,3.8302186,3.697469,3.5647192,3.4319696,3.2992198,2.7838387,2.2645533,1.7491722,1.2298868,0.7106012,0.5700427,0.42557985,0.28502136,0.14055848,0.0,0.078088045,0.15617609,0.23426414,0.30844778,0.38653582,0.5114767,0.63251317,0.75354964,0.8784905,0.999527,1.1361811,1.2689307,1.4055848,1.5383345,1.6749885,1.8584955,2.0459068,2.2294137,2.416825,2.6003318,2.6471848,2.6940374,2.7408905,2.7916477,2.8385005,3.1391394,3.4436827,3.7443218,4.0488653,4.349504,4.2753205,4.2011366,4.123049,4.0488653,3.9746814,4.2323723,4.4900627,4.747753,5.0054436,5.263134,5.2318993,5.196759,5.165524,5.134289,5.099149,4.548629,3.998108,3.4514916,2.900971,2.35045,2.5690966,2.7838387,3.0024853,3.2211318,3.435874,3.1977055,2.9556324,2.717464,2.4792955,2.2372224,2.2957885,2.3543546,2.4090161,2.4675822,2.5261483,3.213323,3.9044023,4.5954814,5.2865605,5.9737353,5.3177958,4.661856,4.0020123,3.3460727,2.6862288,2.8463092,3.0024853,3.1586614,3.3187418,3.474918,4.2557983,5.036679,5.813655,6.5945354,7.375416,6.9264097,6.473499,6.0244927,5.575486,5.12648,4.9742084,4.825841,4.6735697,4.5252023,4.376835,4.5564375,4.73604,4.9156423,5.095245,5.2748475,5.5676775,5.860508,6.153338,6.446168,6.7389984,6.942027,7.1489606,7.3519893,7.558923,7.7619514,7.8634663,7.9610763,8.062591,8.164105,8.261715,8.519405,8.777096,9.034787,9.292478,9.550168,10.124115,10.694158,11.268105,11.838148,12.412095,11.416472,10.416945,9.421323,8.421796,7.426173,7.8088045,8.191436,8.574067,8.956698,9.339331,8.511597,7.6838636,6.8561306,6.028397,5.2006636,4.50568,3.8106966,3.1157131,2.4207294,1.7257458,1.678893,1.6281357,1.5812829,1.53443,1.4875772,1.4836729,1.4836729,1.4797685,1.475864,1.475864,3.5803368,5.6848097,7.7892823,9.893755,11.998228,16.41801,20.83389,25.253674,29.669552,34.089336,32.812595,31.535856,30.263021,28.986282,27.713448,30.790115,33.866787,36.943455,40.02403,43.100697,38.212383,33.324074,28.435762,23.551353,18.663042,14.930434,11.197825,7.465217,3.7326086,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3631094,0.7301232,1.0932326,1.4602464,1.8233559,1.6515622,1.475864,1.3001659,1.1244678,0.94876975,1.6906061,2.436347,3.1781836,3.9200199,4.661856,4.841459,5.017157,5.196759,5.3724575,5.548156,6.3056097,7.0630636,7.824422,8.581876,9.339331,10.049932,10.764437,11.475039,12.185639,12.900145,12.0489855,11.20173,10.350571,9.499411,8.648251,8.870802,9.093353,9.315904,9.538455,9.761005,9.2339115,8.702912,8.171914,7.6409154,7.113821,6.8092775,6.5008297,6.196286,5.891743,5.5871997,5.0601053,4.533011,4.0059166,3.4788225,2.951728,2.8775444,2.803361,2.7330816,2.6588979,2.5886188,2.639376,2.6862288,2.736986,2.787743,2.8385005,2.912684,2.9868677,3.0610514,3.1391394,3.213323,2.8892577,2.5612879,2.2372224,1.9131571,1.5890918,1.4016805,1.2181735,1.0307622,0.8472553,0.6637484,1.2572175,1.8506867,2.4480603,3.0415294,3.638903,3.4007344,3.1664703,2.9322062,2.697942,2.463678,2.2567444,2.0459068,1.8389735,1.6320401,1.4251068,1.8311646,2.233318,2.639376,3.0454338,3.4514916,3.1391394,2.8267872,2.514435,2.1981785,1.8858263,1.7530766,1.6242313,1.4914817,1.358732,1.2259823,1.5266213,1.8311646,2.1318035,2.436347,2.736986,2.366068,1.999054,1.6281357,1.2572175,0.8862993,1.2806439,1.678893,2.0732377,2.4675822,2.8619268,2.533957,2.2059872,1.8819219,1.5539521,1.2259823,1.1908426,1.1596074,1.1283722,1.0932326,1.0619974,1.33921,1.6164225,1.893635,2.1708477,2.4480603,2.8189783,3.1859922,3.5530062,3.9200199,4.2870336,3.9278288,3.5686235,3.2094188,2.8463092,2.4871042,2.069333,1.6515622,1.2337911,0.8160201,0.39824903,0.5583295,0.7145056,0.8706817,1.0307622,1.1869383,1.2494087,1.3118792,1.3743496,1.43682,1.4992905,2.2255092,2.951728,3.6740425,4.4002614,5.12648,4.0996222,3.076669,2.0498111,1.0268579,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.031235218,0.03513962,0.039044023,0.046852827,0.05075723,0.058566034,0.06637484,0.07418364,0.078088045,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.30454338,0.30844778,0.31625658,0.32016098,0.3240654,0.7066968,1.0854238,1.4641509,1.8467822,2.2255092,2.5886188,2.9556324,3.3187418,3.6857557,4.0488653,3.49444,2.9400148,2.3855898,1.8311646,1.2767396,1.038571,0.80430686,0.5700427,0.3357786,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.2298868,2.4597735,3.68966,4.919547,6.1494336,6.36808,6.5867267,6.801469,7.0201154,7.238762,7.6135845,7.988407,8.36323,8.738052,9.112875,9.284669,9.456462,9.628256,9.803954,9.975748,8.597494,7.2192397,5.840986,4.466636,3.0883822,4.263607,5.4427366,6.621866,7.7970915,8.976221,10.139732,11.303245,12.470661,13.634172,14.801589,13.856724,12.911859,11.963089,11.018223,10.073358,9.464272,8.855185,8.246098,7.633106,7.0240197,6.930314,6.8366084,6.7389984,6.6452928,6.551587,6.098676,5.645766,5.192855,4.7399445,4.2870336,4.4978714,4.7087092,4.9156423,5.12648,5.337318,5.9268827,6.5164475,7.1060123,7.6955767,8.289046,7.6955767,7.1021075,6.5086384,5.919074,5.3256044,5.181142,5.036679,4.8883114,4.743849,4.5993857,4.4510183,4.298747,4.1503797,3.998108,3.8497405,3.6701381,3.4905357,3.310933,3.1313305,2.951728,3.310933,3.6740425,4.037152,4.4002614,4.7633705,4.263607,3.7638438,3.2640803,2.7643168,2.260649,2.4246337,2.5886188,2.7486992,2.912684,3.076669,2.9165885,2.7565079,2.5964274,2.436347,2.2762666,2.1161861,1.9561055,1.796025,1.6359446,1.475864,1.7608855,2.0498111,2.338737,2.6237583,2.912684,3.1039999,3.2914112,3.4827268,3.6740425,3.8614538,3.7482262,3.631094,3.5178664,3.4007344,3.2875066,2.9478238,2.6081407,2.2684577,1.9287747,1.5890918,1.6008049,1.6164225,1.6320401,1.6476578,1.6632754,0.57394713,0.5622339,0.5505207,0.5388075,0.5231899,0.5114767,0.4958591,0.47633708,0.46071947,0.44119745,0.42557985,0.42557985,0.42557985,0.42557985,0.42557985,0.42557985,0.42167544,0.42167544,0.41777104,0.41386664,0.41386664,0.40605783,0.40215343,0.39824903,0.39434463,0.38653582,0.43729305,0.48805028,0.5388075,0.58566034,0.63641757,0.62860876,0.62079996,0.61689556,0.60908675,0.60127795,0.61689556,0.63641757,0.6520352,0.6715572,0.6871748,0.6637484,0.6442264,0.62079996,0.59737355,0.57394713,0.6832704,0.79649806,0.9058213,1.0151446,1.1244678,1.4055848,1.6906061,1.9717231,2.2567444,2.5378613,2.6159496,2.697942,2.77603,2.8580225,2.9361105,2.5730011,2.2059872,1.8428779,1.475864,1.1127546,1.097137,1.0815194,1.0659018,1.0541886,1.038571,0.8316377,0.62079996,0.41386664,0.20693332,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6559396,1.3157835,1.9717231,2.631567,3.2875066,3.06886,2.854118,2.6354716,2.416825,2.1981785,1.8545911,1.5110037,1.1635119,0.8199245,0.47633708,0.37872702,0.28502136,0.19131571,0.093705654,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.5388075,0.78088045,1.0190489,1.261122,1.4992905,1.5149081,1.5305257,1.5461433,1.5617609,1.5734742,1.7530766,1.9287747,2.1083772,2.2840753,2.463678,2.4792955,2.4910088,2.5066261,2.522244,2.5378613,2.9087796,3.2836022,3.6545205,4.029343,4.4002614,4.251894,4.0996222,3.951255,3.7989833,3.6506162,3.9161155,4.185519,4.4510183,4.7204223,4.985922,4.9937305,5.001539,5.009348,5.017157,5.024966,4.564246,4.0996222,3.638903,3.174279,2.7135596,3.0337205,3.3538816,3.6740425,3.9942036,4.3143644,3.8653584,3.416352,2.97125,2.522244,2.0732377,2.0810463,2.084951,2.0888553,2.096664,2.1005683,2.6862288,3.2718892,3.853645,4.4393053,5.024966,4.5447245,4.0644827,3.5842414,3.1039999,2.6237583,2.7057507,2.7838387,2.8658314,2.9439192,3.0259118,3.6818514,4.3416953,4.997635,5.6535745,6.3134184,5.989353,5.661383,5.337318,5.0132523,4.689187,4.5876727,4.4861584,4.388548,4.2870336,4.1894236,4.271416,4.3534083,4.435401,4.5173936,4.5993857,5.0327744,5.466163,5.8956475,6.329036,6.7624245,6.996689,7.2270484,7.461313,7.6916723,7.9259367,7.9610763,8.00012,8.039165,8.074304,8.113348,8.32809,8.546737,8.765383,8.98403,9.198771,9.651682,10.104593,10.557504,11.010414,11.4633255,10.534078,9.608734,8.679486,7.7541428,6.824895,7.2426662,7.660437,8.078208,8.495979,8.913751,8.203149,7.492548,6.7819467,6.0713453,5.3607445,4.657952,3.951255,3.2484627,2.541766,1.8389735,1.7491722,1.6593709,1.5656652,1.475864,1.3860629,1.4016805,1.4172981,1.4329157,1.4485333,1.4641509,2.8580225,4.251894,5.645766,7.043542,8.437413,12.220779,16.004145,19.783606,23.566973,27.350338,27.951616,28.548988,29.150267,29.751545,30.348919,35.186474,40.020123,44.853775,49.691326,54.52498,46.485813,38.450554,30.411388,22.37613,14.336966,11.471134,8.601398,5.735567,2.8658314,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3357786,0.6715572,1.0034313,1.33921,1.6749885,1.5266213,1.3743496,1.2259823,1.0737107,0.92534333,1.8194515,2.7135596,3.611572,4.50568,5.3997884,5.735567,6.0713453,6.4032197,6.7389984,7.0747766,7.7307167,8.386656,9.0386915,9.694631,10.350571,11.873287,13.399908,14.92653,16.449247,17.975868,16.761599,15.551234,14.336966,13.1266,11.912332,11.8654785,11.818625,11.771772,11.721016,11.674163,10.865952,10.061645,9.253433,8.445222,7.6370106,7.2426662,6.8483214,6.453977,6.055728,5.661383,5.001539,4.3416953,3.6818514,3.0220075,2.3621633,2.4480603,2.533957,2.6159496,2.7018464,2.787743,2.8892577,2.9868677,3.0883822,3.1859922,3.2875066,3.5608149,3.8380275,4.1113358,4.388548,4.661856,4.0761957,3.4866312,2.900971,2.3114061,1.7257458,1.5461433,1.3704453,1.1908426,1.0151446,0.8394465,1.5305257,2.2216048,2.9165885,3.6076677,4.298747,3.998108,3.6935644,3.3929255,3.0883822,2.787743,2.4714866,2.1513257,1.8350691,1.5188124,1.1986516,1.6437533,2.0888553,2.533957,2.979059,3.4241607,3.049338,2.6745155,2.2996929,1.9248703,1.5500476,1.4680552,1.3899672,1.3118792,1.2298868,1.1517987,1.5227169,1.893635,2.2684577,2.639376,3.0141985,2.5456703,2.077142,1.6086137,1.1439898,0.6754616,1.2064602,1.7335546,2.2645533,2.795552,3.3265507,2.9634414,2.6042364,2.2450314,1.8858263,1.5266213,1.4680552,1.4133936,1.358732,1.3040704,1.2494087,1.5461433,1.8467822,2.1435168,2.4402514,2.736986,2.9322062,3.1274261,3.3226464,3.5178664,3.7130866,3.5100577,3.3070288,3.1039999,2.900971,2.7018464,2.2177005,1.7335546,1.2533131,0.76916724,0.28892577,0.40605783,0.5231899,0.64032197,0.75745404,0.8745861,1.0268579,1.175225,1.3235924,1.475864,1.6242313,2.8385005,4.0488653,5.263134,6.473499,7.687768,6.1494336,4.6110992,3.076669,1.5383345,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.046852827,0.05075723,0.058566034,0.06637484,0.07418364,0.078088045,0.08589685,0.08980125,0.093705654,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.24597734,0.28892577,0.3357786,0.37872702,0.42557985,0.6949836,0.96438736,1.2337911,1.5031948,1.7765031,2.6354716,3.49444,4.3534083,5.2162814,6.0752497,5.2436123,4.40807,3.5764325,2.7447948,1.9131571,1.5617609,1.2064602,0.8550641,0.5036679,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.94486535,1.8897307,2.8345962,3.7794614,4.7243266,5.1460023,5.563773,5.985449,6.4032197,6.824895,7.7619514,8.699008,9.636065,10.573121,11.514082,11.615597,11.717112,11.818625,11.924045,12.025558,10.4286585,8.831758,7.230953,5.6340523,4.037152,5.0210614,6.008875,6.9927845,7.9766936,8.960603,10.2100115,11.455516,12.704925,13.954333,15.199838,14.106606,13.013372,11.924045,10.8308115,9.737579,8.898132,8.058686,7.2192397,6.375889,5.5364423,5.407597,5.278752,5.1460023,5.017157,4.8883114,4.575959,4.267512,3.959064,3.6467118,3.338264,3.541293,3.7443218,3.9434462,4.1464753,4.349504,4.9468775,5.5442514,6.141625,6.7389984,7.336372,6.629675,5.9229784,5.2162814,4.50568,3.7989833,3.8965936,3.9902992,4.084005,4.181615,4.2753205,4.298747,4.3260775,4.349504,4.376835,4.4002614,4.2557983,4.1113358,3.9668727,3.8185053,3.6740425,3.8887846,4.0996222,4.3143644,4.5252023,4.73604,4.3612175,3.9863946,3.611572,3.2367494,2.8619268,2.900971,2.9361105,2.9751544,3.0141985,3.049338,2.8619268,2.6706111,2.4792955,2.2918842,2.1005683,2.0107672,1.9209659,1.8311646,1.7413634,1.6515622,1.901444,2.1513257,2.4012074,2.6510892,2.900971,3.1118085,3.3187418,3.5295796,3.7404175,3.951255,3.7130866,3.4788225,3.2445583,3.0102942,2.77603,2.5261483,2.280171,2.0341935,1.7843118,1.5383345,1.6086137,1.6827974,1.7530766,1.8272603,1.901444,0.60127795,0.58566034,0.57394713,0.5622339,0.5505207,0.5388075,0.5231899,0.5075723,0.49195468,0.47633708,0.46071947,0.46071947,0.46071947,0.46071947,0.46071947,0.46071947,0.45681506,0.44900626,0.44119745,0.43338865,0.42557985,0.42167544,0.42167544,0.41777104,0.41386664,0.41386664,0.47633708,0.5388075,0.60127795,0.6637484,0.7262188,0.7145056,0.7066968,0.6949836,0.6832704,0.6754616,0.6910792,0.7066968,0.71841,0.7340276,0.74964523,0.7340276,0.7145056,0.698888,0.679366,0.6637484,0.75354964,0.8472553,0.94096094,1.0307622,1.1244678,1.4485333,1.7686942,2.0927596,2.416825,2.736986,2.8658314,2.9907722,3.1196175,3.2484627,3.3734035,2.9439192,2.5105307,2.077142,1.6437533,1.2142692,1.1674163,1.1205635,1.077615,1.0307622,0.9878138,0.78868926,0.59346914,0.39434463,0.19912452,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5231899,1.0463798,1.5656652,2.0888553,2.612045,2.3114061,2.0068626,1.7062237,1.4016805,1.1010414,0.92924774,0.75354964,0.58175594,0.40996224,0.23816854,0.19131571,0.14055848,0.093705654,0.046852827,0.0,0.042948425,0.08589685,0.12884527,0.1717937,0.21083772,0.5700427,0.92924774,1.2845483,1.6437533,1.999054,1.893635,1.7882162,1.6867018,1.5812829,1.475864,1.6437533,1.815547,1.9834363,2.15523,2.3231194,2.3075018,2.2918842,2.2723622,2.2567444,2.2372224,2.67842,3.1235218,3.5647192,4.0059166,4.4510183,4.224563,3.998108,3.775557,3.5491016,3.3265507,3.6037633,3.8809757,4.1581883,4.435401,4.7126136,4.759466,4.806319,4.853172,4.903929,4.950782,4.575959,4.2011366,3.8263142,3.4514916,3.076669,3.4983444,3.9200199,4.3416953,4.7633705,5.1889505,4.533011,3.8770714,3.2211318,2.5690966,1.9131571,1.8663043,1.8194515,1.7686942,1.7218413,1.6749885,2.15523,2.6354716,3.1157131,3.5959544,4.0761957,3.7716527,3.4710135,3.1664703,2.8658314,2.5612879,2.5651922,2.5690966,2.5690966,2.5730011,2.5769055,3.1118085,3.6467118,4.181615,4.716518,5.251421,5.0483923,4.8492675,4.650143,4.4510183,4.251894,4.2011366,4.1503797,4.0996222,4.0488653,3.998108,3.9863946,3.970777,3.9551594,3.9395418,3.9239242,4.4978714,5.0718184,5.6418614,6.2158084,6.785851,7.0474463,7.309041,7.5667315,7.8283267,8.086017,8.062591,8.039165,8.011833,7.988407,7.9610763,8.140678,8.316377,8.495979,8.671678,8.85128,9.183154,9.515028,9.846903,10.178777,10.510651,9.655587,8.796618,7.941554,7.082586,6.223617,6.676528,7.1294384,7.5823493,8.03526,8.488171,7.8947015,7.3012323,6.7116675,6.1181984,5.5247293,4.8102236,4.095718,3.3812122,2.6667068,1.9482968,1.8194515,1.6867018,1.5539521,1.4212024,1.2884527,1.319688,1.3509232,1.3860629,1.4172981,1.4485333,2.135708,2.8189783,3.506153,4.1894236,4.8765984,8.023546,11.170495,14.317443,17.464392,20.61134,23.086731,25.562122,28.037512,30.512903,32.988297,39.578926,46.173462,52.76409,59.358627,65.94926,54.763145,43.577034,32.387016,21.200905,10.010887,8.011833,6.008875,4.0059166,2.0029583,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.30454338,0.60908675,0.9136301,1.2181735,1.5266213,1.4016805,1.2767396,1.1517987,1.0268579,0.9019169,1.9482968,2.9946766,4.041056,5.0913405,6.13772,6.629675,7.1216297,7.6135845,8.109444,8.601398,9.151918,9.706344,10.256865,10.81129,11.361811,13.700547,16.039284,18.374117,20.712854,23.05159,21.474213,19.900738,18.32336,16.749886,15.176412,14.856251,14.539994,14.223738,13.903577,13.58732,12.501896,11.416472,10.331048,9.245625,8.164105,7.676055,7.191909,6.707763,6.223617,5.735567,4.9468775,4.154284,3.3616903,2.5690966,1.7765031,2.018576,2.260649,2.5027218,2.7447948,2.9868677,3.1391394,3.2875066,3.435874,3.5881457,3.736513,4.21285,4.689187,5.1616197,5.6379566,6.114294,5.263134,4.4119744,3.5608149,2.7135596,1.8623998,1.6906061,1.5227169,1.3509232,1.183034,1.0112402,1.8038338,2.592523,3.3812122,4.173806,4.9624953,4.591577,4.220659,3.853645,3.4827268,3.1118085,2.6862288,2.2567444,1.8311646,1.4016805,0.97610056,1.4602464,1.9443923,2.4285383,2.9165885,3.4007344,2.9634414,2.5261483,2.0888553,1.6515622,1.2142692,1.1869383,1.1557031,1.1283722,1.1010414,1.0737107,1.5188124,1.9600099,2.4012074,2.8463092,3.2875066,2.7213683,2.1591344,1.5929961,1.0268579,0.46071947,1.1283722,1.7921207,2.455869,3.1235218,3.78727,3.39683,3.0024853,2.6081407,2.2177005,1.8233559,1.7491722,1.6710842,1.5929961,1.5149081,1.43682,1.7530766,2.0732377,2.3894942,2.7057507,3.0259118,3.049338,3.06886,3.0922866,3.1157131,3.1391394,3.0922866,3.049338,3.0024853,2.9556324,2.912684,2.366068,1.8194515,1.2689307,0.7223144,0.1756981,0.25378615,0.3318742,0.40605783,0.48414588,0.5622339,0.80040246,1.038571,1.2767396,1.5110037,1.7491722,3.4514916,5.1499066,6.8483214,8.550641,10.249056,8.1992445,6.1494336,4.0996222,2.0498111,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.058566034,0.07027924,0.078088045,0.08980125,0.10151446,0.10151446,0.10541886,0.10932326,0.10932326,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.1835069,0.26940376,0.3553006,0.44119745,0.5231899,0.6832704,0.8433509,1.0034313,1.1635119,1.3235924,2.67842,4.0332475,5.3919797,6.746807,8.101635,6.98888,5.8800297,4.7711797,3.6584249,2.5495746,2.0810463,1.6086137,1.1400855,0.6715572,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.659844,1.319688,1.979532,2.639376,3.2992198,3.9239242,4.5447245,5.169429,5.7902284,6.4110284,7.914223,9.413514,10.912805,12.412095,13.911386,13.946525,13.97776,14.008995,14.044135,14.07537,12.2559185,10.4403715,8.62092,6.805373,4.985922,5.7785153,6.571109,7.363703,8.156297,8.94889,10.280292,11.611692,12.939189,14.27059,15.598087,14.360392,13.118792,11.881096,10.639496,9.4018,8.32809,7.2582836,6.1884775,5.1186714,4.0488653,3.8848803,3.7208953,3.5569105,3.3890212,3.2250361,3.057147,2.8892577,2.7213683,2.5534792,2.3855898,2.5808098,2.77603,2.97125,3.1664703,3.3616903,3.9668727,4.572055,5.1772375,5.7824197,6.387602,5.563773,4.743849,3.9200199,3.096191,2.2762666,2.6081407,2.9439192,3.279698,3.6154766,3.951255,4.1503797,4.349504,4.548629,4.7516575,4.950782,4.841459,4.728231,4.618908,4.5095844,4.4002614,4.462732,4.5252023,4.5876727,4.650143,4.7126136,4.462732,4.21285,3.9629683,3.7130866,3.4632049,3.3734035,3.2875066,3.2016098,3.1118085,3.0259118,2.803361,2.5847144,2.366068,2.1435168,1.9248703,1.9053483,1.8858263,1.8663043,1.8467822,1.8233559,2.0380979,2.2489357,2.463678,2.6745155,2.8892577,3.1157131,3.3460727,3.5764325,3.8067923,4.037152,3.6818514,3.3265507,2.97125,2.6159496,2.260649,2.1083772,1.9522011,1.796025,1.6437533,1.4875772,1.6164225,1.7491722,1.8780174,2.0068626,2.135708,0.62470436,0.61299115,0.60127795,0.58566034,0.57394713,0.5622339,0.5505207,0.5388075,0.5231899,0.5114767,0.4997635,0.4997635,0.4997635,0.4997635,0.4997635,0.4997635,0.48805028,0.47633708,0.46071947,0.44900626,0.43729305,0.43729305,0.43729305,0.43729305,0.43729305,0.43729305,0.5114767,0.58566034,0.6637484,0.737932,0.81211567,0.80040246,0.78868926,0.77307165,0.76135844,0.74964523,0.76135844,0.77307165,0.78868926,0.80040246,0.81211567,0.80040246,0.78868926,0.77307165,0.76135844,0.74964523,0.8238289,0.9019169,0.97610056,1.0502841,1.1244678,1.4875772,1.8506867,2.2137961,2.5769055,2.9361105,3.1118085,3.2875066,3.4632049,3.638903,3.8106966,3.310933,2.8111696,2.3114061,1.8116426,1.3118792,1.2376955,1.1635119,1.0893283,1.0112402,0.93705654,0.74964523,0.5622339,0.37482262,0.18741131,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.38653582,0.77307165,1.1635119,1.5500476,1.9365835,1.5500476,1.1635119,0.77307165,0.38653582,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.60127795,1.0737107,1.5500476,2.0263848,2.4988174,2.2762666,2.0498111,1.8233559,1.6008049,1.3743496,1.5383345,1.698415,1.8623998,2.0263848,2.1864653,2.135708,2.0888553,2.0380979,1.9873407,1.9365835,2.4480603,2.9634414,3.474918,3.9863946,4.5017757,4.2011366,3.900498,3.5998588,3.2992198,2.998581,3.2875066,3.5764325,3.8614538,4.1503797,4.4393053,4.5252023,4.6110992,4.7009,4.786797,4.8765984,4.5876727,4.298747,4.0137253,3.7247996,3.435874,3.9629683,4.4861584,5.0132523,5.5364423,6.0635366,5.2006636,4.337791,3.474918,2.612045,1.7491722,1.6515622,1.5500476,1.4485333,1.3509232,1.2494087,1.6242313,1.999054,2.3738766,2.7486992,3.1235218,2.998581,2.87364,2.7486992,2.6237583,2.4988174,2.4246337,2.35045,2.2762666,2.1981785,2.1239948,2.5378613,2.951728,3.3616903,3.775557,4.1894236,4.1113358,4.037152,3.9629683,3.8887846,3.8106966,3.8106966,3.8106966,3.8106966,3.8106966,3.8106966,3.7013733,3.5881457,3.474918,3.3616903,3.2484627,3.9629683,4.6735697,5.388075,6.098676,6.813182,7.098203,7.387129,7.676055,7.9610763,8.250002,8.164105,8.074304,7.988407,7.898606,7.812709,7.9493628,8.086017,8.226576,8.36323,8.499884,8.710721,8.925464,9.136301,9.351044,9.561881,8.773191,7.988407,7.1997175,6.4110284,5.6262436,6.114294,6.5984397,7.08649,7.57454,8.062591,7.5862536,7.113821,6.6374836,6.1611466,5.688714,4.9624953,4.2362766,3.513962,2.787743,2.0615244,1.8858263,1.7140326,1.5383345,1.3626363,1.1869383,1.2376955,1.2884527,1.33921,1.3860629,1.43682,1.4133936,1.3860629,1.3626363,1.33921,1.3118792,3.8263142,6.336845,8.85128,11.361811,13.8762455,18.22575,22.575254,26.924759,31.274261,35.623768,43.97528,52.322895,60.67441,69.025925,77.37354,63.036575,48.699608,34.362644,20.025679,5.688714,4.548629,3.4124475,2.2762666,1.1361811,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.27330816,0.5505207,0.8238289,1.1010414,1.3743496,1.2767396,1.175225,1.0737107,0.97610056,0.8745861,2.0732377,3.2757936,4.474445,5.6730967,6.8756523,7.523783,8.175818,8.823949,9.475985,10.124115,10.573121,11.0260315,11.475039,11.924045,12.373051,15.523903,18.674755,21.82561,24.976461,28.12341,26.186827,24.250242,22.31366,20.37317,18.436588,17.850927,17.261362,16.675701,16.086138,15.500477,14.13784,12.775204,11.412568,10.049932,8.687295,8.113348,7.5394006,6.9615493,6.387602,5.813655,4.8883114,3.9629683,3.0376248,2.1122816,1.1869383,1.5890918,1.9873407,2.3855898,2.787743,3.1859922,3.3890212,3.5881457,3.78727,3.9863946,4.1894236,4.860981,5.5364423,6.211904,6.8873653,7.562827,6.4500723,5.337318,4.224563,3.1118085,1.999054,1.8389735,1.6749885,1.5110037,1.3509232,1.1869383,2.0732377,2.9634414,3.8497405,4.73604,5.6262436,5.1889505,4.7516575,4.3143644,3.873167,3.435874,2.900971,2.3621633,1.8233559,1.2884527,0.74964523,1.2767396,1.7999294,2.3231194,2.8502135,3.3734035,2.87364,2.3738766,1.8741131,1.3743496,0.8745861,0.9019169,0.92534333,0.94876975,0.97610056,0.999527,1.5110037,2.0263848,2.5378613,3.049338,3.5608149,2.900971,2.2372224,1.5734742,0.9136301,0.24988174,1.0502841,1.8506867,2.6510892,3.4514916,4.251894,3.8263142,3.4007344,2.9751544,2.5495746,2.1239948,2.0263848,1.9248703,1.8233559,1.7257458,1.6242313,1.9639144,2.2996929,2.639376,2.9751544,3.310933,3.1625657,3.0141985,2.8619268,2.7135596,2.5612879,2.6745155,2.787743,2.900971,3.0141985,3.1235218,2.5105307,1.901444,1.2884527,0.6754616,0.062470436,0.10151446,0.13665408,0.1756981,0.21083772,0.24988174,0.57394713,0.9019169,1.2259823,1.5500476,1.8741131,4.0644827,6.250948,8.437413,10.6238785,12.814248,10.249056,7.687768,5.12648,2.5612879,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,0.6754616,0.7262188,0.77307165,0.8238289,0.8745861,2.7252727,4.575959,6.426646,8.273428,10.124115,8.738052,7.3519893,5.9620223,4.575959,3.1859922,2.6003318,2.0107672,1.4251068,0.8355421,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.37482262,0.74964523,1.1244678,1.4992905,1.8741131,2.7018464,3.5256753,4.349504,5.173333,6.001066,8.062591,10.124115,12.185639,14.251068,16.312593,16.273548,16.238409,16.199366,16.164225,16.125181,14.087084,12.0489855,10.010887,7.9766936,5.938596,6.5359693,7.137247,7.7385254,8.335898,8.937177,10.350571,11.763964,13.173453,14.586847,16.00024,14.614178,13.224211,11.838148,10.44818,9.062118,7.7619514,6.461786,5.1616197,3.8614538,2.5612879,2.3621633,2.1630387,1.9639144,1.7608855,1.5617609,1.5383345,1.5110037,1.4875772,1.4641509,1.43682,1.6242313,1.8116426,1.999054,2.1864653,2.3738766,2.9868677,3.5998588,4.21285,4.825841,5.4388323,4.5017757,3.5608149,2.6237583,1.6867018,0.74964523,1.3235924,1.901444,2.475391,3.049338,3.6232853,3.998108,4.376835,4.7516575,5.12648,5.5013027,5.423215,5.349031,5.2748475,5.2006636,5.12648,5.036679,4.950782,4.860981,4.775084,4.689187,4.564246,4.4393053,4.3143644,4.1894236,4.0605783,3.8497405,3.638903,3.4241607,3.213323,2.998581,2.7486992,2.4988174,2.2489357,1.999054,1.7491722,1.7999294,1.8506867,1.901444,1.9482968,1.999054,2.174752,2.35045,2.5261483,2.7018464,2.87364,3.1235218,3.3734035,3.6232853,3.873167,4.123049,3.6506162,3.174279,2.7018464,2.2255092,1.7491722,1.6867018,1.6242313,1.5617609,1.4992905,1.43682,1.6242313,1.8116426,1.999054,2.1864653,2.3738766,0.62470436,0.61299115,0.60127795,0.58566034,0.57394713,0.5622339,0.5544251,0.5427119,0.5309987,0.5231899,0.5114767,0.5114767,0.5114767,0.5114767,0.5114767,0.5114767,0.5036679,0.4958591,0.48805028,0.48414588,0.47633708,0.46852827,0.46462387,0.46071947,0.45681506,0.44900626,0.5309987,0.61689556,0.698888,0.78088045,0.8628729,0.8511597,0.8433509,0.8316377,0.8238289,0.81211567,0.8316377,0.8511597,0.8706817,0.8941081,0.9136301,0.92143893,0.92924774,0.93315214,0.94096094,0.94876975,1.0073358,1.0659018,1.1205635,1.1791295,1.2376955,1.7491722,2.260649,2.77603,3.2875066,3.7989833,3.8185053,3.8419318,3.8614538,3.8809757,3.900498,3.4905357,3.0805733,2.6706111,2.260649,1.8506867,1.6320401,1.4133936,1.1986516,0.98000497,0.76135844,0.60908675,0.45681506,0.30454338,0.15227169,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5075723,1.0151446,1.5227169,2.0302892,2.5378613,2.0302892,1.5227169,1.0151446,0.5075723,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.26159495,0.26940376,0.28111696,0.28892577,0.30063897,0.659844,1.0190489,1.3782539,1.7413634,2.1005683,1.9443923,1.7843118,1.6281357,1.4680552,1.3118792,1.4094892,1.5070993,1.6047094,1.7023194,1.7999294,1.7725986,1.7452679,1.717937,1.6906061,1.6632754,2.096664,2.533957,2.9673457,3.4007344,3.8380275,3.6857557,3.533484,3.3812122,3.2289407,3.076669,3.3148375,3.5569105,3.795079,4.0332475,4.2753205,4.388548,4.5017757,4.6110992,4.7243266,4.8375545,4.579864,4.322173,4.0644827,3.8067923,3.5491016,3.9161155,4.283129,4.6540475,5.0210614,5.388075,4.716518,4.041056,3.3694992,2.697942,2.0263848,2.0927596,2.1591344,2.2294137,2.2957885,2.3621633,2.5573835,2.7526035,2.9478238,3.1430438,3.338264,3.1391394,2.9439192,2.7447948,2.5456703,2.35045,2.2957885,2.241127,2.1864653,2.1318035,2.0732377,2.377781,2.67842,2.9829633,3.2836022,3.5881457,3.6037633,3.619381,3.631094,3.6467118,3.6623292,3.7013733,3.7443218,3.7833657,3.8224099,3.8614538,3.8263142,3.7911747,3.7560349,3.7208953,3.6857557,4.482254,5.278752,6.0713453,6.8678436,7.6643414,7.871275,8.078208,8.285142,8.492075,8.699008,8.453031,8.203149,7.957172,7.7111945,7.461313,7.601871,7.7424297,7.882988,8.023546,8.164105,8.382751,8.601398,8.823949,9.042596,9.261242,8.648251,8.031356,7.4183645,6.801469,6.1884775,6.6140575,7.0357327,7.461313,7.8868923,8.312472,7.758047,7.2036223,6.649197,6.0908675,5.5364423,4.9742084,4.4119744,3.8497405,3.2875066,2.7252727,2.6588979,2.5964274,2.5300527,2.463678,2.4012074,2.330928,2.2645533,2.1981785,2.1318035,2.0615244,2.0341935,2.0068626,1.979532,1.9522011,1.9248703,4.165997,6.4110284,8.652155,10.893282,13.138313,18.093,23.05159,28.010181,32.968773,37.92346,45.158318,52.393173,59.631935,66.86679,74.101654,62.353306,50.604958,38.856613,27.108265,15.363823,12.412095,9.464272,6.5125427,3.5608149,0.61299115,0.49195468,0.3670138,0.24597734,0.12103647,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.38653582,0.6871748,0.9878138,1.2884527,1.5890918,1.456342,1.3235924,1.1908426,1.0580931,0.92534333,2.7799344,4.6345253,6.4891167,8.343708,10.198298,11.303245,12.408191,13.513136,14.621986,15.726933,16.42582,17.124708,17.823597,18.526388,19.225277,20.775324,22.325373,23.87542,25.425468,26.975515,25.097498,23.21948,21.341463,19.463446,17.589333,17.175465,16.761599,16.351637,15.93777,15.523903,14.3682,13.216402,12.0606985,10.904996,9.749292,9.140205,8.531119,7.918128,7.309041,6.699954,5.7394714,4.7789884,3.8185053,2.8619268,1.901444,2.4597735,3.018103,3.5803368,4.138666,4.7009,4.7633705,4.825841,4.8883114,4.950782,5.0132523,5.493494,5.9776397,6.461786,6.942027,7.426173,6.3329406,5.239708,4.1464753,3.0532427,1.9639144,1.9482968,1.9326792,1.9170616,1.901444,1.8858263,2.6667068,3.4436827,4.220659,4.997635,5.774611,5.2592297,4.743849,4.2284675,3.7130866,3.2016098,2.690133,2.1786566,1.6710842,1.1596074,0.6481308,1.0893283,1.5266213,1.9639144,2.4012074,2.8385005,2.4090161,1.9834363,1.5539521,1.1283722,0.698888,0.71841,0.7418364,0.76135844,0.78088045,0.80040246,1.4485333,2.096664,2.7408905,3.3890212,4.037152,3.310933,2.5886188,1.8623998,1.1361811,0.41386664,1.0698062,1.7257458,2.3855898,3.0415294,3.7013733,3.3070288,2.9165885,2.522244,2.1318035,1.737459,1.6632754,1.5890918,1.5110037,1.43682,1.3626363,1.6242313,1.8819219,2.1435168,2.4012074,2.6628022,2.6042364,2.5456703,2.4910088,2.4324427,2.3738766,2.494913,2.6159496,2.7330816,2.854118,2.9751544,2.397303,1.8194515,1.2415999,0.6637484,0.08589685,0.14055848,0.19131571,0.24597734,0.29673457,0.3513962,0.6637484,0.98000497,1.2962615,1.6086137,1.9248703,3.7443218,5.559869,7.37932,9.194867,11.014318,8.81614,6.617962,4.4197836,2.2216048,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.031235218,0.039044023,0.046852827,0.05466163,0.062470436,0.078088045,0.093705654,0.10932326,0.12103647,0.13665408,0.14055848,0.14055848,0.14446288,0.14836729,0.14836729,0.19131571,0.23426414,0.27721256,0.32016098,0.3631094,0.29673457,0.22645533,0.16008049,0.093705654,0.023426414,0.05075723,0.078088045,0.10932326,0.13665408,0.1639849,0.12884527,0.09761006,0.06637484,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.5388075,0.58175594,0.62079996,0.659844,0.698888,2.1786566,3.6584249,5.138193,6.621866,8.101635,7.008402,5.9151692,4.8219366,3.7287042,2.639376,2.1513257,1.6632754,1.175225,0.6871748,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.38653582,0.74964523,1.1127546,1.475864,1.8389735,2.5027218,3.1664703,3.8341231,4.4978714,5.1616197,6.79366,8.421796,10.053836,11.681972,13.314012,13.368673,13.427239,13.4858055,13.544372,13.599033,12.306676,11.010414,9.714153,8.421796,7.125534,7.191909,7.2582836,7.328563,7.394938,7.461313,8.699008,9.932799,11.166591,12.404286,13.638077,12.728352,11.818625,10.9089,9.999174,9.089449,7.9220324,6.75852,5.591104,4.4275923,3.2640803,2.979059,2.697942,2.416825,2.1318035,1.8506867,2.1122816,2.3738766,2.639376,2.900971,3.1625657,3.2289407,3.2992198,3.3655949,3.4319696,3.4983444,3.873167,4.251894,4.6267166,5.001539,5.376362,4.521298,3.6662338,2.8111696,1.9561055,1.1010414,1.5149081,1.9287747,2.3465457,2.7604125,3.174279,3.5842414,3.9902992,4.396357,4.806319,5.212377,5.278752,5.349031,5.4154058,5.481781,5.548156,5.466163,5.380266,5.2943697,5.2084727,5.12648,4.9663997,4.8102236,4.6540475,4.493967,4.337791,4.0801005,3.8224099,3.5647192,3.3070288,3.049338,2.9439192,2.8345962,2.7291772,2.619854,2.514435,2.4988174,2.4831998,2.4675822,2.4519646,2.436347,2.4910088,2.5456703,2.6042364,2.6588979,2.7135596,2.912684,3.1118085,3.310933,3.513962,3.7130866,3.3538816,2.9907722,2.631567,2.2723622,1.9131571,1.815547,1.7218413,1.6281357,1.53443,1.43682,1.5851873,1.7335546,1.8819219,2.0263848,2.174752,0.62470436,0.61299115,0.60127795,0.58566034,0.57394713,0.5622339,0.5544251,0.5466163,0.5388075,0.5309987,0.5231899,0.5231899,0.5231899,0.5231899,0.5231899,0.5231899,0.5231899,0.5192855,0.5192855,0.5153811,0.5114767,0.5036679,0.49195468,0.48414588,0.47243267,0.46071947,0.5544251,0.6442264,0.7340276,0.8238289,0.9136301,0.9058213,0.8980125,0.8902037,0.8823949,0.8745861,0.9019169,0.92924774,0.95657855,0.98390937,1.0112402,1.038571,1.0659018,1.0932326,1.1205635,1.1517987,1.1908426,1.2298868,1.2689307,1.3118792,1.3509232,2.0107672,2.6745155,3.338264,3.998108,4.661856,4.5291066,4.3924527,4.2557983,4.123049,3.9863946,3.6662338,3.3460727,3.0259118,2.7057507,2.3855898,2.0263848,1.6671798,1.3079748,0.94876975,0.58566034,0.46852827,0.3513962,0.23426414,0.11713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.62860876,1.2533131,1.8819219,2.5105307,3.1391394,2.5105307,1.8819219,1.2533131,0.62860876,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.4958591,0.48805028,0.48414588,0.48024148,0.47633708,0.71841,0.96438736,1.2103647,1.456342,1.698415,1.6086137,1.5188124,1.4290112,1.33921,1.2494087,1.2806439,1.3157835,1.3470187,1.3782539,1.4133936,1.4055848,1.4016805,1.397776,1.3938715,1.3860629,1.7452679,2.1005683,2.4597735,2.8189783,3.174279,3.1703746,3.1664703,3.1586614,3.154757,3.1508527,3.3421683,3.533484,3.7287042,3.9200199,4.1113358,4.251894,4.388548,4.5252023,4.661856,4.7985106,4.572055,4.3455997,4.1191444,3.8887846,3.6623292,3.873167,4.084005,4.290938,4.5017757,4.7126136,4.2284675,3.7482262,3.2640803,2.7838387,2.2996929,2.533957,2.7682211,3.0063896,3.240654,3.474918,3.4905357,3.506153,3.521771,3.533484,3.5491016,3.279698,3.0102942,2.7408905,2.4714866,2.1981785,2.1669433,2.1318035,2.096664,2.0615244,2.0263848,2.2177005,2.4090161,2.6042364,2.795552,2.9868677,3.0922866,3.1977055,3.3031244,3.408543,3.513962,3.59205,3.6740425,3.7521305,3.8341231,3.912211,3.9551594,3.998108,4.041056,4.084005,4.126953,5.001539,5.8800297,6.75852,7.633106,8.511597,8.640442,8.769287,8.894228,9.023073,9.151918,8.741957,8.335898,7.9259367,7.519879,7.113821,7.2543793,7.3988423,7.5394006,7.6838636,7.824422,8.050878,8.281238,8.507692,8.734148,8.960603,8.519405,8.078208,7.633106,7.191909,6.7507114,7.113821,7.47693,7.8361354,8.1992445,8.562354,7.9259367,7.2934237,6.657006,6.0205884,5.388075,4.985922,4.5876727,4.1894236,3.78727,3.3890212,3.4319696,3.4788225,3.521771,3.5686235,3.611572,3.4280653,3.240654,3.057147,2.87364,2.6862288,2.6588979,2.6276627,2.5964274,2.5690966,2.5378613,4.5095844,6.481308,8.456935,10.4286585,12.400381,17.964155,23.527927,29.095606,34.659378,40.223152,46.345253,52.46345,58.585556,64.70375,70.82586,61.66613,52.510307,43.35058,34.194756,25.03893,20.27556,15.51219,10.748819,5.989353,1.2259823,0.98000497,0.7340276,0.48805028,0.24597734,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.4997635,0.8238289,1.1517987,1.475864,1.7999294,1.6359446,1.4680552,1.3040704,1.1400855,0.97610056,3.4866312,5.9932575,8.503788,11.014318,13.524849,15.086611,16.644466,18.206228,19.764084,21.325846,22.274614,23.223385,24.17606,25.124828,26.073599,26.026745,25.975988,25.925232,25.874474,25.823717,24.00817,22.188719,20.37317,18.553719,16.738173,16.500004,16.261835,16.023666,15.789403,15.551234,14.602465,13.653695,12.708829,11.760059,10.81129,10.167064,9.522837,8.878611,8.234385,7.5862536,6.590631,5.5989127,4.60329,3.6076677,2.612045,3.3343596,4.0527697,4.7711797,5.493494,6.211904,6.13772,6.0635366,5.989353,5.911265,5.8370814,6.126007,6.4188375,6.707763,6.996689,7.2856145,6.2158084,5.142098,4.068387,2.998581,1.9248703,2.05762,2.1903696,2.3231194,2.455869,2.5886188,3.2562714,3.9239242,4.591577,5.2592297,5.9268827,5.3334136,4.7399445,4.1464753,3.5569105,2.9634414,2.4792955,1.999054,1.5149081,1.0307622,0.5505207,0.9019169,1.2494087,1.6008049,1.9482968,2.2996929,1.9443923,1.5890918,1.2337911,0.8784905,0.5231899,0.5388075,0.5544251,0.5700427,0.58566034,0.60127795,1.3821584,2.1630387,2.9478238,3.7287042,4.513489,3.7247996,2.9361105,2.1513257,1.3626363,0.57394713,1.0893283,1.6047094,2.1200905,2.6354716,3.1508527,2.7916477,2.4285383,2.069333,1.7101282,1.3509232,1.3001659,1.2494087,1.1986516,1.1517987,1.1010414,1.2806439,1.4641509,1.6476578,1.8311646,2.0107672,2.0459068,2.0810463,2.1161861,2.1513257,2.1864653,2.3153105,2.4441557,2.5690966,2.697942,2.8267872,2.2840753,1.7413634,1.1986516,0.6559396,0.113227665,0.1796025,0.24597734,0.31625658,0.38263142,0.44900626,0.75354964,1.0580931,1.3665408,1.6710842,1.9756275,3.4241607,4.8687897,6.3173227,7.7658563,9.21439,7.37932,5.548156,3.7130866,1.8819219,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.06637484,0.078088045,0.093705654,0.10932326,0.12494087,0.14055848,0.16008049,0.1756981,0.19522011,0.21083772,0.20693332,0.19912452,0.19131571,0.1835069,0.1756981,0.26159495,0.3435874,0.42948425,0.5153811,0.60127795,0.48805028,0.37872702,0.26940376,0.16008049,0.05075723,0.093705654,0.13665408,0.1756981,0.21864653,0.26159495,0.21083772,0.15617609,0.10541886,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.40605783,0.43338865,0.46462387,0.4958591,0.5231899,1.6359446,2.7447948,3.853645,4.9663997,6.0752497,5.278752,4.478349,3.6818514,2.8853533,2.0888553,1.698415,1.3118792,0.92534333,0.5388075,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.39824903,0.74964523,1.1010414,1.4485333,1.7999294,2.3035975,2.8111696,3.3148375,3.8185053,4.3260775,5.520825,6.719476,7.918128,9.116779,10.311526,10.4637985,10.61607,10.768341,10.920613,11.076789,10.522364,9.971844,9.4174185,8.866898,8.312472,7.8478484,7.3832245,6.918601,6.453977,5.989353,7.043542,8.101635,9.159728,10.217821,11.275913,10.8425255,10.409137,9.975748,9.546264,9.112875,8.082112,7.0513506,6.0205884,4.9937305,3.9629683,3.5959544,3.232845,2.8658314,2.5027218,2.135708,2.6862288,3.2367494,3.78727,4.337791,4.8883114,4.83365,4.7828927,4.728231,4.677474,4.6267166,4.7633705,4.900025,5.036679,5.173333,5.3138914,4.5408196,3.767748,2.9946766,2.2216048,1.4485333,1.7062237,1.9600099,2.2137961,2.4714866,2.7252727,3.1664703,3.6037633,4.044961,4.4861584,4.9234514,5.134289,5.3451266,5.5559645,5.7668023,5.9737353,5.891743,5.8097506,5.727758,5.645766,5.563773,5.3724575,5.181142,4.9937305,4.802415,4.6110992,4.31046,4.0059166,3.7052777,3.4007344,3.1000953,3.135235,3.1703746,3.2055142,3.240654,3.2757936,3.193801,3.1157131,3.0337205,2.9556324,2.87364,2.8111696,2.7447948,2.67842,2.6159496,2.5495746,2.7018464,2.8502135,2.998581,3.1508527,3.2992198,3.0532427,2.8111696,2.5651922,2.3192148,2.0732377,1.9482968,1.8194515,1.6906061,1.5656652,1.43682,1.5461433,1.6515622,1.7608855,1.8663043,1.9756275,0.62470436,0.61299115,0.60127795,0.58566034,0.57394713,0.5622339,0.5583295,0.5544251,0.5466163,0.5427119,0.5388075,0.5388075,0.5388075,0.5388075,0.5388075,0.5388075,0.5388075,0.5427119,0.5466163,0.5466163,0.5505207,0.5349031,0.5192855,0.5036679,0.48805028,0.47633708,0.57394713,0.6715572,0.76916724,0.8667773,0.96438736,0.95657855,0.95267415,0.94876975,0.94096094,0.93705654,0.97219616,1.0073358,1.0424755,1.077615,1.1127546,1.1596074,1.2064602,1.2533131,1.3040704,1.3509232,1.3743496,1.3938715,1.4172981,1.4407244,1.4641509,2.2762666,3.0883822,3.900498,4.7126136,5.5247293,5.2358036,4.9468775,4.6540475,4.365122,4.0761957,3.8458362,3.6154766,3.3851168,3.154757,2.9243972,2.4207294,1.9209659,1.4172981,0.9136301,0.41386664,0.3318742,0.24597734,0.1639849,0.08199245,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.74574083,1.4953861,2.241127,2.9907722,3.736513,2.9907722,2.241127,1.4953861,0.74574083,0.0,0.0,0.0,0.0,0.0,0.0,0.14836729,0.30063897,0.44900626,0.60127795,0.74964523,0.7301232,0.7106012,0.6910792,0.6715572,0.6481308,0.78088045,0.9097257,1.038571,1.1713207,1.3001659,1.2767396,1.2533131,1.2337911,1.2103647,1.1869383,1.1557031,1.1205635,1.0893283,1.0580931,1.0268579,1.0424755,1.0580931,1.077615,1.0932326,1.1127546,1.3938715,1.6710842,1.9522011,2.233318,2.514435,2.6549935,2.795552,2.9400148,3.0805733,3.2250361,3.3694992,3.513962,3.6584249,3.8067923,3.951255,4.1113358,4.2753205,4.4393053,4.5993857,4.7633705,4.564246,4.369026,4.169902,3.970777,3.775557,3.8263142,3.8809757,3.9317331,3.9863946,4.037152,3.7443218,3.4514916,3.1586614,2.8658314,2.5769055,2.979059,3.3812122,3.7833657,4.185519,4.5876727,4.423688,4.2557983,4.0918136,3.9278288,3.7638438,3.4202564,3.076669,2.7330816,2.3933985,2.0498111,2.0341935,2.018576,2.0068626,1.9912452,1.9756275,2.05762,2.1396124,2.2216048,2.3035975,2.3855898,2.5808098,2.77603,2.97125,3.1664703,3.3616903,3.4827268,3.6037633,3.7208953,3.8419318,3.9629683,4.084005,4.2011366,4.322173,4.4432096,4.564246,5.520825,6.481308,7.4417906,8.402273,9.362757,9.40961,9.456462,9.503315,9.554072,9.600925,9.030883,8.464745,7.898606,7.328563,6.7624245,6.9068875,7.0513506,7.195813,7.3441806,7.4886436,7.7229075,7.957172,8.191436,8.4257,8.663869,8.39056,8.121157,7.8517528,7.5823493,7.3129454,7.6135845,7.914223,8.210958,8.511597,8.812236,8.097731,7.3832245,6.6687193,5.9542136,5.2358036,5.001539,4.7633705,4.5252023,4.2870336,4.0488653,4.2050414,4.3612175,4.513489,4.6696653,4.825841,4.521298,4.220659,3.9161155,3.6154766,3.310933,3.279698,3.2484627,3.213323,3.182088,3.1508527,4.853172,6.5554914,8.257811,9.96013,11.66245,17.83531,24.00817,30.18103,36.35389,42.52675,47.52829,52.533733,57.539177,62.54462,67.550064,60.98286,54.415653,47.84845,41.281246,34.71404,28.139027,21.564014,14.989,8.413987,1.8389735,1.4680552,1.1010414,0.7340276,0.3670138,0.0,0.05075723,0.10541886,0.15617609,0.21083772,0.26159495,0.61299115,0.96438736,1.3118792,1.6632754,2.0107672,1.815547,1.6164225,1.4212024,1.2220778,1.0268579,4.1894236,7.355894,10.518459,13.68493,16.8514,18.866072,20.880743,22.895414,24.910086,26.924759,28.12341,29.325966,30.524616,31.723269,32.925823,31.274261,29.626604,27.975042,26.32348,24.675823,22.91884,21.16186,19.400974,17.643993,15.8870125,15.824542,15.762072,15.699601,15.637131,15.57466,14.836729,14.0948925,13.353056,12.615124,11.873287,11.193921,10.514555,9.835189,9.155824,8.476458,7.445695,6.4149327,5.3841705,4.3534083,3.3265507,4.2050414,5.083532,5.9659266,6.844417,7.726812,7.5120697,7.3012323,7.08649,6.8756523,6.66091,6.75852,6.8561306,6.9537406,7.0513506,7.1489606,6.098676,5.044488,3.9942036,2.9400148,1.8858263,2.1669433,2.4480603,2.7291772,3.0063896,3.2875066,3.8458362,4.4041657,4.958591,5.5169206,6.0752497,5.4036927,4.73604,4.0644827,3.39683,2.7252727,2.2684577,1.815547,1.358732,0.9058213,0.44900626,0.7106012,0.97610056,1.2376955,1.4992905,1.7608855,1.4797685,1.1986516,0.9136301,0.63251317,0.3513962,0.359205,0.3709182,0.37872702,0.39044023,0.39824903,1.3157835,2.233318,3.1508527,4.068387,4.985922,4.138666,3.2875066,2.436347,1.5890918,0.737932,1.1088502,1.4836729,1.8545911,2.2294137,2.6003318,2.2723622,1.9443923,1.6164225,1.2884527,0.96438736,0.93705654,0.9136301,0.8862993,0.8628729,0.8394465,0.94096094,1.0463798,1.1517987,1.2572175,1.3626363,1.4914817,1.6164225,1.7452679,1.8741131,1.999054,2.135708,2.2684577,2.4051118,2.541766,2.6745155,2.1669433,1.6593709,1.1517987,0.6442264,0.13665408,0.21864653,0.30063897,0.38653582,0.46852827,0.5505207,0.8433509,1.1400855,1.43682,1.7296503,2.0263848,3.1039999,4.181615,5.2592297,6.336845,7.4144597,5.9464045,4.478349,3.0102942,1.542239,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.09761006,0.12103647,0.14055848,0.1639849,0.18741131,0.20693332,0.22645533,0.24597734,0.26940376,0.28892577,0.26940376,0.25378615,0.23426414,0.21864653,0.19912452,0.3279698,0.45681506,0.58175594,0.7106012,0.8394465,0.6832704,0.5309987,0.37872702,0.22645533,0.07418364,0.13274968,0.19131571,0.24597734,0.30454338,0.3631094,0.28892577,0.21864653,0.14446288,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.26940376,0.28892577,0.30844778,0.3318742,0.3513962,1.0893283,1.8311646,2.5690966,3.310933,4.0488653,3.5491016,3.0454338,2.541766,2.0380979,1.5383345,1.2494087,0.96438736,0.6754616,0.38653582,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.41386664,0.74964523,1.0893283,1.4251068,1.7608855,2.1083772,2.4519646,2.7994564,3.1430438,3.4866312,4.251894,5.017157,5.7824197,6.547683,7.3129454,7.558923,7.8088045,8.054782,8.300759,8.550641,8.741957,8.929368,9.120684,9.308095,9.499411,8.503788,7.504261,6.5086384,5.5091114,4.513489,5.3919797,6.2743745,7.152865,8.031356,8.913751,8.956698,9.0035515,9.0465,9.093353,9.136301,8.242193,7.348085,6.453977,5.5559645,4.661856,4.2167544,3.767748,3.3187418,2.87364,2.4246337,3.2640803,4.0996222,4.939069,5.774611,6.6140575,6.4383593,6.266566,6.094772,5.9229784,5.7511845,5.64967,5.548156,5.4505453,5.349031,5.251421,4.560342,3.8692627,3.1781836,2.4910088,1.7999294,1.893635,1.9912452,2.084951,2.1786566,2.2762666,2.7486992,3.2211318,3.6935644,4.165997,4.6384296,4.989826,5.3412223,5.6965227,6.0479193,6.3993154,6.321227,6.239235,6.1611466,6.0791545,6.001066,5.7785153,5.5559645,5.3334136,5.1108627,4.8883114,4.5408196,4.193328,3.8458362,3.4983444,3.1508527,3.3265507,3.506153,3.6818514,3.8614538,4.037152,3.892689,3.7482262,3.6037633,3.4593005,3.310933,3.1274261,2.9439192,2.7565079,2.5730011,2.3855898,2.4871042,2.5886188,2.6862288,2.787743,2.8892577,2.7565079,2.6276627,2.4988174,2.366068,2.2372224,2.077142,1.9170616,1.756981,1.5969005,1.43682,1.5031948,1.5734742,1.639849,1.7062237,1.7765031,0.62470436,0.61299115,0.60127795,0.58566034,0.57394713,0.5622339,0.5583295,0.5583295,0.5544251,0.5544251,0.5505207,0.5505207,0.5505207,0.5505207,0.5505207,0.5505207,0.5583295,0.5661383,0.57394713,0.58175594,0.58566034,0.5661383,0.5466163,0.5270943,0.5075723,0.48805028,0.59346914,0.698888,0.80430686,0.9058213,1.0112402,1.0112402,1.0073358,1.0034313,1.0034313,0.999527,1.0424755,1.0854238,1.1283722,1.1713207,1.2142692,1.2806439,1.3470187,1.4133936,1.4836729,1.5500476,1.5539521,1.5617609,1.5656652,1.5695697,1.5734742,2.5378613,3.4983444,4.462732,5.423215,6.387602,5.9425,5.4973984,5.0522966,4.607195,4.1620927,4.0215344,3.8809757,3.7443218,3.6037633,3.4632049,2.8189783,2.1708477,1.5266213,0.8823949,0.23816854,0.19131571,0.14055848,0.093705654,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.8667773,1.7335546,2.6042364,3.4710135,4.337791,3.4710135,2.6042364,1.7335546,0.8667773,0.0,0.0,0.0,0.0,0.0,0.0,0.19912452,0.39824903,0.60127795,0.80040246,0.999527,0.96438736,0.92924774,0.8941081,0.8589685,0.8238289,0.8394465,0.8550641,0.8706817,0.8862993,0.9019169,0.94486535,0.9917182,1.0346665,1.0815194,1.1244678,1.0268579,0.92924774,0.8316377,0.7340276,0.63641757,0.679366,0.71841,0.75745404,0.79649806,0.8394465,1.038571,1.2415999,1.4446288,1.6476578,1.8506867,2.1396124,2.4285383,2.7213683,3.0102942,3.2992198,3.39683,3.49444,3.59205,3.68966,3.78727,3.9746814,4.1620927,4.349504,4.5369153,4.7243266,4.5564375,4.388548,4.220659,4.056674,3.8887846,3.7833657,3.677947,3.5725281,3.4671092,3.3616903,3.260176,3.1586614,3.0532427,2.951728,2.8502135,3.4202564,3.9902992,4.560342,5.1303844,5.700427,5.35684,5.009348,4.6657605,4.318269,3.9746814,3.5608149,3.1469483,2.7291772,2.3153105,1.901444,1.9053483,1.9092526,1.9131571,1.9209659,1.9248703,1.8975395,1.8702087,1.8428779,1.815547,1.7882162,2.0732377,2.358259,2.6432803,2.9283018,3.213323,3.3734035,3.533484,3.6935644,3.853645,4.0137253,4.2089458,4.40807,4.60329,4.802415,5.001539,6.044015,7.08649,8.128965,9.171441,10.213917,10.178777,10.147541,10.116306,10.081166,10.049932,9.323712,8.59359,7.8673706,7.141152,6.4110284,6.559396,6.707763,6.8561306,7.000593,7.1489606,7.3910336,7.633106,7.8790836,8.121157,8.36323,8.265619,8.16801,8.070399,7.9727893,7.8751793,8.113348,8.351517,8.58578,8.823949,9.062118,8.265619,7.473026,6.676528,5.883934,5.087436,5.0132523,4.939069,4.860981,4.786797,4.7126136,4.9781127,5.2436123,5.5091114,5.7707067,6.036206,5.618435,5.196759,4.7789884,4.357313,3.9356375,3.9044023,3.8692627,3.8341231,3.7989833,3.7638438,5.196759,6.6257706,8.058686,9.491602,10.924518,17.706465,24.484507,31.266453,38.044495,44.826443,48.715225,52.60401,56.4967,60.385487,64.27427,60.295685,56.321003,52.342415,48.36383,44.38915,35.99859,27.611933,19.225277,10.838621,2.4480603,1.9600099,1.4719596,0.98000497,0.48805028,0.0,0.07027924,0.14055848,0.21083772,0.28111696,0.3513962,0.7262188,1.1010414,1.475864,1.8506867,2.2255092,1.9951496,1.7647898,1.53443,1.3040704,1.0737107,4.8961205,8.714626,12.537036,16.355541,20.174046,22.645533,25.113115,27.584602,30.05609,32.52367,33.97611,35.42464,36.87708,38.32561,39.774147,36.525684,33.273315,30.024853,26.77639,23.524023,21.82561,20.131098,18.432684,16.734268,15.035853,15.14908,15.262308,15.375536,15.488764,15.598087,15.067088,14.53609,14.001186,13.470188,12.939189,12.220779,11.506273,10.791768,10.077262,9.362757,8.296855,7.230953,6.168956,5.1030536,4.037152,5.0757227,6.1181984,7.1567693,8.1992445,9.237816,8.886419,8.538928,8.187531,7.8361354,7.4886436,7.3910336,7.297328,7.2036223,7.1060123,7.012306,5.9815445,4.9468775,3.9161155,2.8814487,1.8506867,2.2762666,2.7057507,3.1313305,3.5608149,3.9863946,4.435401,4.884407,5.3295093,5.7785153,6.223617,5.477876,4.728231,3.9824903,3.2367494,2.4871042,2.0615244,1.6320401,1.2064602,0.77697605,0.3513962,0.5231899,0.698888,0.8745861,1.0502841,1.2259823,1.0151446,0.80430686,0.59346914,0.38653582,0.1756981,0.1796025,0.1835069,0.19131571,0.19522011,0.19912452,1.2533131,2.3035975,3.357786,4.40807,5.462259,4.548629,3.638903,2.7252727,1.8116426,0.9019169,1.1283722,1.358732,1.5890918,1.8194515,2.0498111,1.7530766,1.4602464,1.1635119,0.8706817,0.57394713,0.57394713,0.57394713,0.57394713,0.57394713,0.57394713,0.60127795,0.62860876,0.6559396,0.6832704,0.7106012,0.93315214,1.1517987,1.3743496,1.5929961,1.8116426,1.9561055,2.096664,2.241127,2.3816853,2.5261483,2.0537157,1.5812829,1.1088502,0.63641757,0.1639849,0.26159495,0.359205,0.45681506,0.5544251,0.6481308,0.93315214,1.2181735,1.5031948,1.7882162,2.0732377,2.7838387,3.4905357,4.1972322,4.903929,5.610626,4.5095844,3.408543,2.3035975,1.2025559,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.12884527,0.16008049,0.19131571,0.21864653,0.24988174,0.27330816,0.29673457,0.31625658,0.339683,0.3631094,0.3357786,0.30844778,0.28111696,0.25378615,0.22645533,0.39434463,0.5661383,0.7340276,0.9058213,1.0737107,0.8784905,0.6832704,0.48805028,0.29673457,0.10151446,0.1717937,0.24597734,0.31625658,0.39044023,0.46071947,0.3709182,0.27721256,0.1835069,0.093705654,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.13665408,0.14446288,0.15617609,0.1639849,0.1756981,0.5466163,0.9136301,1.2845483,1.6554666,2.0263848,1.815547,1.6086137,1.4016805,1.1947471,0.9878138,0.80040246,0.61299115,0.42557985,0.23816854,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.42557985,0.74964523,1.0737107,1.4016805,1.7257458,1.9092526,2.096664,2.280171,2.463678,2.6510892,2.9829633,3.3148375,3.6467118,3.978586,4.3143644,4.6540475,4.997635,5.3412223,5.6809053,6.0244927,6.957645,7.890797,8.823949,9.753197,10.686349,9.155824,7.629202,6.098676,4.5681505,3.0376248,3.7404175,4.4432096,5.1460023,5.8487945,6.551587,7.0708723,7.5940623,8.117252,8.640442,9.163632,8.402273,7.6409154,6.883461,6.1221027,5.3607445,4.83365,4.3026514,3.7716527,3.240654,2.7135596,3.8380275,4.9624953,6.086963,7.211431,8.335898,8.043069,7.7541428,7.461313,7.168483,6.8756523,6.5359693,6.2001905,5.8644123,5.5247293,5.1889505,4.579864,3.970777,3.3655949,2.7565079,2.1513257,2.084951,2.018576,1.9561055,1.8897307,1.8233559,2.330928,2.8345962,3.338264,3.8458362,4.349504,4.845363,5.3412223,5.833177,6.329036,6.824895,6.746807,6.6687193,6.590631,6.5164475,6.4383593,6.180669,5.9268827,5.6730967,5.4193106,5.1616197,4.7711797,4.376835,3.9863946,3.59205,3.2016098,3.521771,3.8419318,4.1581883,4.478349,4.7985106,4.591577,4.380739,4.169902,3.959064,3.7482262,3.4436827,3.1391394,2.8345962,2.5300527,2.2255092,2.2762666,2.3231194,2.3738766,2.4246337,2.475391,2.4597735,2.4441557,2.4285383,2.416825,2.4012074,2.2059872,2.0146716,1.8233559,1.6281357,1.43682,1.4641509,1.4914817,1.5188124,1.5461433,1.5734742,0.62470436,0.61299115,0.60127795,0.58566034,0.57394713,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.57394713,0.58566034,0.60127795,0.61299115,0.62470436,0.60127795,0.57394713,0.5505207,0.5231899,0.4997635,0.61299115,0.7262188,0.8394465,0.94876975,1.0619974,1.0619974,1.0619974,1.0619974,1.0619974,1.0619974,1.1127546,1.1635119,1.2142692,1.261122,1.3118792,1.4016805,1.4875772,1.5734742,1.6632754,1.7491722,1.737459,1.7257458,1.7140326,1.698415,1.6867018,2.7994564,3.912211,5.024966,6.13772,7.250475,6.649197,6.0518236,5.4505453,4.8492675,4.251894,4.2011366,4.1503797,4.0996222,4.0488653,3.998108,3.213323,2.4246337,1.6359446,0.8511597,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.9878138,1.9756275,2.9634414,3.951255,4.939069,3.951255,2.9634414,1.9756275,0.9878138,0.0,0.0,0.0,0.0,0.0,0.0,0.24988174,0.4997635,0.74964523,0.999527,1.2494087,1.1986516,1.1517987,1.1010414,1.0502841,0.999527,0.9019169,0.80040246,0.698888,0.60127795,0.4997635,0.61299115,0.7262188,0.8394465,0.94876975,1.0619974,0.9019169,0.737932,0.57394713,0.41386664,0.24988174,0.31235218,0.37482262,0.43729305,0.4997635,0.5622339,0.6871748,0.81211567,0.93705654,1.0619974,1.1869383,1.6242313,2.0615244,2.4988174,2.9361105,3.3734035,3.4241607,3.474918,3.5256753,3.5764325,3.6232853,3.8380275,4.0488653,4.263607,4.474445,4.689187,4.548629,4.4119744,4.2753205,4.138666,3.998108,3.736513,3.474918,3.213323,2.951728,2.6862288,2.77603,2.8619268,2.951728,3.0376248,3.1235218,3.8614538,4.5993857,5.337318,6.0752497,6.813182,6.2860875,5.7628975,5.2358036,4.7126136,4.1894236,3.7013733,3.213323,2.7252727,2.2372224,1.7491722,1.7765031,1.7999294,1.8233559,1.8506867,1.8741131,1.737459,1.6008049,1.4641509,1.3235924,1.1869383,1.5617609,1.9365835,2.3114061,2.6862288,3.0610514,3.2640803,3.4632049,3.6623292,3.8614538,4.0605783,4.337791,4.6110992,4.8883114,5.1616197,5.4388323,6.5633,7.687768,8.812236,9.936704,11.061172,10.951848,10.838621,10.725393,10.612165,10.498938,9.612638,8.726339,7.8361354,6.949836,6.0635366,6.211904,6.364176,6.5125427,6.66091,6.813182,7.0630636,7.3129454,7.562827,7.812709,8.062591,8.136774,8.210958,8.289046,8.36323,8.437413,8.6131115,8.78881,8.960603,9.136301,9.311999,8.437413,7.562827,6.688241,5.813655,4.939069,5.024966,5.1108627,5.2006636,5.2865605,5.376362,5.7511845,6.126007,6.5008297,6.8756523,7.250475,6.7116675,6.1767645,5.6379566,5.099149,4.564246,4.5252023,4.4861584,4.4510183,4.4119744,4.376835,5.5364423,6.699954,7.8634663,9.023073,10.186585,17.573715,24.960844,32.351875,39.739006,47.126137,49.898262,52.67429,55.45032,58.226353,60.998478,59.612415,58.226353,56.836384,55.45032,54.06426,43.862057,33.663757,23.461554,13.263254,3.0610514,2.4480603,1.8389735,1.2259823,0.61299115,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.8355421,1.2376955,1.6359446,2.0380979,2.436347,2.174752,1.9131571,1.6515622,1.3860629,1.1244678,5.5989127,10.073358,14.551707,19.026152,23.500597,26.424995,29.349392,32.27379,35.198185,38.126488,39.8249,41.52332,43.225636,44.924053,46.626373,41.7732,36.92393,32.074665,27.225397,22.37613,20.73628,19.100336,17.464392,15.824542,14.188598,14.473619,14.762545,15.051471,15.336493,15.625418,15.3013525,14.973383,14.649317,14.325252,14.001186,13.251541,12.501896,11.748346,10.998701,10.249056,9.148014,8.050878,6.949836,5.8487945,4.7516575,5.950309,7.1489606,8.351517,9.550168,10.748819,10.260769,9.776623,9.288573,8.800523,8.312472,8.023546,7.7385254,7.4495993,7.1606736,6.8756523,5.860508,4.8492675,3.8380275,2.8267872,1.8116426,2.3855898,2.9634414,3.5373883,4.1113358,4.689187,5.024966,5.3607445,5.700427,6.036206,6.375889,5.548156,4.7243266,3.900498,3.076669,2.2489357,1.8506867,1.4485333,1.0502841,0.6481308,0.24988174,0.3357786,0.42557985,0.5114767,0.60127795,0.6871748,0.5505207,0.41386664,0.27330816,0.13665408,0.0,0.0,0.0,0.0,0.0,0.0,1.1869383,2.3738766,3.5608149,4.7516575,5.938596,4.9624953,3.9863946,3.0141985,2.0380979,1.0619974,1.1517987,1.2376955,1.3235924,1.4133936,1.4992905,1.2376955,0.97610056,0.7106012,0.44900626,0.18741131,0.21083772,0.23816854,0.26159495,0.28892577,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.37482262,0.6871748,0.999527,1.3118792,1.6242313,1.7765031,1.9248703,2.0732377,2.2255092,2.3738766,1.9365835,1.4992905,1.0619974,0.62470436,0.18741131,0.30063897,0.41386664,0.5231899,0.63641757,0.74964523,1.0268579,1.3001659,1.5734742,1.8506867,2.1239948,2.463678,2.7994564,3.1391394,3.474918,3.8106966,3.076669,2.338737,1.6008049,0.8628729,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.1639849,0.19912452,0.23816854,0.27330816,0.31235218,0.3357786,0.3631094,0.38653582,0.41386664,0.43729305,0.39824903,0.3631094,0.3240654,0.28892577,0.24988174,0.46071947,0.6754616,0.8862993,1.1010414,1.3118792,1.0737107,0.8394465,0.60127795,0.3631094,0.12494087,0.21083772,0.30063897,0.38653582,0.47633708,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.3513962,0.26159495,0.1756981,0.08589685,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.43729305,0.74964523,1.0619974,1.3743496,1.6867018,1.7140326,1.737459,1.7608855,1.7882162,1.8116426,1.7140326,1.6125181,1.5110037,1.4133936,1.3118792,1.7491722,2.1864653,2.6237583,3.0610514,3.4983444,5.173333,6.8483214,8.52331,10.198298,11.873287,9.811763,7.7502384,5.688714,3.6232853,1.5617609,2.0888553,2.612045,3.1391394,3.6623292,4.1894236,5.1889505,6.1884775,7.1880045,8.187531,9.187058,8.562354,7.9376497,7.3129454,6.688241,6.0635366,5.4505453,4.8375545,4.224563,3.611572,2.998581,4.4119744,5.825368,7.238762,8.648251,10.061645,9.651682,9.237816,8.823949,8.413987,8.00012,7.426173,6.8483214,6.2743745,5.700427,5.12648,4.5993857,4.0761957,3.5491016,3.0259118,2.4988174,2.2762666,2.0498111,1.8233559,1.6008049,1.3743496,1.9131571,2.4519646,2.9868677,3.5256753,4.0605783,4.7009,5.337318,5.9737353,6.6140575,7.250475,7.1762915,7.098203,7.0240197,6.949836,6.8756523,6.5867267,6.3017054,6.012779,5.7238536,5.4388323,5.001539,4.564246,4.123049,3.6857557,3.2484627,3.7130866,4.173806,4.6384296,5.099149,5.563773,5.2865605,5.0132523,4.73604,4.462732,4.1894236,3.7638438,3.338264,2.912684,2.4871042,2.0615244,2.0615244,2.0615244,2.0615244,2.0615244,2.0615244,2.1630387,2.260649,2.3621633,2.463678,2.5612879,2.338737,2.1122816,1.8858263,1.6632754,1.43682,1.4251068,1.4133936,1.4016805,1.3860629,1.3743496,0.62470436,0.61299115,0.60127795,0.58566034,0.57394713,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.5583295,0.5583295,0.5544251,0.5544251,0.5505207,0.5661383,0.58175594,0.59346914,0.60908675,0.62470436,0.60127795,0.58175594,0.5583295,0.5349031,0.5114767,0.6442264,0.77697605,0.9097257,1.0424755,1.175225,1.1908426,1.2103647,1.2259823,1.2455044,1.261122,1.2415999,1.2220778,1.2025559,1.183034,1.1635119,1.2962615,1.4290112,1.5617609,1.6906061,1.8233559,1.9639144,2.1044729,2.2450314,2.3855898,2.5261483,3.638903,4.7516575,5.8644123,6.9732623,8.086017,7.519879,6.9537406,6.3836975,5.8175592,5.251421,5.12648,5.001539,4.8765984,4.7516575,4.6267166,3.7091823,2.795552,1.8819219,0.96438736,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.1717937,0.25769055,0.3435874,0.42557985,0.5114767,0.40996224,0.30844778,0.20693332,0.10151446,0.0,0.78868926,1.5812829,2.3699722,3.1586614,3.951255,3.1586614,2.3699722,1.5812829,0.78868926,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.41386664,0.8160201,1.2181735,1.6242313,2.0263848,1.7804074,1.53443,1.2884527,1.0463798,0.80040246,0.7223144,0.6442264,0.5661383,0.48805028,0.41386664,0.5036679,0.59737355,0.6910792,0.78088045,0.8745861,0.75745404,0.64032197,0.5231899,0.40605783,0.28892577,0.3435874,0.40215343,0.46071947,0.5192855,0.57394713,0.7340276,0.8902037,1.0463798,1.2064602,1.3626363,1.7140326,2.0615244,2.4129205,2.7643168,3.1118085,3.2055142,3.2992198,3.3890212,3.4827268,3.5764325,3.6662338,3.7560349,3.8458362,3.9356375,4.025439,3.9902992,3.9551594,3.9200199,3.8848803,3.8497405,3.6271896,3.4046388,3.182088,2.959537,2.736986,2.893162,3.0532427,3.2094188,3.3655949,3.5256753,4.087909,4.650143,5.212377,5.774611,6.336845,5.9737353,5.610626,5.251421,4.8883114,4.5252023,4.1074314,3.68966,3.2718892,2.854118,2.436347,2.3543546,2.2684577,2.182561,2.096664,2.0107672,1.8467822,1.6827974,1.5188124,1.3509232,1.1869383,1.5227169,1.8584955,2.194274,2.5261483,2.8619268,3.0063896,3.1508527,3.2992198,3.4436827,3.5881457,3.8302186,4.0722914,4.3143644,4.5564375,4.7985106,5.786324,6.7702336,7.7541428,8.741957,9.725866,9.768814,9.811763,9.850807,9.893755,9.936704,9.21439,8.488171,7.7619514,7.0357327,6.3134184,6.3017054,6.2860875,6.2743745,6.262661,6.250948,6.524256,6.79366,7.066968,7.3402762,7.6135845,7.6135845,7.6135845,7.6135845,7.6135845,7.6135845,7.719003,7.8283267,7.9337454,8.043069,8.148487,7.433982,6.715572,5.997162,5.278752,4.564246,4.677474,4.7907014,4.9078336,5.0210614,5.138193,5.446641,5.7511845,6.0596323,6.36808,6.676528,6.2587566,5.84489,5.4310236,5.0132523,4.5993857,4.5017757,4.4041657,4.3065557,4.2089458,4.1113358,5.044488,5.9776397,6.910792,7.843944,8.773191,16.46877,24.16044,31.852114,39.543785,47.239365,48.67618,50.113003,51.549824,52.986645,54.423462,52.775806,51.124245,49.476585,47.825024,46.173462,37.681385,29.189312,20.697237,12.205161,3.7130866,3.0141985,2.3114061,1.6125181,0.9136301,0.21083772,0.25769055,0.30063897,0.3474918,0.39434463,0.43729305,0.81211567,1.1869383,1.5617609,1.9365835,2.3114061,2.4324427,2.5534792,2.6706111,2.7916477,2.912684,7.3129454,11.713207,16.113468,20.51373,24.91399,27.826675,30.743263,33.65595,36.572536,39.489124,39.719482,39.953747,40.18411,40.418373,40.64873,36.900505,33.148376,29.400148,25.648018,21.899792,20.747993,19.6001,18.448301,17.300406,16.148607,16.531239,16.91387,17.296501,17.679134,18.061766,16.827974,15.594183,14.356487,13.122696,11.888905,11.43209,10.979179,10.522364,10.065549,9.612638,8.847376,8.082112,7.3168497,6.551587,5.786324,6.7624245,7.7385254,8.710721,9.686822,10.662923,10.170968,9.682918,9.190963,8.702912,8.210958,8.1992445,8.183627,8.16801,8.152391,8.136774,7.039637,5.9425,4.845363,3.7482262,2.6510892,3.1235218,3.5959544,4.068387,4.5408196,5.0132523,5.2006636,5.388075,5.575486,5.7628975,5.950309,5.153811,4.3612175,3.5647192,2.7682211,1.9756275,1.620327,1.2650263,0.9097257,0.5544251,0.19912452,0.26940376,0.339683,0.40996224,0.48024148,0.5505207,0.44119745,0.3318742,0.21864653,0.10932326,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.96048295,1.9092526,2.854118,3.802888,4.7516575,3.970777,3.1898966,2.4090161,1.6281357,0.8511597,0.93315214,1.0151446,1.097137,1.1791295,1.261122,1.0580931,0.8511597,0.6481308,0.44119745,0.23816854,0.25378615,0.26940376,0.28111696,0.29673457,0.31235218,0.27330816,0.23426414,0.19131571,0.15227169,0.113227665,0.37872702,0.6442264,0.9058213,1.1713207,1.43682,1.5734742,1.7140326,1.8506867,1.9873407,2.1239948,1.7530766,1.3860629,1.0151446,0.6442264,0.27330816,0.3513962,0.42557985,0.4997635,0.57394713,0.6481308,1.116659,1.5812829,2.0459068,2.5105307,2.9751544,2.9907722,3.0063896,3.018103,3.0337205,3.049338,2.475391,1.901444,1.3235924,0.74964523,0.1756981,0.31625658,0.46071947,0.60127795,0.74574083,0.8862993,1.0815194,1.2728351,1.4641509,1.6593709,1.8506867,1.5773785,1.3040704,1.0307622,0.76135844,0.48805028,0.46852827,0.44900626,0.42557985,0.40605783,0.38653582,0.5388075,0.6910792,0.8433509,0.9956226,1.1517987,0.98390937,0.8199245,0.6559396,0.48805028,0.3240654,0.39044023,0.45681506,0.5192855,0.58566034,0.6481308,0.5388075,0.42948425,0.32016098,0.21083772,0.10151446,0.3709182,0.6442264,0.91753453,1.1908426,1.4641509,1.1791295,0.8980125,0.61689556,0.3318742,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.07027924,0.14055848,0.21083772,0.28111696,0.3513962,0.28111696,0.21083772,0.14055848,0.07027924,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.1756981,0.58956474,1.0034313,1.4212024,1.8350691,2.2489357,2.366068,2.4792955,2.5964274,2.7096553,2.8267872,2.7408905,2.6588979,2.5769055,2.494913,2.4129205,2.639376,2.8619268,3.0883822,3.310933,3.5373883,4.83365,6.126007,7.422269,8.718531,10.010887,8.331994,6.6531014,4.9742084,3.2914112,1.6125181,2.0615244,2.514435,2.9634414,3.4124475,3.8614538,4.73604,5.610626,6.4891167,7.363703,8.238289,7.773665,7.309041,6.844417,6.375889,5.911265,5.376362,4.8375545,4.298747,3.7638438,3.2250361,4.423688,5.618435,6.817086,8.015738,9.21439,9.066022,8.917655,8.769287,8.62092,8.476458,7.8205175,7.168483,6.5164475,5.8644123,5.212377,4.911738,4.607195,4.3065557,4.0020123,3.7013733,3.4007344,3.1000953,2.7994564,2.4988174,2.1981785,2.7135596,3.2289407,3.7443218,4.2597027,4.775084,5.251421,5.7316628,6.2079997,6.6843367,7.1606736,6.984976,6.8092775,6.629675,6.453977,6.2743745,6.0752497,5.8761253,5.6730967,5.473972,5.2748475,4.9351645,4.5954814,4.2557983,3.9161155,3.5764325,3.9356375,4.298747,4.661856,5.024966,5.388075,5.181142,4.9781127,4.7711797,4.5681505,4.3612175,3.8653584,3.3655949,2.8697357,2.3738766,1.8741131,1.9443923,2.0107672,2.077142,2.1435168,2.2137961,2.330928,2.4480603,2.5651922,2.6823244,2.7994564,2.6237583,2.4441557,2.2684577,2.0888553,1.9131571,1.7530766,1.5929961,1.4329157,1.2728351,1.1127546,0.62470436,0.61299115,0.60127795,0.58566034,0.57394713,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.5583295,0.5544251,0.5466163,0.5427119,0.5388075,0.5544251,0.57394713,0.58956474,0.60908675,0.62470436,0.60518235,0.58566034,0.5661383,0.5466163,0.5231899,0.679366,0.8316377,0.98390937,1.1361811,1.2884527,1.3235924,1.358732,1.3938715,1.4290112,1.4641509,1.3743496,1.2806439,1.1908426,1.1010414,1.0112402,1.1908426,1.3665408,1.5461433,1.7218413,1.901444,2.194274,2.4831998,2.77603,3.06886,3.3616903,4.474445,5.5871997,6.699954,7.812709,8.925464,8.39056,7.8556576,7.320754,6.785851,6.250948,6.0518236,5.8487945,5.64967,5.4505453,5.251421,4.2089458,3.1664703,2.1239948,1.0815194,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.3435874,0.5153811,0.6832704,0.8550641,1.0268579,0.8199245,0.61689556,0.40996224,0.20693332,0.0,0.59346914,1.183034,1.7765031,2.3699722,2.9634414,2.3699722,1.7765031,1.183034,0.59346914,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.58175594,1.1361811,1.6906061,2.2450314,2.7994564,2.358259,1.9209659,1.4797685,1.038571,0.60127795,0.5466163,0.48805028,0.43338865,0.37872702,0.3240654,0.39824903,0.46852827,0.5427119,0.61689556,0.6871748,0.61689556,0.5427119,0.46852827,0.39824903,0.3240654,0.37872702,0.42948425,0.48414588,0.5349031,0.58566034,0.77697605,0.96829176,1.1557031,1.3470187,1.5383345,1.7999294,2.0615244,2.3231194,2.5886188,2.8502135,2.9868677,3.1196175,3.2562714,3.3890212,3.5256753,3.49444,3.4593005,3.4280653,3.39683,3.3616903,3.4280653,3.4983444,3.5647192,3.631094,3.7013733,3.5178664,3.3343596,3.1508527,2.97125,2.787743,3.0141985,3.240654,3.4710135,3.697469,3.9239242,4.3143644,4.7009,5.087436,5.473972,5.8644123,5.661383,5.462259,5.263134,5.0640097,4.860981,4.513489,4.165997,3.8185053,3.4710135,3.1235218,2.9283018,2.7330816,2.541766,2.3465457,2.1513257,1.9561055,1.7647898,1.5734742,1.3782539,1.1869383,1.4836729,1.7765031,2.0732377,2.366068,2.6628022,2.7526035,2.8424048,2.9322062,3.0220075,3.1118085,3.3226464,3.533484,3.7443218,3.951255,4.1620927,5.009348,5.852699,6.6960497,7.5433054,8.386656,8.58578,8.781001,8.980125,9.17925,9.37447,8.812236,8.250002,7.687768,7.125534,6.5633,6.387602,6.211904,6.036206,5.8644123,5.688714,5.9815445,6.278279,6.571109,6.8678436,7.1606736,7.08649,7.012306,6.9381227,6.8639393,6.785851,6.8287997,6.8678436,6.9068875,6.9459314,6.98888,6.426646,5.8683167,5.3060827,4.747753,4.1894236,4.3299823,4.474445,4.6150036,4.755562,4.900025,5.138193,5.380266,5.618435,5.860508,6.098676,5.805846,5.5169206,5.22409,4.93126,4.6384296,4.478349,4.322173,4.165997,4.0059166,3.8497405,4.552533,5.2553253,5.958118,6.66091,7.363703,15.359919,23.356134,31.356255,39.35247,47.348686,47.4502,47.551716,47.649326,47.75084,47.84845,45.939198,44.02604,42.112885,40.199726,38.286568,31.500717,24.718771,17.93292,11.147068,4.3612175,3.5764325,2.787743,1.999054,1.2142692,0.42557985,0.42557985,0.42948425,0.43338865,0.43338865,0.43729305,0.78868926,1.1361811,1.4875772,1.8389735,2.1864653,2.690133,3.193801,3.6935644,4.1972322,4.7009,9.023073,13.349152,17.675228,22.001307,26.32348,29.228355,32.133232,35.04201,37.946884,40.85176,39.614067,38.380276,37.146484,35.908787,34.674995,32.023907,29.376722,26.725634,24.074545,21.423454,20.76361,20.099863,19.436115,18.77627,18.112522,18.58886,19.069101,19.545437,20.021774,20.498112,18.354595,16.211079,14.063657,11.92014,9.776623,9.616543,9.456462,9.296382,9.136301,8.976221,8.546737,8.113348,7.6838636,7.2543793,6.824895,7.57454,8.324185,9.073831,9.823476,10.573121,10.081166,9.589212,9.097258,8.605303,8.113348,8.371038,8.628729,8.886419,9.14411,9.4018,8.218767,7.0357327,5.852699,4.6696653,3.4866312,3.8575494,4.2284675,4.5993857,4.9663997,5.337318,5.376362,5.4115014,5.4505453,5.4856853,5.5247293,4.759466,3.9942036,3.2289407,2.463678,1.698415,1.3899672,1.0815194,0.76916724,0.46071947,0.14836729,0.20302892,0.25378615,0.30844778,0.359205,0.41386664,0.3318742,0.24597734,0.1639849,0.08199245,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.7340276,1.4407244,2.1474214,2.854118,3.5608149,2.979059,2.3933985,1.8077383,1.2220778,0.63641757,0.7145056,0.79259366,0.8706817,0.94876975,1.0268579,0.8784905,0.7301232,0.58175594,0.43338865,0.28892577,0.29283017,0.29673457,0.30063897,0.30844778,0.31235218,0.28111696,0.25378615,0.22255093,0.19131571,0.1639849,0.37872702,0.59737355,0.8160201,1.0307622,1.2494087,1.3743496,1.4992905,1.6242313,1.7491722,1.8741131,1.5734742,1.2689307,0.96829176,0.6637484,0.3631094,0.39824903,0.43729305,0.47633708,0.5114767,0.5505207,1.2064602,1.8584955,2.514435,3.1703746,3.8263142,3.5178664,3.2094188,2.900971,2.5964274,2.2879796,1.8741131,1.4641509,1.0502841,0.63641757,0.22645533,0.5114767,0.79649806,1.0815194,1.3665408,1.6515622,1.999054,2.3465457,2.6940374,3.0415294,3.3890212,2.8189783,2.2489357,1.678893,1.1088502,0.5388075,0.5349031,0.5309987,0.5309987,0.5270943,0.5231899,0.61689556,0.7106012,0.80430686,0.8941081,0.9878138,0.8941081,0.80430686,0.7106012,0.61689556,0.5231899,0.5661383,0.60908675,0.6520352,0.6949836,0.737932,0.62860876,0.5231899,0.41386664,0.30844778,0.19912452,0.74574083,1.2884527,1.8350691,2.3816853,2.9243972,2.358259,1.796025,1.2298868,0.6637484,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10541886,0.15617609,0.21083772,0.26159495,0.21083772,0.15617609,0.10541886,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.12494087,0.14836729,0.1756981,0.19912452,0.22645533,0.7418364,1.261122,1.7765031,2.2957885,2.8111696,3.018103,3.2211318,3.4280653,3.631094,3.8380275,3.7716527,3.7091823,3.6428072,3.5764325,3.513962,3.5256753,3.5373883,3.5491016,3.5608149,3.5764325,4.4900627,5.4036927,6.321227,7.2348576,8.148487,6.852226,5.5559645,4.2557983,2.959537,1.6632754,2.0380979,2.4129205,2.787743,3.1625657,3.5373883,4.2870336,5.036679,5.786324,6.5359693,7.2856145,6.9810715,6.676528,6.3719845,6.067441,5.7628975,5.298274,4.8375545,4.376835,3.912211,3.4514916,4.4314966,5.4154058,6.3993154,7.37932,8.36323,8.480362,8.597494,8.714626,8.831758,8.94889,8.218767,7.4886436,6.75852,6.028397,5.298274,5.2201858,5.138193,5.0601053,4.9781127,4.900025,4.5252023,4.1503797,3.775557,3.4007344,3.0259118,3.5178664,4.009821,4.5017757,4.9937305,5.4856853,5.805846,6.1221027,6.4383593,6.75852,7.0747766,6.79366,6.5164475,6.2353306,5.9542136,5.6730967,5.563773,5.4505453,5.337318,5.22409,5.1108627,4.8687897,4.6267166,4.3846436,4.142571,3.900498,4.1620927,4.423688,4.689187,4.950782,5.212377,5.0757227,4.942973,4.806319,4.6735697,4.5369153,3.9668727,3.39683,2.8267872,2.2567444,1.6867018,1.8233559,1.9561055,2.0927596,2.2294137,2.3621633,2.4988174,2.631567,2.7682211,2.900971,3.0376248,2.9087796,2.77603,2.6471848,2.5183394,2.3855898,2.0810463,1.7725986,1.4641509,1.1557031,0.8511597,0.62470436,0.61299115,0.60127795,0.58566034,0.57394713,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.5544251,0.5466163,0.5388075,0.5309987,0.5231899,0.5466163,0.5661383,0.58566034,0.60518235,0.62470436,0.60908675,0.58956474,0.57394713,0.5544251,0.5388075,0.7106012,0.8823949,1.0541886,1.2259823,1.4016805,1.4524376,1.5031948,1.5578566,1.6086137,1.6632754,1.5031948,1.3431144,1.183034,1.0229534,0.8628729,1.0854238,1.3079748,1.5305257,1.7530766,1.9756275,2.4207294,2.8658314,3.310933,3.7560349,4.2011366,5.3138914,6.426646,7.5394006,8.648251,9.761005,9.261242,8.757574,8.253906,7.7541428,7.250475,6.9732623,6.699954,6.426646,6.1494336,5.8761253,4.704805,3.533484,2.366068,1.1947471,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.05075723,0.10541886,0.15617609,0.21083772,0.26159495,0.5192855,0.77307165,1.0268579,1.2806439,1.5383345,1.2298868,0.92143893,0.61689556,0.30844778,0.0,0.39434463,0.78868926,1.1869383,1.5812829,1.9756275,1.5812829,1.1869383,0.78868926,0.39434463,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.74574083,1.4524376,2.1591344,2.8658314,3.5764325,2.9400148,2.3035975,1.6710842,1.0346665,0.39824903,0.3670138,0.3357786,0.30063897,0.26940376,0.23816854,0.28892577,0.3435874,0.39434463,0.44900626,0.4997635,0.47243267,0.44510186,0.41777104,0.39044023,0.3631094,0.40996224,0.45681506,0.5036679,0.5544251,0.60127795,0.8238289,1.0463798,1.2689307,1.4914817,1.7140326,1.8858263,2.0615244,2.2372224,2.4129205,2.5886188,2.7643168,2.9439192,3.1196175,3.2992198,3.474918,3.3187418,3.1664703,3.0102942,2.854118,2.7018464,2.8697357,3.0415294,3.2094188,3.3812122,3.5491016,3.408543,3.2640803,3.1235218,2.979059,2.8385005,3.135235,3.4319696,3.7287042,4.029343,4.3260775,4.5369153,4.7516575,4.9624953,5.173333,5.388075,5.349031,5.3138914,5.2748475,5.2358036,5.2006636,4.9234514,4.646239,4.369026,4.0918136,3.8106966,3.506153,3.2016098,2.8970666,2.592523,2.2879796,2.069333,1.8467822,1.6281357,1.4055848,1.1869383,1.4407244,1.698415,1.9522011,2.2059872,2.463678,2.4988174,2.533957,2.5690966,2.6042364,2.639376,2.815074,2.9907722,3.1703746,3.3460727,3.5256753,4.2284675,4.9351645,5.6418614,6.3446536,7.0513506,7.4027467,7.7541428,8.109444,8.460839,8.812236,8.413987,8.011833,7.6135845,7.211431,6.813182,6.473499,6.13772,5.801942,5.462259,5.12648,5.4427366,5.758993,6.0791545,6.395411,6.7116675,6.5633,6.4110284,6.262661,6.114294,5.9620223,5.9346914,5.9073606,5.8800297,5.852699,5.825368,5.423215,5.0210614,4.618908,4.2167544,3.8106966,3.9824903,4.154284,4.322173,4.493967,4.661856,4.83365,5.009348,5.181142,5.3529353,5.5247293,5.35684,5.185046,5.0132523,4.845363,4.6735697,4.4588275,4.240181,4.0215344,3.8067923,3.5881457,4.0605783,4.533011,5.0054436,5.477876,5.950309,14.251068,22.555733,30.856491,39.161156,47.461914,46.224216,44.986523,43.74883,42.51113,41.273438,39.098682,36.92393,34.74918,32.57443,30.399675,25.323954,20.244326,15.168603,10.088976,5.0132523,4.138666,3.2640803,2.3855898,1.5110037,0.63641757,0.59737355,0.5583295,0.5192855,0.47633708,0.43729305,0.76135844,1.0893283,1.4133936,1.737459,2.0615244,2.9478238,3.8341231,4.716518,5.602817,6.4891167,10.737106,14.989,19.23699,23.488884,27.736874,30.63394,33.527103,36.424168,39.31733,42.214397,39.508648,36.8068,34.104954,31.403107,28.701262,27.151213,25.601166,24.051117,22.50107,20.951023,20.775324,20.599627,20.423927,20.24823,20.076437,20.646479,21.220427,21.794373,22.364416,22.938364,19.881216,16.827974,13.770826,10.717585,7.6643414,7.7970915,7.9337454,8.066495,8.203149,8.335898,8.242193,8.148487,8.050878,7.957172,7.8634663,8.386656,8.913751,9.43694,9.964035,10.487225,9.991365,9.499411,9.0035515,8.507692,8.011833,8.542832,9.073831,9.600925,10.131924,10.662923,9.393991,8.128965,6.860035,5.591104,4.3260775,4.591577,4.860981,5.12648,5.395884,5.661383,5.548156,5.4388323,5.3256044,5.212377,5.099149,4.365122,3.631094,2.893162,2.1591344,1.4251068,1.1596074,0.8941081,0.62860876,0.3631094,0.10151446,0.13665408,0.1717937,0.20693332,0.23816854,0.27330816,0.21864653,0.1639849,0.10932326,0.05466163,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.5036679,0.97219616,1.4407244,1.9092526,2.3738766,1.9834363,1.5969005,1.2064602,0.8160201,0.42557985,0.4958591,0.5700427,0.6442264,0.7145056,0.78868926,0.698888,0.60908675,0.5192855,0.42557985,0.3357786,0.3318742,0.3279698,0.3240654,0.31625658,0.31235218,0.29283017,0.27330816,0.25378615,0.23426414,0.21083772,0.38263142,0.5544251,0.7223144,0.8941081,1.0619974,1.175225,1.2884527,1.4016805,1.5110037,1.6242313,1.3899672,1.1557031,0.92143893,0.6832704,0.44900626,0.44900626,0.44900626,0.44900626,0.44900626,0.44900626,1.2962615,2.1396124,2.9868677,3.8302186,4.6735697,4.044961,3.416352,2.7838387,2.15523,1.5266213,1.2767396,1.0268579,0.77307165,0.5231899,0.27330816,0.7027924,1.1283722,1.5578566,1.9834363,2.4129205,2.9165885,3.416352,3.9200199,4.423688,4.9234514,4.056674,3.1898966,2.3231194,1.456342,0.58566034,0.60127795,0.61689556,0.63251317,0.6481308,0.6637484,0.6949836,0.7262188,0.76135844,0.79259366,0.8238289,0.80430686,0.78478485,0.76526284,0.74574083,0.7262188,0.74574083,0.76526284,0.78478485,0.80430686,0.8238289,0.71841,0.61689556,0.5114767,0.40605783,0.30063897,1.116659,1.9365835,2.7526035,3.5686235,4.388548,3.541293,2.6940374,1.8467822,0.9956226,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.1756981,0.19912452,0.22645533,0.24988174,0.27330816,0.8941081,1.5149081,2.135708,2.7565079,3.3734035,3.6701381,3.9668727,4.2597027,4.5564375,4.8492675,4.802415,4.755562,4.7087092,4.661856,4.6110992,4.4119744,4.21285,4.0137253,3.8106966,3.611572,4.1464753,4.6813784,5.2162814,5.7511845,6.2860875,5.3724575,4.4588275,3.541293,2.6276627,1.7140326,2.0107672,2.3114061,2.612045,2.912684,3.213323,3.8380275,4.462732,5.087436,5.7121406,6.336845,6.192382,6.0479193,5.903456,5.758993,5.610626,5.22409,4.8375545,4.4510183,4.0605783,3.6740425,4.4432096,5.2084727,5.9776397,6.746807,7.5120697,7.8947015,8.277332,8.659965,9.042596,9.425227,8.617016,7.8088045,7.000593,6.196286,5.388075,5.5286336,5.6730967,5.813655,5.958118,6.098676,5.64967,5.2006636,4.7516575,4.298747,3.8497405,4.318269,4.7907014,5.2592297,5.7316628,6.2001905,6.356367,6.5164475,6.6726236,6.8287997,6.98888,6.606249,6.223617,5.840986,5.4583545,5.0757227,5.0483923,5.024966,5.001539,4.9742084,4.950782,4.806319,4.661856,4.513489,4.369026,4.224563,4.388548,4.548629,4.7126136,4.8765984,5.036679,4.9742084,4.9078336,4.841459,4.7789884,4.7126136,4.068387,3.4280653,2.7838387,2.1435168,1.4992905,1.7023194,1.9053483,2.1083772,2.3114061,2.514435,2.6667068,2.8189783,2.97125,3.1235218,3.2757936,3.193801,3.1118085,3.0259118,2.9439192,2.8619268,2.4090161,1.9522011,1.4992905,1.0424755,0.58566034,0.62470436,0.61299115,0.60127795,0.58566034,0.57394713,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.5544251,0.5427119,0.5309987,0.5231899,0.5114767,0.5349031,0.5583295,0.58175594,0.60127795,0.62470436,0.60908675,0.59346914,0.58175594,0.5661383,0.5505207,0.7418364,0.93315214,1.1283722,1.319688,1.5110037,1.5812829,1.6515622,1.7218413,1.7921207,1.8623998,1.6320401,1.4016805,1.1713207,0.94096094,0.7106012,0.98000497,1.2494087,1.5149081,1.7843118,2.0498111,2.6471848,3.2445583,3.8419318,4.4393053,5.036679,6.1494336,7.262188,8.374943,9.487698,10.600452,10.131924,9.659492,9.190963,8.718531,8.250002,7.898606,7.551114,7.1997175,6.8483214,6.5008297,5.2006636,3.9044023,2.6081407,1.3118792,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.07027924,0.14055848,0.21083772,0.28111696,0.3513962,0.6910792,1.0307622,1.3704453,1.7101282,2.0498111,1.639849,1.2298868,0.8199245,0.40996224,0.0,0.19912452,0.39434463,0.59346914,0.78868926,0.9878138,0.78868926,0.59346914,0.39434463,0.19912452,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.9097257,1.7686942,2.631567,3.4905357,4.349504,3.521771,2.690133,1.8584955,1.0307622,0.19912452,0.19131571,0.1796025,0.1717937,0.16008049,0.14836729,0.1835069,0.21474212,0.24597734,0.28111696,0.31235218,0.3318742,0.3474918,0.3631094,0.38263142,0.39824903,0.44119745,0.48414588,0.5270943,0.5700427,0.61299115,0.8667773,1.1205635,1.3782539,1.6320401,1.8858263,1.9756275,2.0615244,2.1513257,2.2372224,2.3231194,2.5456703,2.7643168,2.9868677,3.2055142,3.4241607,3.1469483,2.8697357,2.592523,2.3153105,2.0380979,2.3114061,2.5808098,2.854118,3.1274261,3.4007344,3.2992198,3.193801,3.0922866,2.9907722,2.8892577,3.2562714,3.6232853,3.9902992,4.357313,4.7243266,4.7633705,4.7985106,4.8375545,4.8765984,4.911738,5.036679,5.1616197,5.2865605,5.4115014,5.5364423,5.3295093,5.1225758,4.9156423,4.7087092,4.5017757,4.084005,3.6701381,3.2562714,2.8385005,2.4246337,2.1786566,1.9287747,1.6827974,1.43682,1.1869383,1.4016805,1.6164225,1.8311646,2.0459068,2.260649,2.241127,2.2216048,2.2020829,2.182561,2.1630387,2.3075018,2.4519646,2.5964274,2.7408905,2.8892577,3.4514916,4.01763,4.5837684,5.1460023,5.7121406,6.2197127,6.727285,7.2348576,7.7424297,8.250002,8.011833,7.773665,7.5394006,7.3012323,7.0630636,6.5633,6.0635366,5.563773,5.0640097,4.564246,4.903929,5.2436123,5.5832953,5.9229784,6.262661,6.036206,5.813655,5.5871997,5.3607445,5.138193,5.040583,4.9468775,4.853172,4.755562,4.661856,4.415879,4.173806,3.9278288,3.6818514,3.435874,3.6349986,3.8341231,4.029343,4.2284675,4.423688,4.5291066,4.6345253,4.7399445,4.845363,4.950782,4.903929,4.853172,4.806319,4.759466,4.7126136,4.435401,4.1581883,3.8809757,3.6037633,3.3265507,3.5686235,3.8106966,4.0527697,4.2948427,4.5369153,13.146122,21.751425,30.360632,38.965935,47.57514,44.998238,42.425236,39.848328,37.27533,34.69842,32.262077,29.82573,27.385477,24.949131,22.512783,19.143284,15.773785,12.404286,9.030883,5.661383,4.7009,3.736513,2.77603,1.8116426,0.8511597,0.76916724,0.6832704,0.60127795,0.5192855,0.43729305,0.737932,1.038571,1.33921,1.6359446,1.9365835,3.2055142,4.4705405,5.7394714,7.008402,8.273428,12.4511385,16.624945,20.79875,24.976461,29.150267,32.03562,34.920975,37.806328,40.69168,43.573128,39.40323,35.233326,31.063425,26.893522,22.723621,22.274614,21.82561,21.376602,20.92369,20.474686,20.787037,21.09939,21.411741,21.724094,22.036446,22.7041,23.371752,24.039404,24.707058,25.37471,21.407837,17.44487,13.477997,9.515028,5.548156,5.9815445,6.4110284,6.8405128,7.269997,7.699481,7.941554,8.179723,8.421796,8.659965,8.898132,9.198771,9.499411,9.80005,10.100689,10.401327,9.901564,9.405705,8.905942,8.410083,7.914223,8.714626,9.518932,10.319335,11.123642,11.924045,10.573121,9.218294,7.8673706,6.5164475,5.1616197,5.3256044,5.493494,5.657479,5.8214636,5.989353,5.7238536,5.462259,5.2006636,4.939069,4.6735697,3.970777,3.2640803,2.5612879,1.8545911,1.1517987,0.92924774,0.7106012,0.48805028,0.26940376,0.05075723,0.06637484,0.08589685,0.10151446,0.12103647,0.13665408,0.10932326,0.08199245,0.05466163,0.027330816,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.27721256,0.5036679,0.7340276,0.96048295,1.1869383,0.9917182,0.79649806,0.60127795,0.40605783,0.21083772,0.28111696,0.3474918,0.41386664,0.48414588,0.5505207,0.5192855,0.48414588,0.45291066,0.42167544,0.38653582,0.3709182,0.359205,0.3435874,0.3279698,0.31235218,0.30063897,0.29283017,0.28111696,0.27330816,0.26159495,0.38653582,0.5075723,0.62860876,0.75354964,0.8745861,0.97610056,1.0737107,1.175225,1.2767396,1.3743496,1.2064602,1.038571,0.8706817,0.7066968,0.5388075,0.4997635,0.46071947,0.42557985,0.38653582,0.3513962,1.3860629,2.4207294,3.455396,4.4900627,5.5247293,4.572055,3.619381,2.6667068,1.7140326,0.76135844,0.6754616,0.58566034,0.4997635,0.41386664,0.3240654,0.8941081,1.4641509,2.0341935,2.6042364,3.174279,3.8341231,4.4900627,5.1460023,5.805846,6.461786,5.298274,4.1308575,2.9673457,1.8038338,0.63641757,0.6715572,0.7027924,0.7340276,0.76916724,0.80040246,0.77307165,0.74574083,0.71841,0.6910792,0.6637484,0.7145056,0.76916724,0.8199245,0.8706817,0.92534333,0.92143893,0.92143893,0.91753453,0.9136301,0.9136301,0.80821127,0.7066968,0.60518235,0.5036679,0.39824903,1.4914817,2.5808098,3.6701381,4.759466,5.8487945,4.7204223,3.5881457,2.4597735,1.3314011,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.22645533,0.24988174,0.27330816,0.30063897,0.3240654,1.0463798,1.7686942,2.4910088,3.213323,3.9356375,4.322173,4.7087092,5.0913405,5.477876,5.8644123,5.833177,5.801942,5.7707067,5.743376,5.7121406,5.298274,4.8883114,4.474445,4.0605783,3.6506162,3.8067923,3.959064,4.11524,4.271416,4.423688,3.892689,3.3616903,2.8267872,2.2957885,1.7608855,1.9873407,2.2137961,2.436347,2.6628022,2.8892577,3.3890212,3.8887846,4.388548,4.8883114,5.388075,5.4036927,5.4193106,5.4310236,5.446641,5.462259,5.1499066,4.8375545,4.5252023,4.21285,3.900498,4.4510183,5.0054436,5.5559645,6.1103897,6.66091,7.309041,7.957172,8.605303,9.253433,9.901564,9.0152645,8.128965,7.2465706,6.3602715,5.473972,5.840986,6.2040954,6.571109,6.9342184,7.3012323,6.774138,6.250948,5.7238536,5.2006636,4.6735697,5.1225758,5.571582,6.016684,6.46569,6.910792,6.910792,6.9068875,6.9068875,6.902983,6.899079,6.4149327,5.930787,5.446641,4.958591,4.474445,4.5369153,4.5993857,4.661856,4.7243266,4.786797,4.7399445,4.6930914,4.646239,4.5993857,4.548629,4.6110992,4.6735697,4.73604,4.7985106,4.860981,4.8687897,4.872694,4.8765984,4.884407,4.8883114,4.173806,3.4593005,2.7408905,2.0263848,1.3118792,1.5812829,1.8506867,2.1239948,2.3933985,2.6628022,2.8306916,3.0024853,3.174279,3.3421683,3.513962,3.4788225,3.4436827,3.408543,3.3734035,3.338264,2.7330816,2.1318035,1.5305257,0.92924774,0.3240654,0.62470436,0.61299115,0.60127795,0.58566034,0.57394713,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.5505207,0.5388075,0.5231899,0.5114767,0.4997635,0.5231899,0.5505207,0.57394713,0.60127795,0.62470436,0.61299115,0.60127795,0.58566034,0.57394713,0.5622339,0.77307165,0.9878138,1.1986516,1.4133936,1.6242313,1.7140326,1.7999294,1.8858263,1.9756275,2.0615244,1.7608855,1.4641509,1.1635119,0.8628729,0.5622339,0.8745861,1.1869383,1.4992905,1.8116426,2.1239948,2.87364,3.6232853,4.376835,5.12648,5.8761253,6.98888,8.101635,9.21439,10.323239,11.435994,10.998701,10.561408,10.124115,9.686822,9.249529,8.823949,8.398369,7.9766936,7.551114,7.125534,5.700427,4.2753205,2.8502135,1.4251068,0.0,0.0,0.0,0.0,0.0,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.8628729,1.2884527,1.7140326,2.135708,2.5612879,2.0498111,1.5383345,1.0268579,0.5114767,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,1.0737107,2.0888553,3.1000953,4.1113358,5.12648,4.0996222,3.076669,2.0498111,1.0268579,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.18741131,0.24988174,0.31235218,0.37482262,0.43729305,0.47633708,0.5114767,0.5505207,0.58566034,0.62470436,0.9136301,1.1986516,1.4875772,1.7765031,2.0615244,2.0615244,2.0615244,2.0615244,2.0615244,2.0615244,2.3231194,2.5886188,2.8502135,3.1118085,3.3734035,2.9751544,2.5769055,2.174752,1.7765031,1.3743496,1.7491722,2.1239948,2.4988174,2.87364,3.2484627,3.1859922,3.1235218,3.0610514,2.998581,2.9361105,3.3734035,3.8106966,4.251894,4.689187,5.12648,4.985922,4.8492675,4.7126136,4.575959,4.4393053,4.7243266,5.0132523,5.298274,5.5871997,5.8761253,5.735567,5.5989127,5.462259,5.3256044,5.1889505,4.661856,4.138666,3.611572,3.0883822,2.5612879,2.2879796,2.0107672,1.737459,1.4641509,1.1869383,1.3626363,1.5383345,1.7140326,1.8858263,2.0615244,1.9873407,1.9131571,1.8389735,1.7608855,1.6867018,1.7999294,1.9131571,2.0263848,2.135708,2.2489357,2.6745155,3.1000953,3.5256753,3.951255,4.376835,5.036679,5.700427,6.364176,7.0240197,7.687768,7.6135845,7.5394006,7.461313,7.387129,7.3129454,6.649197,5.989353,5.3256044,4.661856,3.998108,4.3612175,4.7243266,5.087436,5.4505453,5.813655,5.5130157,5.212377,4.911738,4.6110992,4.3143644,4.1503797,3.9863946,3.8263142,3.6623292,3.4983444,3.4124475,3.3265507,3.2367494,3.1508527,3.0610514,3.2875066,3.513962,3.736513,3.9629683,4.1894236,4.224563,4.263607,4.298747,4.337791,4.376835,4.4510183,4.5252023,4.5993857,4.6735697,4.7516575,4.4119744,4.0761957,3.736513,3.4007344,3.0610514,3.076669,3.0883822,3.1000953,3.1118085,3.1235218,12.037272,20.951023,29.860868,38.77462,47.68837,43.776157,39.86395,35.951736,32.03562,28.12341,25.425468,22.723621,20.025679,17.323833,14.625891,12.962616,11.29934,9.636065,7.9766936,6.3134184,5.263134,4.21285,3.1625657,2.1122816,1.0619974,0.93705654,0.81211567,0.6871748,0.5622339,0.43729305,0.7106012,0.9878138,1.261122,1.5383345,1.8116426,3.4632049,5.1108627,6.7624245,8.413987,10.061645,14.161267,18.26089,22.364416,26.464039,30.563662,33.4373,36.31094,39.188484,42.062126,44.935764,39.29781,33.663757,28.025799,22.387842,16.749886,17.40192,18.05005,18.698183,19.350218,19.998348,20.79875,21.599154,22.399555,23.199959,24.00036,24.761719,25.523077,26.28834,27.049698,27.811058,22.938364,18.061766,13.189071,8.312472,3.435874,4.1620927,4.8883114,5.610626,6.336845,7.0630636,7.6370106,8.210958,8.78881,9.362757,9.936704,10.010887,10.088976,10.163159,10.237343,10.311526,9.811763,9.311999,8.812236,8.312472,7.812709,8.886419,9.964035,11.037745,12.111456,13.189071,11.748346,10.311526,8.874706,7.437886,6.001066,6.0635366,6.126007,6.1884775,6.250948,6.3134184,5.899552,5.4856853,5.0757227,4.661856,4.251894,3.5764325,2.900971,2.2255092,1.5500476,0.8745861,0.698888,0.5231899,0.3513962,0.1756981,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.3357786,0.3631094,0.38653582,0.41386664,0.43729305,0.41386664,0.38653582,0.3631094,0.3357786,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.38653582,0.46071947,0.5388075,0.61299115,0.6871748,0.77307165,0.8628729,0.94876975,1.038571,1.1244678,1.0268579,0.92534333,0.8238289,0.7262188,0.62470436,0.5505207,0.47633708,0.39824903,0.3240654,0.24988174,1.475864,2.7018464,3.9239242,5.1499066,6.375889,5.099149,3.8263142,2.5495746,1.2767396,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,1.0893283,1.7999294,2.514435,3.2250361,3.9356375,4.7516575,5.563773,6.375889,7.1880045,8.00012,6.5359693,5.0757227,3.611572,2.1513257,0.6871748,0.737932,0.78868926,0.8394465,0.8862993,0.93705654,0.8511597,0.76135844,0.6754616,0.58566034,0.4997635,0.62470436,0.74964523,0.8745861,0.999527,1.1244678,1.1010414,1.0737107,1.0502841,1.0268579,0.999527,0.9019169,0.80040246,0.698888,0.60127795,0.4997635,1.8623998,3.2250361,4.5876727,5.950309,7.3129454,5.899552,4.4861584,3.076669,1.6632754,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.27330816,0.30063897,0.3240654,0.3513962,0.37482262,1.1986516,2.0263848,2.8502135,3.6740425,4.5017757,4.9742084,5.4505453,5.9268827,6.3993154,6.8756523,6.8639393,6.8483214,6.8366084,6.824895,6.813182,6.1884775,5.563773,4.939069,4.3143644,3.6857557,3.4632049,3.2367494,3.0141985,2.787743,2.5612879,2.4129205,2.260649,2.1122816,1.9639144,1.8116426,1.9639144,2.1122816,2.260649,2.4129205,2.5612879,2.9361105,3.310933,3.6857557,4.0605783,4.4393053,4.6110992,4.786797,4.9624953,5.138193,5.3138914,5.0757227,4.8375545,4.5993857,4.3612175,4.123049,4.462732,4.7985106,5.138193,5.473972,5.813655,6.7233806,7.6370106,8.550641,9.464272,10.373997,9.413514,8.449126,7.4886436,6.524256,5.563773,6.1494336,6.7389984,7.3246584,7.914223,8.499884,7.898606,7.3012323,6.699954,6.098676,5.5013027,5.9268827,6.348558,6.774138,7.1997175,7.6252975,7.461313,7.3012323,7.137247,6.9732623,6.813182,6.223617,5.6379566,5.0483923,4.462732,3.873167,4.025439,4.173806,4.3260775,4.474445,4.6267166,4.6735697,4.7243266,4.775084,4.825841,4.8765984,4.8375545,4.7985106,4.7633705,4.7243266,4.689187,4.7633705,4.8375545,4.911738,4.985922,5.0640097,4.2753205,3.4866312,2.7018464,1.9131571,1.1244678,1.4641509,1.7999294,2.135708,2.475391,2.8111696,2.998581,3.1859922,3.3734035,3.5608149,3.7482262,3.7638438,3.775557,3.78727,3.7989833,3.8106966,3.0610514,2.3114061,1.5617609,0.81211567,0.062470436,0.62470436,0.61689556,0.60518235,0.59346914,0.58566034,0.57394713,0.58175594,0.58956474,0.59737355,0.60518235,0.61299115,0.60127795,0.58566034,0.57394713,0.5622339,0.5505207,0.58175594,0.60908675,0.64032197,0.6715572,0.698888,0.71841,0.7340276,0.75354964,0.76916724,0.78868926,1.0112402,1.2376955,1.4641509,1.6867018,1.9131571,1.9834363,2.05762,2.1318035,2.2020829,2.2762666,2.0498111,1.8233559,1.6008049,1.3743496,1.1517987,1.33921,1.5305257,1.7218413,1.9092526,2.1005683,2.87364,3.6467118,4.415879,5.1889505,5.9620223,7.0786815,8.1992445,9.315904,10.432563,11.549222,11.084598,10.619974,10.155351,9.690726,9.226103,9.261242,9.300286,9.339331,9.37447,9.413514,7.562827,5.7121406,3.8614538,2.0107672,0.1639849,0.12884527,0.09761006,0.06637484,0.031235218,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.9097257,1.4446288,1.979532,2.514435,3.049338,2.4402514,1.8311646,1.2181735,0.60908675,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.14446288,0.22645533,0.30844778,0.39434463,0.47633708,0.39824903,0.32016098,0.24207294,0.1639849,0.08589685,0.8941081,1.698415,2.5027218,3.3070288,4.1113358,3.408543,2.7057507,2.0068626,1.3040704,0.60127795,0.76526284,0.92924774,1.0932326,1.261122,1.4251068,1.2962615,1.1635119,1.0346665,0.9058213,0.77307165,0.8355421,0.8941081,0.95657855,1.0151446,1.0737107,1.0346665,0.9956226,0.95657855,0.9136301,0.8745861,1.1205635,1.3704453,1.6164225,1.8663043,2.1122816,2.1083772,2.1083772,2.1044729,2.1005683,2.1005683,2.2996929,2.4988174,2.7018464,2.900971,3.1000953,2.8463092,2.5886188,2.3348327,2.0810463,1.8233559,2.0459068,2.2684577,2.4910088,2.7135596,2.9361105,2.9634414,2.9868677,3.0141985,3.0376248,3.0610514,3.4632049,3.8614538,4.263607,4.661856,5.0640097,4.892216,4.7243266,4.552533,4.380739,4.21285,4.4393053,4.661856,4.8883114,5.1108627,5.337318,5.239708,5.142098,5.044488,4.9468775,4.8492675,4.423688,3.9942036,3.5686235,3.1391394,2.7135596,2.397303,2.0810463,1.7686942,1.4524376,1.1361811,1.2415999,1.3431144,1.4446288,1.5461433,1.6515622,1.6008049,1.5539521,1.5070993,1.4602464,1.4133936,1.5500476,1.6867018,1.8233559,1.9639144,2.1005683,2.4207294,2.7447948,3.06886,3.3890212,3.7130866,4.3612175,5.009348,5.6535745,6.3017054,6.949836,6.9927845,7.0357327,7.0786815,7.1216297,7.1606736,6.6413884,6.1221027,5.602817,5.083532,4.564246,4.8648853,5.169429,5.4700675,5.7707067,6.0752497,5.7902284,5.505207,5.2201858,4.9351645,4.650143,4.4588275,4.263607,4.0722914,3.8809757,3.6857557,3.5842414,3.4827268,3.3812122,3.2757936,3.174279,3.3616903,3.5451972,3.7287042,3.9161155,4.0996222,4.271416,4.4432096,4.618908,4.7907014,4.9624953,5.001539,5.036679,5.0757227,5.1108627,5.1499066,4.7985106,4.4510183,4.0996222,3.7482262,3.4007344,3.4905357,3.5803368,3.6701381,3.7599394,3.8497405,11.842052,19.834364,27.826675,35.818985,43.8113,40.8869,37.9625,35.038105,32.11371,29.189312,25.921326,22.653341,19.385357,16.117373,12.849388,11.674163,10.498938,9.323712,8.148487,6.9732623,6.3017054,5.630148,4.958591,4.283129,3.611572,3.533484,3.4514916,3.3734035,3.2914112,3.213323,3.5569105,3.8965936,4.240181,4.5837684,4.9234514,7.375416,9.823476,12.27544,14.723501,17.175465,19.98273,22.789995,25.597261,28.404526,31.211792,33.070286,34.928783,36.783375,38.64187,40.500366,35.8307,31.161034,26.49137,21.821705,17.148134,17.640089,18.12814,18.620094,19.108145,19.6001,20.63867,21.681147,22.719717,23.758287,24.800762,25.452799,26.104834,26.756868,27.408903,28.06094,23.047686,18.034433,13.017277,8.0040245,2.9868677,3.6623292,4.337791,5.0132523,5.688714,6.364176,7.0474463,7.7307167,8.4178915,9.101162,9.788337,9.792241,9.796145,9.803954,9.807858,9.811763,9.815667,9.823476,9.82738,9.8312845,9.839094,10.760532,11.681972,12.603411,13.528754,14.450192,12.86891,11.283723,9.702439,8.121157,6.5359693,6.348558,6.1611466,5.9737353,5.786324,5.5989127,5.173333,4.7516575,4.3260775,3.900498,3.474918,2.920493,2.366068,1.8116426,1.2533131,0.698888,0.5583295,0.42167544,0.28111696,0.14055848,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.07418364,0.07027924,0.06637484,0.06637484,0.062470436,0.06637484,0.06637484,0.07027924,0.07418364,0.07418364,0.12884527,0.1835069,0.23816854,0.29673457,0.3513962,0.3709182,0.39044023,0.40996224,0.42948425,0.44900626,0.42948425,0.40996224,0.39044023,0.3709182,0.3513962,0.3513962,0.3513962,0.3513962,0.3513962,0.3513962,0.40605783,0.46462387,0.5231899,0.58175594,0.63641757,0.6949836,0.75354964,0.80821127,0.8667773,0.92534333,0.8433509,0.76526284,0.6832704,0.60518235,0.5231899,0.47243267,0.42167544,0.3670138,0.31625658,0.26159495,1.2572175,2.25284,3.2484627,4.2440853,5.2358036,4.533011,3.8341231,3.1313305,2.4285383,1.7257458,1.4407244,1.1557031,0.8706817,0.58566034,0.30063897,0.9058213,1.5110037,2.1161861,2.7213683,3.3265507,4.126953,4.9234514,5.7238536,6.524256,7.3246584,6.0518236,4.775084,3.4983444,2.2255092,0.94876975,1.0034313,1.0541886,1.1088502,1.1596074,1.2142692,1.0854238,0.95657855,0.8316377,0.7027924,0.57394713,0.76526284,0.95657855,1.1439898,1.3353056,1.5266213,1.456342,1.3860629,1.3157835,1.2455044,1.175225,1.5070993,1.8389735,2.1708477,2.5066261,2.8385005,3.7326086,4.6267166,5.520825,6.4188375,7.3129454,5.9464045,4.5837684,3.2172275,1.8506867,0.48805028,0.41777104,0.3474918,0.27721256,0.20693332,0.13665408,0.10932326,0.08199245,0.05466163,0.027330816,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.21864653,0.23816854,0.26159495,0.28111696,0.30063897,0.96048295,1.620327,2.280171,2.9400148,3.5998588,4.084005,4.5681505,5.056201,5.5403466,6.0244927,6.098676,6.1767645,6.250948,6.3251314,6.3993154,5.938596,5.473972,5.0132523,4.548629,4.087909,3.853645,3.6232853,3.3890212,3.1586614,2.9243972,2.795552,2.6706111,2.541766,2.416825,2.2879796,2.338737,2.3855898,2.436347,2.4871042,2.5378613,2.912684,3.2875066,3.6623292,4.037152,4.4119744,4.5017757,4.5876727,4.6735697,4.7633705,4.8492675,4.6267166,4.4002614,4.173806,3.951255,3.7247996,4.2479897,4.7711797,5.2943697,5.813655,6.336845,6.9732623,7.6135845,8.250002,8.886419,9.526741,8.734148,7.941554,7.1489606,6.356367,5.563773,5.9737353,6.3836975,6.79366,7.2036223,7.6135845,7.238762,6.8639393,6.4891167,6.114294,5.735567,5.9659266,6.192382,6.4188375,6.649197,6.8756523,6.832704,6.7897553,6.746807,6.703859,6.66091,6.165051,5.6691923,5.169429,4.6735697,4.173806,4.1464753,4.1191444,4.0918136,4.0644827,4.037152,4.087909,4.138666,4.1894236,4.2362766,4.2870336,4.2362766,4.181615,4.1308575,4.0761957,4.025439,4.087909,4.1503797,4.21285,4.2753205,4.337791,3.6818514,3.0259118,2.3738766,1.717937,1.0619974,1.4212024,1.7843118,2.1435168,2.5027218,2.8619268,2.97125,3.076669,3.1859922,3.2914112,3.4007344,3.5491016,3.6935644,3.8419318,3.9902992,4.138666,3.6818514,3.2211318,2.7643168,2.3075018,1.8506867,0.62470436,0.61689556,0.60908675,0.60127795,0.59346914,0.58566034,0.60127795,0.61689556,0.63251317,0.6481308,0.6637484,0.6481308,0.63641757,0.62470436,0.61299115,0.60127795,0.63641757,0.6715572,0.7066968,0.7418364,0.77307165,0.8238289,0.8706817,0.91753453,0.96438736,1.0112402,1.2494087,1.4875772,1.7257458,1.9639144,2.1981785,2.2567444,2.3153105,2.3738766,2.4285383,2.4871042,2.338737,2.1864653,2.0380979,1.8858263,1.737459,1.8038338,1.8741131,1.9404879,2.0068626,2.0732377,2.8697357,3.6662338,4.4588275,5.2553253,6.0518236,7.172387,8.296855,9.4174185,10.541886,11.66245,11.170495,10.67854,10.186585,9.690726,9.198771,9.698535,10.198298,10.701966,11.20173,11.701493,9.425227,7.1489606,4.8765984,2.6003318,0.3240654,0.26159495,0.19522011,0.12884527,0.06637484,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.95657855,1.6008049,2.2489357,2.893162,3.5373883,2.8306916,2.1239948,1.4133936,0.7066968,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.28892577,0.45681506,0.62079996,0.78478485,0.94876975,0.78088045,0.61689556,0.44900626,0.28111696,0.113227665,0.7106012,1.3079748,1.9053483,2.5027218,3.1000953,2.7213683,2.338737,1.9600099,1.5812829,1.1986516,1.5188124,1.8350691,2.1513257,2.4714866,2.787743,2.514435,2.241127,1.9717231,1.698415,1.4251068,1.4836729,1.5383345,1.5969005,1.6554666,1.7140326,1.5969005,1.475864,1.358732,1.2415999,1.1244678,1.3314011,1.5383345,1.7491722,1.9561055,2.1630387,2.1591344,2.1513257,2.1474214,2.1435168,2.135708,2.2762666,2.4129205,2.5495746,2.6862288,2.8267872,2.7135596,2.6042364,2.494913,2.3855898,2.2762666,2.3465457,2.416825,2.4831998,2.5534792,2.6237583,2.736986,2.8502135,2.9634414,3.076669,3.1859922,3.5491016,3.912211,4.2753205,4.6384296,5.001539,4.7985106,4.5954814,4.3924527,4.1894236,3.9863946,4.1503797,4.3143644,4.474445,4.6384296,4.7985106,4.743849,4.6852827,4.6267166,4.5681505,4.513489,4.181615,3.853645,3.521771,3.193801,2.8619268,2.5066261,2.1513257,1.796025,1.4407244,1.0893283,1.116659,1.1478943,1.1791295,1.2064602,1.2376955,1.2181735,1.1986516,1.1791295,1.1557031,1.1361811,1.3001659,1.4641509,1.6242313,1.7882162,1.9482968,2.1708477,2.3894942,2.6081407,2.8306916,3.049338,3.6818514,4.3143644,4.9468775,5.579391,6.211904,6.3719845,6.532065,6.6921453,6.852226,7.012306,6.6335793,6.2587566,5.8800297,5.5013027,5.12648,5.368553,5.610626,5.852699,6.094772,6.336845,6.067441,5.7980375,5.5286336,5.2592297,4.985922,4.7633705,4.5408196,4.318269,4.095718,3.873167,3.7560349,3.638903,3.521771,3.4046388,3.2875066,3.4319696,3.5764325,3.7208953,3.8692627,4.0137253,4.318269,4.6267166,4.9351645,5.2436123,5.548156,5.548156,5.548156,5.548156,5.548156,5.548156,5.1889505,4.825841,4.462732,4.0996222,3.736513,3.9044023,4.0722914,4.240181,4.40807,4.575959,11.6468315,18.72161,25.79248,32.863354,39.93813,38.00155,36.061058,34.124477,32.187893,30.251308,26.41328,22.579159,18.745035,14.9109125,11.076789,10.38571,9.698535,9.01136,8.324185,7.6370106,7.3441806,7.0474463,6.7507114,6.4578815,6.1611466,6.126007,6.0908675,6.055728,6.0205884,5.989353,6.3993154,6.8092775,7.2192397,7.629202,8.039165,11.287627,14.53609,17.788456,21.036919,24.289286,25.804195,27.319103,28.834011,30.348919,31.863827,32.703274,33.54272,34.382168,35.22161,36.061058,32.359688,28.658312,24.953035,21.251661,17.550287,17.878258,18.210133,18.538101,18.869976,19.20185,20.47859,21.759233,23.039877,24.320522,25.601166,26.143877,26.68659,27.229301,27.768108,28.310822,23.15701,18.003199,12.845484,7.6916723,2.5378613,3.1625657,3.78727,4.4119744,5.036679,5.661383,6.4578815,7.2543793,8.046973,8.843472,9.636065,9.573594,9.507219,9.440845,9.378374,9.311999,9.823476,10.331048,10.8425255,11.354002,11.861574,12.630741,13.403813,14.17298,14.942147,15.711315,13.985569,12.2559185,10.530173,8.804427,7.0747766,6.6374836,6.2001905,5.7628975,5.3256044,4.8883114,4.4510183,4.0137253,3.5764325,3.1391394,2.7018464,2.2645533,1.8311646,1.3938715,0.96048295,0.5231899,0.42167544,0.31625658,0.21083772,0.10541886,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.093705654,0.10151446,0.10932326,0.11713207,0.12494087,0.12884527,0.13665408,0.14055848,0.14446288,0.14836729,0.19912452,0.24597734,0.29283017,0.339683,0.38653582,0.40215343,0.41777104,0.43338865,0.44900626,0.46071947,0.44900626,0.43338865,0.41777104,0.40215343,0.38653582,0.38653582,0.38653582,0.38653582,0.38653582,0.38653582,0.42557985,0.46852827,0.5075723,0.5466163,0.58566034,0.61689556,0.6442264,0.6715572,0.698888,0.7262188,0.6637484,0.60518235,0.5466163,0.48414588,0.42557985,0.39434463,0.3631094,0.3357786,0.30454338,0.27330816,1.038571,1.8038338,2.5690966,3.3343596,4.0996222,3.970777,3.8419318,3.7091823,3.5803368,3.4514916,2.803361,2.1591344,1.5149081,0.8706817,0.22645533,0.7223144,1.2181735,1.717937,2.2137961,2.7135596,3.4983444,4.2870336,5.0757227,5.8644123,6.649197,5.563773,4.474445,3.3890212,2.2996929,1.2142692,1.2689307,1.3235924,1.3782539,1.4329157,1.4875772,1.319688,1.1517987,0.98390937,0.8160201,0.6481308,0.9058213,1.1596074,1.4133936,1.6710842,1.9248703,1.8116426,1.6945106,1.5812829,1.4641509,1.3509232,2.1161861,2.8814487,3.6467118,4.4119744,5.173333,5.602817,6.028397,6.4578815,6.883461,7.3129454,5.9932575,4.677474,3.3616903,2.0420024,0.7262188,0.63641757,0.5466163,0.45681506,0.3631094,0.27330816,0.21864653,0.1639849,0.10932326,0.05466163,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.1639849,0.1796025,0.19522011,0.21083772,0.22645533,0.71841,1.2142692,1.7101282,2.2059872,2.7018464,3.193801,3.68966,4.185519,4.6813784,5.173333,5.337318,5.5013027,5.661383,5.825368,5.989353,5.688714,5.388075,5.087436,4.786797,4.4861584,4.2479897,4.0059166,3.767748,3.5256753,3.2875066,3.182088,3.076669,2.97125,2.8658314,2.7643168,2.7135596,2.6628022,2.612045,2.5612879,2.514435,2.8892577,3.2640803,3.638903,4.0137253,4.388548,4.388548,4.388548,4.388548,4.388548,4.388548,4.173806,3.9629683,3.7482262,3.5373883,3.3265507,4.0332475,4.7399445,5.446641,6.153338,6.8639393,7.223144,7.5862536,7.9493628,8.312472,8.675582,8.050878,7.4300776,6.8092775,6.184573,5.563773,5.794133,6.028397,6.2587566,6.493021,6.7233806,6.575013,6.426646,6.2743745,6.126007,5.9737353,6.0049706,6.036206,6.0635366,6.094772,6.126007,6.2040954,6.278279,6.356367,6.434455,6.5125427,6.1064854,5.6965227,5.290465,4.884407,4.474445,4.271416,4.0644827,3.8614538,3.6545205,3.4514916,3.4983444,3.5491016,3.5998588,3.6506162,3.7013733,3.631094,3.5647192,3.4983444,3.4280653,3.3616903,3.4124475,3.4632049,3.513962,3.5608149,3.611572,3.0883822,2.5690966,2.0459068,1.5227169,0.999527,1.3821584,1.7647898,2.1474214,2.5300527,2.912684,2.9400148,2.9673457,2.9946766,3.0220075,3.049338,3.3343596,3.6154766,3.8965936,4.181615,4.462732,4.298747,4.1308575,3.9668727,3.802888,3.638903,0.62470436,0.62079996,0.61689556,0.60908675,0.60518235,0.60127795,0.62079996,0.6442264,0.6676528,0.6910792,0.7106012,0.698888,0.6871748,0.6754616,0.6637484,0.6481308,0.6910792,0.7301232,0.76916724,0.80821127,0.8511597,0.92924774,1.0034313,1.0815194,1.1596074,1.2376955,1.4875772,1.737459,1.9873407,2.2372224,2.4871042,2.5300527,2.5730011,2.6159496,2.6588979,2.7018464,2.6237583,2.5495746,2.475391,2.4012074,2.3231194,2.2684577,2.2137961,2.1591344,2.1044729,2.0498111,2.8658314,3.6857557,4.5017757,5.3217,6.13772,7.266093,8.39056,9.518932,10.647305,11.775677,11.256392,10.733202,10.213917,9.694631,9.175345,10.135828,11.100216,12.0606985,13.025085,13.985569,11.287627,8.58578,5.8878384,3.1859922,0.48805028,0.39044023,0.29283017,0.19522011,0.09761006,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,1.0034313,1.7608855,2.514435,3.2718892,4.025439,3.2211318,2.416825,1.6086137,0.80430686,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.43338865,0.6832704,0.92924774,1.1791295,1.4251068,1.1674163,0.9097257,0.6520352,0.39434463,0.13665408,0.5270943,0.91753453,1.3079748,1.698415,2.0888553,2.0302892,1.9717231,1.9131571,1.8584955,1.7999294,2.2684577,2.7408905,3.2094188,3.6818514,4.1503797,3.736513,3.3187418,2.9048753,2.4910088,2.0732377,2.1318035,2.1864653,2.241127,2.2957885,2.35045,2.15523,1.9600099,1.7647898,1.5695697,1.3743496,1.542239,1.7101282,1.8780174,2.0459068,2.2137961,2.2059872,2.1981785,2.1903696,2.182561,2.174752,2.2489357,2.3231194,2.4012074,2.475391,2.5495746,2.5847144,2.619854,2.6549935,2.690133,2.7252727,2.6432803,2.5612879,2.4792955,2.3933985,2.3114061,2.514435,2.7135596,2.912684,3.1118085,3.310933,3.638903,3.9629683,4.2870336,4.6110992,4.939069,4.7009,4.466636,4.2323723,3.998108,3.7638438,3.8614538,3.9629683,4.0605783,4.1620927,4.263607,4.2440853,4.2284675,4.2089458,4.193328,4.173806,3.9434462,3.7091823,3.4788225,3.2445583,3.0141985,2.6159496,2.2216048,1.8272603,1.4329157,1.038571,0.9956226,0.95267415,0.9097257,0.8667773,0.8238289,0.8316377,0.8394465,0.8472553,0.8550641,0.8628729,1.0502841,1.2376955,1.4251068,1.6125181,1.7999294,1.9170616,2.0341935,2.1513257,2.2684577,2.3855898,3.0063896,3.6232853,4.240181,4.8570766,5.473972,5.7511845,6.028397,6.3056097,6.5867267,6.8639393,6.6257706,6.3915067,6.1572423,5.9229784,5.688714,5.8683167,6.0518236,6.2353306,6.4188375,6.5984397,6.3446536,6.0908675,5.833177,5.579391,5.3256044,5.0718184,4.8219366,4.5681505,4.3143644,4.0605783,3.9317331,3.7989833,3.6662338,3.533484,3.4007344,3.506153,3.611572,3.7130866,3.8185053,3.9239242,4.369026,4.8102236,5.251421,5.6965227,6.13772,6.098676,6.0635366,6.0244927,5.989353,5.950309,5.575486,5.2006636,4.825841,4.4510183,4.0761957,4.318269,4.564246,4.8102236,5.056201,5.298274,11.4516115,17.60495,23.758287,29.911625,36.061058,35.11229,34.16352,33.210846,32.262077,31.313307,26.90914,22.508879,18.104713,13.700547,9.300286,9.101162,8.898132,8.699008,8.499884,8.300759,8.382751,8.464745,8.546737,8.628729,8.710721,8.722435,8.734148,8.741957,8.75367,8.761478,9.24172,9.718058,10.194394,10.670732,11.150972,15.199838,19.248703,23.301472,27.350338,31.399202,31.621754,31.844305,32.066856,32.289406,32.51196,32.336258,32.15666,31.980959,31.801357,31.625658,28.888672,26.15559,23.418604,20.685524,17.948538,18.12033,18.28822,18.460014,18.631807,18.799696,20.31851,21.841227,23.360039,24.87885,26.401567,26.831053,27.26444,27.69783,28.131218,28.560703,23.266333,17.971964,12.677594,7.3832245,2.0888553,2.6628022,3.2367494,3.8106966,4.388548,4.9624953,5.8683167,6.774138,7.676055,8.581876,9.487698,9.351044,9.218294,9.081639,8.94889,8.812236,9.82738,10.8425255,11.85767,12.872814,13.887959,14.504854,15.12175,15.738646,16.359446,16.976341,15.102228,13.228115,11.357906,9.483793,7.6135845,6.9264097,6.239235,5.548156,4.860981,4.173806,3.7247996,3.2757936,2.8267872,2.3738766,1.9248703,1.6086137,1.2962615,0.98000497,0.6637484,0.3513962,0.28111696,0.21083772,0.14055848,0.07027924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.11713207,0.13665408,0.15227169,0.1717937,0.18741131,0.19522011,0.20302892,0.21083772,0.21864653,0.22645533,0.26549935,0.30454338,0.3435874,0.38653582,0.42557985,0.43338865,0.44510186,0.45681506,0.46462387,0.47633708,0.46462387,0.45681506,0.44510186,0.43338865,0.42557985,0.42557985,0.42557985,0.42557985,0.42557985,0.42557985,0.44900626,0.46852827,0.49195468,0.5153811,0.5388075,0.5349031,0.5309987,0.5309987,0.5270943,0.5231899,0.48414588,0.44510186,0.40605783,0.3631094,0.3240654,0.31625658,0.30844778,0.30063897,0.29673457,0.28892577,0.8238289,1.358732,1.893635,2.4285383,2.9634414,3.4046388,3.8458362,4.290938,4.732136,5.173333,4.169902,3.1664703,2.1591344,1.1557031,0.14836729,0.5388075,0.92924774,1.319688,1.7101282,2.1005683,2.87364,3.6506162,4.423688,5.2006636,5.9737353,5.0757227,4.173806,3.2757936,2.3738766,1.475864,1.53443,1.5890918,1.6476578,1.7062237,1.7608855,1.5539521,1.3470187,1.1400855,0.93315214,0.7262188,1.0463798,1.3665408,1.6867018,2.0068626,2.3231194,2.1630387,2.0068626,1.8467822,1.6867018,1.5266213,2.7213683,3.9200199,5.1186714,6.3134184,7.5120697,7.473026,7.433982,7.3910336,7.3519893,7.3129454,6.044015,4.7711797,3.5022488,2.233318,0.96438736,0.8511597,0.7418364,0.63251317,0.5231899,0.41386664,0.3318742,0.24597734,0.1639849,0.08199245,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.10932326,0.12103647,0.12884527,0.14055848,0.14836729,0.48024148,0.80821127,1.1400855,1.4719596,1.7999294,2.3035975,2.8111696,3.3148375,3.8185053,4.3260775,4.575959,4.825841,5.0757227,5.3256044,5.575486,5.4388323,5.298274,5.1616197,5.024966,4.8883114,4.6384296,4.3924527,4.1464753,3.8965936,3.6506162,3.5686235,3.4866312,3.4007344,3.3187418,3.2367494,3.0883822,2.9361105,2.787743,2.639376,2.4871042,2.8619268,3.2367494,3.611572,3.9863946,4.3612175,4.2753205,4.1894236,4.0996222,4.0137253,3.9239242,3.7247996,3.5256753,3.3265507,3.1235218,2.9243972,3.8185053,4.7087092,5.602817,6.493021,7.387129,7.47693,7.562827,7.648724,7.7385254,7.824422,7.3715115,6.918601,6.46569,6.016684,5.563773,5.618435,5.6730967,5.727758,5.7824197,5.8370814,5.911265,5.989353,6.0635366,6.13772,6.211904,6.044015,5.8761253,5.708236,5.5442514,5.376362,5.571582,5.7707067,5.9659266,6.165051,6.364176,6.044015,5.727758,5.4115014,5.0913405,4.775084,4.3924527,4.009821,3.6271896,3.2445583,2.8619268,2.912684,2.9634414,3.0141985,3.0610514,3.1118085,3.0298162,2.9478238,2.8658314,2.7838387,2.7018464,2.736986,2.77603,2.8111696,2.8502135,2.8892577,2.4988174,2.1083772,1.717937,1.3274968,0.93705654,1.3431144,1.7491722,2.1513257,2.5573835,2.9634414,2.9087796,2.8580225,2.803361,2.7526035,2.7018464,3.1157131,3.533484,3.951255,4.369026,4.786797,4.9156423,5.040583,5.169429,5.298274,5.423215,0.62470436,0.62079996,0.62079996,0.61689556,0.61689556,0.61299115,0.6442264,0.6715572,0.7027924,0.7340276,0.76135844,0.74964523,0.737932,0.7262188,0.7106012,0.698888,0.74574083,0.78868926,0.8355421,0.8784905,0.92534333,1.0307622,1.1400855,1.2494087,1.3548276,1.4641509,1.7257458,1.9873407,2.2489357,2.514435,2.77603,2.803361,2.8306916,2.8580225,2.8853533,2.912684,2.912684,2.912684,2.912684,2.912684,2.912684,2.7330816,2.5573835,2.3816853,2.2020829,2.0263848,2.8658314,3.7052777,4.5447245,5.3841705,6.223617,7.355894,8.488171,9.6243515,10.756628,11.888905,11.338385,10.791768,10.2451515,9.698535,9.151918,10.573121,11.998228,13.423335,14.848442,16.273548,13.150026,10.0265045,6.899079,3.775557,0.6481308,0.5192855,0.39044023,0.26159495,0.12884527,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,1.0541886,1.9170616,2.7838387,3.6467118,4.513489,3.611572,2.7057507,1.8038338,0.9019169,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.58175594,0.9097257,1.2415999,1.5695697,1.901444,1.5539521,1.2064602,0.8589685,0.5114767,0.1639849,0.3435874,0.5270943,0.7106012,0.8941081,1.0737107,1.33921,1.6047094,1.8702087,2.135708,2.4012074,3.0220075,3.6467118,4.267512,4.8883114,5.5130157,4.9546866,4.396357,3.8419318,3.2836022,2.7252727,2.77603,2.8306916,2.8814487,2.9361105,2.9868677,2.7135596,2.4441557,2.1708477,1.8975395,1.6242313,1.7530766,1.8819219,2.0068626,2.135708,2.260649,2.25284,2.241127,2.233318,2.2216048,2.2137961,2.2255092,2.2372224,2.2489357,2.260649,2.2762666,2.455869,2.6354716,2.815074,2.9946766,3.174279,2.9400148,2.7057507,2.4714866,2.233318,1.999054,2.2879796,2.5769055,2.8619268,3.1508527,3.435874,3.7247996,4.0137253,4.298747,4.5876727,4.8765984,4.607195,4.3416953,4.0722914,3.8067923,3.5373883,3.5764325,3.611572,3.6506162,3.6857557,3.7247996,3.7482262,3.7716527,3.7911747,3.814601,3.8380275,3.7013733,3.5686235,3.4319696,3.2992198,3.1625657,2.7291772,2.2918842,1.8584955,1.4212024,0.9878138,0.8706817,0.75745404,0.6442264,0.5270943,0.41386664,0.44900626,0.48414588,0.5192855,0.5544251,0.58566034,0.80040246,1.0112402,1.2259823,1.43682,1.6515622,1.6632754,1.678893,1.6945106,1.7101282,1.7257458,2.3270237,2.9283018,3.533484,4.134762,4.73604,5.134289,5.5286336,5.9229784,6.3173227,6.7116675,6.621866,6.5281606,6.434455,6.3407493,6.250948,6.3719845,6.4969254,6.617962,6.7389984,6.8639393,6.621866,6.3836975,6.141625,5.903456,5.661383,5.380266,5.099149,4.814128,4.533011,4.251894,4.1035266,3.9551594,3.8067923,3.6584249,3.513962,3.5764325,3.6428072,3.7091823,3.7716527,3.8380275,4.415879,4.9937305,5.571582,6.1494336,6.7233806,6.649197,6.575013,6.5008297,6.426646,6.348558,5.9620223,5.575486,5.1889505,4.7985106,4.4119744,4.73604,5.056201,5.380266,5.704332,6.0244927,11.256392,16.48829,21.724094,26.955994,32.187893,32.22303,32.262077,32.30112,32.336258,32.375305,27.404999,22.434696,17.464392,12.494087,7.523783,7.812709,8.101635,8.386656,8.675582,8.960603,9.421323,9.882042,10.342762,10.803481,11.2642,11.318862,11.373524,11.428185,11.482847,11.537509,12.084125,12.626837,13.173453,13.716166,14.262781,19.11205,23.961317,28.81449,33.663757,38.513023,37.44322,36.373413,35.303604,34.2338,33.163994,31.969246,30.770594,29.575848,28.3811,27.186354,25.421562,23.652868,21.884174,20.119385,18.35069,18.3585,18.370213,18.381926,18.389734,18.401447,20.158428,21.919313,23.6802,25.441086,27.198067,27.522131,27.846197,28.166357,28.490423,28.810585,23.375656,17.94073,12.5058,7.0708723,1.6359446,2.1630387,2.6862288,3.213323,3.736513,4.263607,5.278752,6.2938967,7.309041,8.324185,9.339331,9.132397,8.929368,8.722435,8.519405,8.312472,9.8312845,11.354002,12.872814,14.391626,15.914344,16.378967,16.843592,17.308216,17.772839,18.237463,16.218887,14.204215,12.185639,10.167064,8.148487,7.211431,6.2743745,5.337318,4.4002614,3.4632049,2.998581,2.5378613,2.0732377,1.6125181,1.1517987,0.95657855,0.76135844,0.5661383,0.3709182,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.14055848,0.1678893,0.19522011,0.22255093,0.24988174,0.26159495,0.26940376,0.28111696,0.28892577,0.30063897,0.3318742,0.3631094,0.39824903,0.42948425,0.46071947,0.46852827,0.47243267,0.47633708,0.48414588,0.48805028,0.48414588,0.47633708,0.47243267,0.46852827,0.46071947,0.46071947,0.46071947,0.46071947,0.46071947,0.46071947,0.46852827,0.47243267,0.47633708,0.48414588,0.48805028,0.45681506,0.42167544,0.39044023,0.359205,0.3240654,0.30454338,0.28502136,0.26549935,0.24597734,0.22645533,0.23816854,0.25378615,0.26940376,0.28502136,0.30063897,0.60518235,0.9097257,1.2142692,1.5188124,1.8233559,2.8385005,3.853645,4.8687897,5.883934,6.899079,5.5364423,4.169902,2.803361,1.4407244,0.07418364,0.359205,0.64032197,0.92143893,1.2064602,1.4875772,2.2489357,3.0141985,3.775557,4.5369153,5.298274,4.5876727,3.873167,3.1625657,2.4480603,1.737459,1.796025,1.8584955,1.9170616,1.9756275,2.0380979,1.7882162,1.542239,1.2962615,1.0463798,0.80040246,1.1869383,1.5695697,1.9561055,2.338737,2.7252727,2.5183394,2.3153105,2.1083772,1.9053483,1.698415,3.330455,4.958591,6.590631,8.218767,9.850807,9.343235,8.835662,8.32809,7.8205175,7.3129454,6.0908675,4.8687897,3.6467118,2.4207294,1.1986516,1.0698062,0.94096094,0.80821127,0.679366,0.5505207,0.44119745,0.3318742,0.21864653,0.10932326,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05466163,0.058566034,0.06637484,0.07027924,0.07418364,0.23816854,0.40605783,0.5700427,0.7340276,0.9019169,1.4133936,1.9287747,2.4441557,2.959537,3.474918,3.8106966,4.1503797,4.4861584,4.825841,5.1616197,5.1889505,5.212377,5.2358036,5.263134,5.2865605,5.0327744,4.7789884,4.521298,4.267512,4.0137253,3.951255,3.892689,3.8341231,3.7716527,3.7130866,3.4632049,3.213323,2.9634414,2.7135596,2.463678,2.8385005,3.213323,3.5881457,3.9629683,4.337791,4.1620927,3.9863946,3.8106966,3.638903,3.4632049,3.2757936,3.0883822,2.900971,2.7135596,2.5261483,3.6037633,4.6813784,5.758993,6.8366084,7.914223,7.726812,7.5394006,7.348085,7.1606736,6.9732623,6.6921453,6.4110284,6.126007,5.84489,5.563773,5.4388323,5.3177958,5.196759,5.0718184,4.950782,5.251421,5.548156,5.8487945,6.1494336,6.4500723,6.083059,5.7199492,5.35684,4.989826,4.6267166,4.942973,5.2592297,5.579391,5.8956475,6.211904,5.985449,5.758993,5.5286336,5.3021784,5.0757227,4.513489,3.9551594,3.39683,2.8345962,2.2762666,2.3231194,2.3738766,2.4246337,2.475391,2.5261483,2.4285383,2.330928,2.233318,2.135708,2.0380979,2.0615244,2.0888553,2.1122816,2.135708,2.1630387,1.9053483,1.6476578,1.3899672,1.1322767,0.8745861,1.3040704,1.7296503,2.1591344,2.5847144,3.0141985,2.8814487,2.7486992,2.6159496,2.4831998,2.35045,2.900971,3.455396,4.0059166,4.560342,5.1108627,5.532538,5.9542136,6.3719845,6.79366,7.211431,0.62470436,0.62470436,0.62470436,0.62470436,0.62470436,0.62470436,0.6637484,0.698888,0.737932,0.77307165,0.81211567,0.80040246,0.78868926,0.77307165,0.76135844,0.74964523,0.80040246,0.8511597,0.9019169,0.94876975,0.999527,1.1361811,1.2767396,1.4133936,1.5500476,1.6867018,1.9639144,2.2372224,2.514435,2.787743,3.0610514,3.076669,3.0883822,3.1000953,3.1118085,3.1235218,3.2016098,3.2757936,3.349977,3.4241607,3.4983444,3.2016098,2.900971,2.6003318,2.2996929,1.999054,2.8619268,3.7247996,4.5876727,5.4505453,6.3134184,7.4495993,8.58578,9.725866,10.862047,11.998228,11.424281,10.850334,10.276386,9.698535,9.124588,11.014318,12.900145,14.785972,16.675701,18.56153,15.012426,11.4633255,7.914223,4.3612175,0.81211567,0.6481308,0.48805028,0.3240654,0.1639849,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,1.1010414,2.0732377,3.049338,4.025439,5.001539,3.998108,2.998581,1.999054,0.999527,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.7262188,1.1361811,1.5500476,1.9639144,2.3738766,1.9365835,1.4992905,1.0619974,0.62470436,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.6481308,1.2376955,1.8233559,2.4129205,2.998581,3.775557,4.548629,5.3256044,6.098676,6.8756523,6.1767645,5.473972,4.775084,4.0761957,3.3734035,3.4241607,3.474918,3.5256753,3.5764325,3.6232853,3.2757936,2.9243972,2.5769055,2.2255092,1.8741131,1.9639144,2.0498111,2.135708,2.2255092,2.3114061,2.2996929,2.2879796,2.2762666,2.260649,2.2489357,2.1981785,2.1513257,2.1005683,2.0498111,1.999054,2.3231194,2.6510892,2.9751544,3.2992198,3.6232853,3.2367494,2.8502135,2.463678,2.0732377,1.6867018,2.0615244,2.436347,2.8111696,3.1859922,3.5608149,3.8106966,4.0605783,4.3143644,4.564246,4.814128,4.513489,4.21285,3.912211,3.611572,3.310933,3.2875066,3.2640803,3.2367494,3.213323,3.1859922,3.2484627,3.310933,3.3734035,3.435874,3.4983444,3.4632049,3.4241607,3.3890212,3.349977,3.310933,2.8385005,2.3621633,1.8858263,1.4133936,0.93705654,0.74964523,0.5622339,0.37482262,0.18741131,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.5505207,0.78868926,1.0268579,1.261122,1.4992905,1.4133936,1.3235924,1.2376955,1.1517987,1.0619974,1.6515622,2.2372224,2.8267872,3.4124475,3.998108,4.513489,5.024966,5.5364423,6.0518236,6.5633,6.6140575,6.66091,6.7116675,6.7624245,6.813182,6.8756523,6.9381227,7.000593,7.0630636,7.125534,6.899079,6.676528,6.4500723,6.223617,6.001066,5.688714,5.376362,5.0640097,4.7516575,4.4393053,4.2753205,4.1113358,3.951255,3.78727,3.6232853,3.6506162,3.6740425,3.7013733,3.7247996,3.7482262,4.462732,5.173333,5.8878384,6.5984397,7.3129454,7.1997175,7.08649,6.9732623,6.8639393,6.7507114,6.348558,5.950309,5.548156,5.1499066,4.7516575,5.1499066,5.548156,5.950309,6.348558,6.7507114,11.061172,15.375536,19.685997,24.00036,28.310822,29.337679,30.360632,31.38749,32.41435,33.4373,27.900858,22.364416,16.82407,11.287627,5.7511845,6.524256,7.3012323,8.074304,8.85128,9.6243515,10.4637985,11.29934,12.138786,12.974329,13.813775,13.911386,14.012899,14.114414,14.212025,14.313539,14.92653,15.535617,16.148607,16.761599,17.37459,23.02426,28.673931,34.3236,39.97327,45.626846,43.260777,40.898613,38.53645,36.174286,33.812122,31.598328,29.388435,27.17464,24.960844,22.750952,21.95055,21.150146,20.349745,19.549341,18.74894,18.600573,18.448301,18.299932,18.151566,17.999294,19.998348,22.001307,24.00036,25.999414,27.998468,28.213211,28.42405,28.63879,28.849628,29.064371,23.488884,17.913397,12.337912,6.7624245,1.1869383,1.6632754,2.135708,2.612045,3.0883822,3.5608149,4.689187,5.813655,6.9381227,8.062591,9.187058,8.913751,8.636538,8.36323,8.086017,7.812709,9.839094,11.861574,13.887959,15.914344,17.936825,18.249176,18.56153,18.87388,19.186234,19.498585,17.335546,15.176412,13.013372,10.850334,8.687295,7.5003567,6.3134184,5.12648,3.9356375,2.7486992,2.2762666,1.7999294,1.3235924,0.8511597,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.1639849,0.19912452,0.23816854,0.27330816,0.31235218,0.3240654,0.3357786,0.3513962,0.3631094,0.37482262,0.39824903,0.42557985,0.44900626,0.47633708,0.4997635,0.4997635,0.4997635,0.4997635,0.4997635,0.4997635,0.4997635,0.4997635,0.4997635,0.4997635,0.4997635,0.4997635,0.4997635,0.4997635,0.4997635,0.4997635,0.48805028,0.47633708,0.46071947,0.44900626,0.43729305,0.37482262,0.31235218,0.24988174,0.18741131,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.1639849,0.19912452,0.23816854,0.27330816,0.31235218,0.38653582,0.46071947,0.5388075,0.61299115,0.6871748,2.2762666,3.8614538,5.4505453,7.0357327,8.624825,6.899079,5.173333,3.4514916,1.7257458,0.0,0.1756981,0.3513962,0.5231899,0.698888,0.8745861,1.6242313,2.3738766,3.1235218,3.873167,4.6267166,4.0996222,3.5764325,3.049338,2.5261483,1.999054,2.0615244,2.1239948,2.1864653,2.2489357,2.3114061,2.0263848,1.737459,1.4485333,1.1635119,0.8745861,1.3235924,1.7765031,2.2255092,2.6745155,3.1235218,2.87364,2.6237583,2.3738766,2.1239948,1.8741131,3.9395418,6.001066,8.062591,10.124115,12.185639,11.213444,10.237343,9.261242,8.289046,7.3129454,6.13772,4.9624953,3.78727,2.612045,1.43682,1.2884527,1.1361811,0.9878138,0.8394465,0.6871748,0.5505207,0.41386664,0.27330816,0.13665408,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5231899,1.0502841,1.5734742,2.1005683,2.6237583,3.049338,3.474918,3.900498,4.3260775,4.7516575,4.939069,5.12648,5.3138914,5.5013027,5.688714,5.423215,5.1616197,4.900025,4.6384296,4.376835,4.337791,4.298747,4.263607,4.224563,4.1894236,3.8380275,3.4866312,3.1391394,2.787743,2.436347,2.8111696,3.1859922,3.5608149,3.9356375,4.3143644,4.0488653,3.78727,3.5256753,3.2640803,2.998581,2.8267872,2.6510892,2.475391,2.2996929,2.1239948,3.3890212,4.650143,5.911265,7.1762915,8.437413,7.9766936,7.5120697,7.0513506,6.5867267,6.126007,6.012779,5.899552,5.786324,5.6730967,5.563773,5.263134,4.9624953,4.661856,4.3612175,4.0605783,4.5876727,5.1108627,5.6379566,6.1611466,6.688241,6.126007,5.563773,5.001539,4.4393053,3.873167,4.3143644,4.7516575,5.1889505,5.6262436,6.0635366,5.9268827,5.786324,5.64967,5.5130157,5.376362,4.6384296,3.900498,3.1625657,2.4246337,1.6867018,1.737459,1.7882162,1.8389735,1.8858263,1.9365835,1.8233559,1.7140326,1.6008049,1.4875772,1.3743496,1.3860629,1.4016805,1.4133936,1.4251068,1.43682,1.3118792,1.1869383,1.0619974,0.93705654,0.81211567,1.261122,1.7140326,2.1630387,2.612045,3.0610514,2.8502135,2.639376,2.4246337,2.2137961,1.999054,2.6862288,3.3734035,4.0605783,4.7516575,5.4388323,6.1494336,6.8639393,7.57454,8.289046,8.999647,0.6481308,0.6481308,0.6442264,0.6442264,0.64032197,0.63641757,0.6676528,0.698888,0.7262188,0.75745404,0.78868926,0.78088045,0.77307165,0.76526284,0.75745404,0.74964523,0.80040246,0.8511597,0.9019169,0.94876975,0.999527,1.1205635,1.2455044,1.3665408,1.4914817,1.6125181,1.8467822,2.077142,2.3114061,2.541766,2.77603,2.8385005,2.9048753,2.97125,3.0337205,3.1000953,3.2992198,3.49444,3.6935644,3.8887846,4.087909,3.8067923,3.521771,3.240654,2.9556324,2.6745155,3.416352,4.1581883,4.903929,5.645766,6.387602,7.57454,8.761478,9.948417,11.139259,12.326198,11.814721,11.303245,10.795672,10.284196,9.776623,11.318862,12.861101,14.40334,15.945579,17.487818,14.196406,10.901091,7.60968,4.318269,1.0268579,0.8199245,0.61689556,0.40996224,0.20693332,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.93315214,1.7413634,2.5456703,3.3538816,4.1620927,3.330455,2.4988174,1.6632754,0.8316377,0.0,0.09761006,0.19522011,0.29283017,0.39044023,0.48805028,0.9019169,1.3118792,1.7257458,2.135708,2.5495746,2.1708477,1.796025,1.4172981,1.038571,0.6637484,0.76135844,0.8589685,0.95657855,1.0541886,1.1517987,1.7101282,2.2684577,2.8306916,3.3890212,3.951255,4.5095844,5.0718184,5.630148,6.1884775,6.7507114,6.4383593,6.126007,5.813655,5.5013027,5.1889505,5.278752,5.3724575,5.466163,5.5559645,5.64967,5.251421,4.8492675,4.4510183,4.0488653,3.6506162,3.506153,3.3616903,3.213323,3.06886,2.9243972,2.8619268,2.795552,2.7291772,2.6667068,2.6003318,2.5651922,2.5300527,2.494913,2.4597735,2.4246337,2.736986,3.049338,3.3616903,3.6740425,3.9863946,3.5959544,3.2094188,2.8189783,2.4285383,2.0380979,2.4831998,2.9322062,3.3812122,3.8263142,4.2753205,4.3612175,4.4510183,4.5369153,4.6267166,4.7126136,4.5017757,4.2870336,4.0761957,3.8614538,3.6506162,3.6662338,3.6818514,3.6935644,3.7091823,3.7247996,3.6740425,3.6232853,3.5764325,3.5256753,3.474918,3.4007344,3.3265507,3.2484627,3.174279,3.1000953,2.6940374,2.2918842,1.8858263,1.4797685,1.0737107,0.9917182,0.9058213,0.8199245,0.7340276,0.6481308,0.62079996,0.59346914,0.5661383,0.5388075,0.5114767,0.74574083,0.97610056,1.2103647,1.4407244,1.6749885,1.5734742,1.475864,1.3743496,1.2767396,1.175225,1.6476578,2.1200905,2.592523,3.0649557,3.5373883,3.9863946,4.4393053,4.8883114,5.337318,5.786324,5.8644123,5.938596,6.012779,6.086963,6.1611466,6.223617,6.2860875,6.348558,6.4110284,6.473499,6.36808,6.2587566,6.153338,6.044015,5.938596,5.7980375,5.657479,5.5169206,5.376362,5.2358036,5.02887,4.8180323,4.607195,4.396357,4.1894236,4.1035266,4.0215344,3.9395418,3.8575494,3.775557,4.435401,5.095245,5.755089,6.4149327,7.0747766,6.9654536,6.8561306,6.746807,6.6335793,6.524256,6.1611466,5.801942,5.4388323,5.0757227,4.7126136,5.270943,5.8292727,6.3836975,6.942027,7.5003567,10.912805,14.325252,17.7377,21.150146,24.562595,26.190731,27.822771,29.450907,31.082947,32.711082,27.338625,21.962263,16.585901,11.213444,5.8370814,6.785851,7.7307167,8.679486,9.628256,10.573121,11.931853,13.286681,14.641508,15.996336,17.351164,17.936825,18.51858,19.10424,19.689901,20.27556,20.013966,19.748466,19.486872,19.225277,18.963682,23.4147,27.865719,32.32064,36.77166,41.22658,40.059166,38.895657,37.728237,36.564728,35.401215,33.10152,30.805735,28.50604,26.210253,23.910559,23.09454,22.278519,21.458595,20.642574,19.826555,19.639143,19.451733,19.26432,19.07691,18.885593,20.568392,22.247284,23.926178,25.608974,27.287867,27.198067,27.108265,27.018463,26.928663,26.838861,21.958359,17.08176,12.205161,7.328563,2.4480603,2.5573835,2.6667068,2.7721257,2.8814487,2.9868677,3.9161155,4.841459,5.7707067,6.6960497,7.6252975,7.570636,7.5159745,7.461313,7.406651,7.348085,9.21439,11.080693,12.946998,14.809398,16.675701,17.066143,17.460487,17.850927,18.245272,18.635712,16.527334,14.418958,12.306676,10.198298,8.086017,6.914696,5.743376,4.5681505,3.39683,2.2255092,1.8389735,1.456342,1.0698062,0.6832704,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.039044023,0.06637484,0.093705654,0.12103647,0.14836729,0.1835069,0.21864653,0.25378615,0.28892577,0.3240654,0.3435874,0.359205,0.37872702,0.39434463,0.41386664,0.48414588,0.5583295,0.62860876,0.7027924,0.77307165,0.8589685,0.94096094,1.0229534,1.1049459,1.1869383,1.1400855,1.0932326,1.0463798,0.9956226,0.94876975,0.92143893,0.8941081,0.8667773,0.8394465,0.81211567,0.8589685,0.9019169,0.94876975,0.9917182,1.038571,1.0815194,1.1205635,1.1635119,1.2064602,1.2494087,1.2494087,1.2455044,1.2415999,1.2415999,1.2376955,1.3235924,1.4133936,1.4992905,1.5890918,1.6749885,1.9443923,2.2098918,2.4792955,2.7447948,3.0141985,4.251894,5.493494,6.7311897,7.9727893,9.21439,8.449126,7.6838636,6.918601,6.153338,5.388075,4.4510183,3.5178664,2.5808098,1.6476578,0.7106012,1.4016805,2.0927596,2.7838387,3.4710135,4.1620927,3.7326086,3.3031244,2.87364,2.4441557,2.0107672,2.1981785,2.3855898,2.5769055,2.7643168,2.951728,2.8345962,2.7213683,2.6042364,2.4910088,2.3738766,2.8463092,3.3187418,3.7911747,4.263607,4.73604,4.533011,4.3260775,4.123049,3.9161155,3.7130866,6.083059,8.453031,10.823003,13.192975,15.562947,14.2666855,12.974329,11.678067,10.381805,9.089449,8.36323,7.6409154,6.918601,6.196286,5.473972,4.7126136,3.951255,3.1859922,2.4246337,1.6632754,1.3314011,0.9956226,0.6637484,0.3318742,0.0,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,0.64032197,0.6559396,0.6715572,0.6832704,0.698888,0.63251317,0.5661383,0.4958591,0.42948425,0.3631094,0.28892577,0.21864653,0.14446288,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.45291066,0.8784905,1.3079748,1.7335546,2.1630387,2.5378613,2.912684,3.2875066,3.6623292,4.037152,4.337791,4.6384296,4.939069,5.2358036,5.5364423,5.493494,5.45445,5.4115014,5.368553,5.3256044,5.083532,4.845363,4.60329,4.365122,4.123049,4.0527697,3.978586,3.9083066,3.8341231,3.7638438,4.193328,4.6267166,5.0601053,5.493494,5.9268827,5.3138914,4.704805,4.095718,3.4866312,2.87364,2.6549935,2.436347,2.2137961,1.9951496,1.7765031,2.8658314,3.959064,5.0522966,6.1455293,7.238762,6.89127,6.547683,6.2040954,5.8566036,5.5130157,5.4856853,5.4583545,5.4310236,5.4036927,5.376362,5.2045684,5.036679,4.8648853,4.6930914,4.5252023,4.9781127,5.4310236,5.883934,6.336845,6.785851,6.461786,6.13772,5.813655,5.4856853,5.1616197,5.7199492,6.278279,6.8366084,7.3910336,7.9493628,7.558923,7.164578,6.774138,6.379793,5.989353,5.2553253,4.521298,3.7911747,3.057147,2.3231194,2.3933985,2.463678,2.533957,2.6042364,2.6745155,2.5027218,2.330928,2.1591344,1.9834363,1.8116426,1.7413634,1.6671798,1.5969005,1.5227169,1.4485333,1.33921,1.2259823,1.1127546,0.999527,0.8862993,1.261122,1.6359446,2.0107672,2.3855898,2.7643168,2.5690966,2.3738766,2.1786566,1.9834363,1.7882162,2.533957,3.2836022,4.029343,4.7789884,5.5247293,6.2040954,6.8795567,7.558923,8.234385,8.913751,0.6754616,0.6715572,0.6637484,0.659844,0.6559396,0.6481308,0.6715572,0.6949836,0.71841,0.7418364,0.76135844,0.76135844,0.75745404,0.75354964,0.75354964,0.74964523,0.80040246,0.8511597,0.9019169,0.94876975,0.999527,1.1088502,1.2142692,1.3235924,1.4290112,1.5383345,1.7257458,1.9170616,2.1083772,2.2957885,2.4871042,2.6042364,2.7213683,2.8385005,2.9556324,3.076669,3.39683,3.7130866,4.0332475,4.3534083,4.6735697,4.40807,4.1464753,3.8809757,3.6154766,3.349977,3.970777,4.5954814,5.2162814,5.840986,6.461786,7.699481,8.937177,10.174872,11.412568,12.650263,12.205161,11.760059,11.314958,10.869856,10.424754,11.623405,12.818152,14.016804,15.215456,16.414106,13.376482,10.342762,7.309041,4.271416,1.2376955,0.9917182,0.7418364,0.4958591,0.24597734,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.76526284,1.4055848,2.0459068,2.6862288,3.3265507,2.6588979,1.9951496,1.3314011,0.6637484,0.0,0.13274968,0.26549935,0.39824903,0.5309987,0.6637484,1.0737107,1.4875772,1.901444,2.3114061,2.7252727,2.4090161,2.0888553,1.7725986,1.456342,1.1361811,1.358732,1.5773785,1.796025,2.018576,2.2372224,2.7682211,3.3031244,3.8341231,4.369026,4.900025,5.2436123,5.591104,5.9346914,6.278279,6.6257706,6.699954,6.774138,6.8483214,6.9264097,7.000593,7.1333427,7.269997,7.406651,7.5394006,7.676055,7.223144,6.774138,6.3251314,5.8761253,5.423215,5.0483923,4.6696653,4.290938,3.9161155,3.5373883,3.4202564,3.3031244,3.1859922,3.06886,2.951728,2.9283018,2.9087796,2.8892577,2.8697357,2.8502135,3.1508527,3.4514916,3.7482262,4.0488653,4.349504,3.959064,3.5647192,3.174279,2.7799344,2.3855898,2.9087796,3.4280653,3.9473507,4.466636,4.985922,4.911738,4.8375545,4.7633705,4.689187,4.6110992,4.4861584,4.3612175,4.2362766,4.1113358,3.9863946,4.041056,4.095718,4.154284,4.2089458,4.263607,4.0996222,3.9356375,3.775557,3.611572,3.4514916,3.338264,3.2250361,3.1118085,2.998581,2.8892577,2.5534792,2.2177005,1.8819219,1.5461433,1.2142692,1.2298868,1.2494087,1.2650263,1.2806439,1.3001659,1.183034,1.0659018,0.94876975,0.8316377,0.7106012,0.94096094,1.1674163,1.3938715,1.6242313,1.8506867,1.737459,1.6242313,1.5110037,1.4016805,1.2884527,1.6437533,2.0029583,2.358259,2.717464,3.076669,3.4632049,3.8497405,4.2362766,4.6267166,5.0132523,5.1108627,5.212377,5.3138914,5.4115014,5.5130157,5.575486,5.6379566,5.700427,5.7628975,5.825368,5.833177,5.84489,5.8566036,5.8644123,5.8761253,5.9073606,5.938596,5.9737353,6.0049706,6.036206,5.7785153,5.520825,5.263134,5.009348,4.7516575,4.560342,4.369026,4.181615,3.9902992,3.7989833,4.40807,5.0132523,5.6223392,6.2314262,6.8366084,6.7311897,6.621866,6.5164475,6.407124,6.3017054,5.9737353,5.64967,5.3256044,5.001539,4.6735697,5.388075,6.1064854,6.8209906,7.535496,8.250002,10.760532,13.274967,15.789403,18.299932,20.81437,23.047686,25.281004,27.518227,29.751545,31.988768,26.77639,21.564014,16.351637,11.139259,5.9268827,7.043542,8.164105,9.284669,10.405232,11.525795,13.396004,15.270117,17.14423,19.014439,20.888552,21.958359,23.028164,24.097971,25.167776,26.237583,25.101402,23.961317,22.825136,21.688955,20.548868,23.805141,27.061413,30.31378,33.57005,36.82632,36.85756,36.888794,36.92393,36.955166,36.986404,34.604717,32.22303,29.841347,27.455757,25.074072,24.23853,23.40689,22.57135,21.735807,20.900265,20.67381,20.45126,20.224804,19.998348,19.775797,21.13453,22.493261,23.855898,25.21463,26.573362,26.182922,25.788576,25.398136,25.003792,24.613352,20.431738,16.254026,12.072412,7.890797,3.7130866,3.4514916,3.193801,2.9322062,2.6706111,2.4129205,3.1430438,3.873167,4.60329,5.3334136,6.0635366,6.2275214,6.3915067,6.559396,6.7233806,6.8873653,8.59359,10.295909,12.002132,13.708356,15.410676,15.883108,16.355541,16.831879,17.30431,17.776743,15.719124,13.661504,11.603884,9.546264,7.4886436,6.329036,5.173333,4.0137253,2.8580225,1.698415,1.4055848,1.1088502,0.8160201,0.5192855,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.05466163,0.08589685,0.113227665,0.14446288,0.1756981,0.20693332,0.23816854,0.27330816,0.30454338,0.3357786,0.359205,0.38263142,0.40605783,0.42557985,0.44900626,0.5700427,0.6910792,0.80821127,0.92924774,1.0502841,1.2142692,1.3782539,1.5461433,1.7101282,1.8741131,1.7804074,1.6867018,1.5890918,1.4953861,1.4016805,1.3431144,1.2884527,1.2337911,1.1791295,1.1244678,1.2259823,1.3314011,1.4329157,1.53443,1.6359446,1.7843118,1.9326792,2.0810463,2.2294137,2.3738766,2.3699722,2.366068,2.358259,2.3543546,2.35045,2.4871042,2.6237583,2.7643168,2.900971,3.0376248,3.4983444,3.959064,4.415879,4.8765984,5.337318,6.2314262,7.1216297,8.015738,8.905942,9.80005,9.99527,10.19049,10.38571,10.58093,10.77615,8.730244,6.6843367,4.6384296,2.5964274,0.5505207,1.1791295,1.8116426,2.4402514,3.06886,3.7013733,3.3655949,3.0298162,2.6940374,2.358259,2.0263848,2.338737,2.6510892,2.9634414,3.2757936,3.5881457,3.6467118,3.7013733,3.7599394,3.8185053,3.873167,4.369026,4.8648853,5.3607445,5.8566036,6.348558,6.1884775,6.028397,5.8683167,5.708236,5.548156,8.226576,10.904996,13.583415,16.261835,18.936352,17.323833,15.70741,14.090988,12.47847,10.862047,10.592644,10.323239,10.053836,9.784432,9.511124,8.136774,6.7624245,5.388075,4.0137253,2.639376,2.1083772,1.5812829,1.0541886,0.5270943,0.0,0.24988174,0.4997635,0.74964523,0.999527,1.2494087,1.2806439,1.3118792,1.33921,1.3704453,1.4016805,1.2650263,1.1283722,0.9956226,0.8589685,0.7262188,0.58175594,0.43338865,0.28892577,0.14446288,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.37872702,0.7106012,1.038571,1.3704453,1.698415,2.0263848,2.35045,2.6745155,2.998581,3.3265507,3.736513,4.1503797,4.564246,4.9742084,5.388075,5.563773,5.743376,5.919074,6.098676,6.2743745,5.833177,5.388075,4.9468775,4.50568,4.0605783,4.267512,4.474445,4.677474,4.884407,5.087436,5.579391,6.067441,6.559396,7.0474463,7.5394006,6.578918,5.6223392,4.6657605,3.7091823,2.7486992,2.4831998,2.2216048,1.9561055,1.6906061,1.4251068,2.3465457,3.2718892,4.193328,5.114767,6.036206,5.8097506,5.5832953,5.35684,5.12648,4.900025,4.958591,5.0132523,5.0718184,5.1303844,5.1889505,5.1460023,5.1069584,5.067914,5.02887,4.985922,5.368553,5.74728,6.126007,6.5086384,6.8873653,6.801469,6.7116675,6.6257706,6.5359693,6.4500723,7.1294384,7.8049,8.484266,9.159728,9.839094,9.190963,8.542832,7.8947015,7.2465706,6.5984397,5.872221,5.1460023,4.415879,3.68966,2.9634414,3.0532427,3.1430438,3.232845,3.3226464,3.4124475,3.1781836,2.9478238,2.7135596,2.4831998,2.2489357,2.0927596,1.9365835,1.7765031,1.620327,1.4641509,1.3626363,1.261122,1.1635119,1.0619974,0.96438736,1.261122,1.5617609,1.8623998,2.1630387,2.463678,2.2840753,2.1083772,1.9287747,1.7530766,1.5734742,2.3816853,3.1898966,3.998108,4.806319,5.610626,6.2548523,6.899079,7.5394006,8.183627,8.823949,0.698888,0.6910792,0.6832704,0.679366,0.6715572,0.6637484,0.679366,0.6910792,0.7066968,0.7223144,0.737932,0.7418364,0.7418364,0.74574083,0.74574083,0.74964523,0.80040246,0.8511597,0.9019169,0.94876975,0.999527,1.0932326,1.1869383,1.2767396,1.3704453,1.4641509,1.6086137,1.756981,1.9053483,2.0537157,2.1981785,2.3699722,2.541766,2.7096553,2.8814487,3.049338,3.49444,3.9356375,4.376835,4.8219366,5.263134,5.0132523,4.7672753,4.521298,4.271416,4.025439,4.5291066,5.02887,5.532538,6.036206,6.5359693,7.824422,9.112875,10.401327,11.685876,12.974329,12.595602,12.216875,11.834243,11.455516,11.076789,11.927949,12.779109,13.634172,14.4853325,15.336493,12.560462,9.784432,7.0044975,4.2284675,1.4485333,1.1596074,0.8706817,0.58175594,0.28892577,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.59737355,1.0698062,1.542239,2.0146716,2.4871042,1.9912452,1.4914817,0.9956226,0.4958591,0.0,0.1678893,0.3357786,0.5036679,0.6715572,0.8394465,1.2494087,1.6632754,2.0732377,2.4871042,2.900971,2.6432803,2.3855898,2.1278992,1.8702087,1.6125181,1.9561055,2.2957885,2.639376,2.9829633,3.3265507,3.8302186,4.3338866,4.841459,5.3451266,5.8487945,5.9815445,6.1103897,6.239235,6.36808,6.5008297,6.9615493,7.426173,7.8868923,8.351517,8.812236,8.991838,9.167537,9.343235,9.522837,9.698535,9.198771,8.699008,8.1992445,7.699481,7.1997175,6.590631,5.9815445,5.368553,4.759466,4.1503797,3.978586,3.8106966,3.638903,3.4710135,3.2992198,3.2953155,3.2914112,3.2836022,3.279698,3.2757936,3.5608149,3.8497405,4.138666,4.423688,4.7126136,4.318269,3.9239242,3.5256753,3.1313305,2.736986,3.330455,3.9239242,4.513489,5.1069584,5.700427,5.462259,5.22409,4.985922,4.7516575,4.513489,4.474445,4.4393053,4.4002614,4.3612175,4.3260775,4.4197836,4.513489,4.6110992,4.704805,4.7985106,4.5252023,4.251894,3.9746814,3.7013733,3.4241607,3.2757936,3.1235218,2.9751544,2.8267872,2.6745155,2.4090161,2.1435168,1.8819219,1.6164225,1.3509232,1.4680552,1.5890918,1.7101282,1.8311646,1.9482968,1.7413634,1.53443,1.3274968,1.1205635,0.9136301,1.1361811,1.358732,1.5812829,1.8038338,2.0263848,1.901444,1.7765031,1.6515622,1.5266213,1.4016805,1.6437533,1.8858263,2.1278992,2.3699722,2.612045,2.9361105,3.2640803,3.5881457,3.912211,4.2362766,4.3612175,4.4861584,4.6110992,4.73604,4.860981,4.9234514,4.985922,5.0483923,5.1108627,5.173333,5.3021784,5.4310236,5.5559645,5.6848097,5.813655,6.016684,6.223617,6.426646,6.6335793,6.8366084,6.532065,6.2275214,5.9229784,5.618435,5.3138914,5.0132523,4.716518,4.4197836,4.123049,3.8263142,4.380739,4.9351645,5.4895897,6.044015,6.5984397,6.4969254,6.3915067,6.2860875,6.180669,6.0752497,5.786324,5.5013027,5.212377,4.9234514,4.6384296,5.5091114,6.3836975,7.2543793,8.128965,8.999647,10.612165,12.224684,13.837202,15.449719,17.062239,19.900738,22.743143,25.581644,28.42405,31.262548,26.214157,21.16186,16.113468,11.061172,6.012779,7.3051367,8.597494,9.889851,11.182208,12.4745655,14.864059,17.253553,19.646952,22.036446,24.425941,25.979893,27.533844,29.091702,30.645653,32.199604,30.188839,28.174168,26.163399,24.148727,22.13796,24.195581,26.2532,28.310822,30.36844,32.42606,33.65595,34.885834,36.115723,37.345608,38.575493,36.10791,33.64033,31.172749,28.705166,26.237583,25.386423,24.531359,23.6802,22.82904,21.973976,21.712381,21.450787,21.189192,20.92369,20.662096,21.700668,22.743143,23.781713,24.82419,25.86276,25.167776,24.472794,23.77781,23.082827,22.387842,18.905115,15.422389,11.939662,8.456935,4.9742084,4.3455997,3.7208953,3.0922866,2.463678,1.8389735,2.3699722,2.900971,3.435874,3.9668727,4.5017757,4.884407,5.270943,5.6535745,6.04011,6.426646,7.968885,9.515028,11.061172,12.603411,14.149553,14.703979,15.254499,15.808925,16.359446,16.91387,14.907008,12.90405,10.897186,8.894228,6.8873653,5.743376,4.60329,3.4593005,2.3192148,1.175225,0.96829176,0.76526284,0.5583295,0.3553006,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.07027924,0.10151446,0.13665408,0.1678893,0.19912452,0.23035973,0.26159495,0.28892577,0.32016098,0.3513962,0.37872702,0.40605783,0.43338865,0.46071947,0.48805028,0.6559396,0.8238289,0.9917182,1.1557031,1.3235924,1.5734742,1.8194515,2.069333,2.3153105,2.5612879,2.4207294,2.2762666,2.135708,1.9912452,1.8506867,1.7686942,1.6867018,1.6008049,1.5188124,1.43682,1.5969005,1.756981,1.9170616,2.077142,2.2372224,2.4910088,2.7408905,2.9946766,3.2484627,3.4983444,3.49444,3.4866312,3.4788225,3.4710135,3.4632049,3.6506162,3.8380275,4.025439,4.21285,4.4002614,5.0522966,5.704332,6.356367,7.008402,7.6643414,8.207053,8.75367,9.296382,9.8429985,10.38571,11.541413,12.697116,13.852819,15.008522,16.164225,13.005564,9.850807,6.6960497,3.541293,0.38653582,0.95657855,1.5266213,2.096664,2.6667068,3.2367494,2.998581,2.7565079,2.5183394,2.2762666,2.0380979,2.475391,2.912684,3.349977,3.78727,4.224563,4.454923,4.6852827,4.9156423,5.1460023,5.376362,5.891743,6.4110284,6.9264097,7.445695,7.9610763,7.8478484,7.7307167,7.617489,7.504261,7.387129,10.373997,13.35696,16.343828,19.326792,22.31366,20.377075,18.444397,16.507812,14.571229,12.63855,12.818152,13.001659,13.185166,13.368673,13.548276,11.560935,9.573594,7.5862536,5.5989127,3.611572,2.8892577,2.1669433,1.4446288,0.7223144,0.0,0.37482262,0.74964523,1.1244678,1.4992905,1.8741131,1.9209659,1.9639144,2.0107672,2.0537157,2.1005683,1.8975395,1.6945106,1.4914817,1.2884527,1.0893283,0.8706817,0.6520352,0.43338865,0.21864653,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.30844778,0.5388075,0.77307165,1.0034313,1.2376955,1.5110037,1.7882162,2.0615244,2.338737,2.612045,3.1391394,3.6623292,4.1894236,4.7126136,5.2358036,5.6340523,6.0323014,6.4305506,6.8287997,7.223144,6.578918,5.9346914,5.290465,4.646239,3.998108,4.482254,4.9663997,5.446641,5.930787,6.4110284,6.9615493,7.5081654,8.054782,8.601398,9.151918,7.843944,6.5398736,5.2358036,3.9317331,2.6237583,2.3153105,2.0068626,1.6945106,1.3860629,1.0737107,1.8272603,2.5808098,3.3343596,4.084005,4.8375545,4.728231,4.618908,4.50568,4.396357,4.2870336,4.4314966,4.572055,4.716518,4.8570766,5.001539,5.0913405,5.181142,5.270943,5.3607445,5.4505453,5.758993,6.0635366,6.3719845,6.6804323,6.98888,7.137247,7.2856145,7.437886,7.5862536,7.7385254,8.535024,9.331521,10.131924,10.928422,11.72492,10.823003,9.921086,9.019169,8.113348,7.211431,6.4891167,5.7668023,5.044488,4.322173,3.5998588,3.7091823,3.8185053,3.9317331,4.041056,4.1503797,3.8575494,3.5647192,3.2718892,2.979059,2.6862288,2.4441557,2.2020829,1.9600099,1.717937,1.475864,1.3860629,1.3001659,1.2142692,1.1244678,1.038571,1.261122,1.4875772,1.7140326,1.9365835,2.1630387,2.0029583,1.8428779,1.6827974,1.5227169,1.3626363,2.2294137,3.096191,3.9668727,4.83365,5.700427,6.3056097,6.914696,7.523783,8.128965,8.738052,0.7262188,0.7145056,0.7066968,0.6949836,0.6832704,0.6754616,0.6832704,0.6910792,0.698888,0.7066968,0.7106012,0.71841,0.7262188,0.7340276,0.7418364,0.74964523,0.80040246,0.8511597,0.9019169,0.94876975,0.999527,1.077615,1.1557031,1.2337911,1.3118792,1.3860629,1.4914817,1.5969005,1.7023194,1.8077383,1.9131571,2.135708,2.358259,2.5808098,2.803361,3.0259118,3.5881457,4.154284,4.7204223,5.2865605,5.8487945,5.618435,5.388075,5.1616197,4.93126,4.7009,5.083532,5.466163,5.8487945,6.2314262,6.6140575,7.9493628,9.288573,10.6238785,11.963089,13.298394,12.986042,12.6697855,12.353529,12.041177,11.72492,12.232492,12.740065,13.247637,13.755209,14.262781,11.744442,9.2221985,6.703859,4.181615,1.6632754,1.3314011,0.9956226,0.6637484,0.3318742,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.42948425,0.7340276,1.038571,1.3431144,1.6515622,1.319688,0.9917182,0.659844,0.3318742,0.0,0.20302892,0.40605783,0.60908675,0.80821127,1.0112402,1.4251068,1.8389735,2.2489357,2.6628022,3.076669,2.8775444,2.67842,2.4831998,2.2840753,2.0888553,2.5534792,3.018103,3.4827268,3.9473507,4.4119744,4.8883114,5.368553,5.84489,6.321227,6.801469,6.715572,6.629675,6.5437784,6.461786,6.375889,7.223144,8.074304,8.925464,9.776623,10.6238785,10.84643,11.065076,11.283723,11.506273,11.72492,11.174399,10.6238785,10.073358,9.526741,8.976221,8.13287,7.289519,6.446168,5.606722,4.7633705,4.5408196,4.318269,4.095718,3.873167,3.6506162,3.6584249,3.6701381,3.6818514,3.68966,3.7013733,3.9746814,4.251894,4.5252023,4.7985106,5.0757227,4.677474,4.279225,3.8809757,3.4866312,3.0883822,3.7521305,4.415879,5.083532,5.74728,6.4110284,6.012779,5.610626,5.212377,4.814128,4.4119744,4.462732,4.513489,4.564246,4.6110992,4.661856,4.7985106,4.93126,5.067914,5.2006636,5.337318,4.950782,4.564246,4.173806,3.78727,3.4007344,3.213323,3.0259118,2.8385005,2.6510892,2.463678,2.2684577,2.0732377,1.8780174,1.6827974,1.4875772,1.7101282,1.9326792,2.15523,2.377781,2.6003318,2.3035975,2.0068626,1.7062237,1.4094892,1.1127546,1.3314011,1.5461433,1.7647898,1.9834363,2.1981785,2.0615244,1.9248703,1.7882162,1.6515622,1.5110037,1.639849,1.7686942,1.893635,2.0224805,2.1513257,2.4129205,2.6745155,2.9361105,3.2016098,3.4632049,3.611572,3.7638438,3.912211,4.0605783,4.21285,4.2753205,4.337791,4.4002614,4.462732,4.5252023,4.7711797,5.0132523,5.2592297,5.505207,5.7511845,6.126007,6.504734,6.883461,7.2582836,7.6370106,7.2856145,6.9342184,6.578918,6.2275214,5.8761253,5.4700675,5.0640097,4.661856,4.2557983,3.8497405,4.3534083,4.853172,5.35684,5.860508,6.364176,6.2587566,6.1572423,6.055728,5.9542136,5.8487945,5.5989127,5.349031,5.099149,4.8492675,4.5993857,5.630148,6.66091,7.6916723,8.718531,9.749292,10.4637985,11.174399,11.888905,12.599506,13.314012,16.757694,20.201378,23.648964,27.092648,30.53633,25.651922,20.76361,15.875299,10.986988,6.098676,7.5667315,9.030883,10.495033,11.959184,13.423335,16.332115,19.240894,22.14577,25.05455,27.96333,30.001427,32.04343,34.081528,36.12353,38.16163,35.276276,32.387016,29.501663,26.612406,23.723148,24.586021,25.44499,26.303959,27.16683,28.025799,30.454338,32.87897,35.30751,37.73605,40.160683,37.611107,35.05763,32.50415,29.95067,27.401094,26.530413,25.65973,24.78905,23.918367,23.05159,22.750952,22.450314,22.149673,21.849035,21.548395,22.27071,22.98912,23.711435,24.429846,25.148254,24.152632,23.153105,22.157482,21.16186,20.162333,17.378494,14.590752,11.806912,9.023073,6.239235,5.2436123,4.2479897,3.252367,2.2567444,1.261122,1.5969005,1.9326792,2.2684577,2.6042364,2.9361105,3.541293,4.1464753,4.7516575,5.35684,5.9620223,7.348085,8.734148,10.116306,11.502369,12.888432,13.520945,14.153459,14.785972,15.418485,16.050997,14.098797,12.146595,10.19049,8.238289,6.2860875,5.1616197,4.0332475,2.9048753,1.7765031,0.6481308,0.5349031,0.42167544,0.30454338,0.19131571,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.08589685,0.12103647,0.15617609,0.19131571,0.22645533,0.25378615,0.28111696,0.30844778,0.3357786,0.3631094,0.39434463,0.42557985,0.46071947,0.49195468,0.5231899,0.7418364,0.95657855,1.1713207,1.3860629,1.6008049,1.9287747,2.260649,2.5886188,2.920493,3.2484627,3.0610514,2.8697357,2.67842,2.4910088,2.2996929,2.1903696,2.0810463,1.9717231,1.8584955,1.7491722,1.9678187,2.1864653,2.4012074,2.619854,2.8385005,3.193801,3.5530062,3.9083066,4.267512,4.6267166,4.6150036,4.60329,4.5954814,4.5837684,4.575959,4.814128,5.0483923,5.2865605,5.5247293,5.7628975,6.606249,7.453504,8.296855,9.14411,9.987461,10.186585,10.381805,10.58093,10.77615,10.975275,13.091461,15.203742,17.31993,19.436115,21.548395,17.284788,13.021181,8.75367,4.4900627,0.22645533,0.7340276,1.2455044,1.7530766,2.2645533,2.77603,2.631567,2.4831998,2.338737,2.194274,2.0498111,2.612045,3.174279,3.736513,4.298747,4.860981,5.263134,5.6691923,6.0713453,6.473499,6.8756523,7.4144597,7.9532676,8.495979,9.034787,9.573594,9.503315,9.43694,9.366661,9.296382,9.226103,12.517513,15.808925,19.10424,22.39565,25.687063,23.434223,21.177479,18.920732,16.667892,14.411149,15.047566,15.683984,16.316498,16.952915,17.589333,14.989,12.388668,9.788337,7.1880045,4.5876727,3.6701381,2.7526035,1.8350691,0.91753453,0.0,0.4997635,0.999527,1.4992905,1.999054,2.4988174,2.5612879,2.619854,2.67842,2.7408905,2.7994564,2.5300527,2.260649,1.9912452,1.7218413,1.4485333,1.1596074,0.8706817,0.58175594,0.28892577,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.23426414,0.3709182,0.5036679,0.64032197,0.77307165,0.999527,1.2259823,1.4485333,1.6749885,1.901444,2.5378613,3.174279,3.8106966,4.4510183,5.087436,5.704332,6.321227,6.9381227,7.558923,8.175818,7.328563,6.481308,5.6340523,4.786797,3.9356375,4.6969957,5.4583545,6.2158084,6.9771667,7.7385254,8.343708,8.94889,9.554072,10.159255,10.764437,9.108971,7.4574084,5.805846,4.154284,2.4988174,2.1435168,1.7882162,1.43682,1.0815194,0.7262188,1.3079748,1.8897307,2.4714866,3.0532427,3.638903,3.6467118,3.6506162,3.6584249,3.6662338,3.6740425,3.9044023,4.1308575,4.357313,4.5837684,4.814128,5.0327744,5.251421,5.473972,5.6926184,5.911265,6.1494336,6.3836975,6.617962,6.852226,7.08649,7.47693,7.8634663,8.250002,8.636538,9.023073,9.944512,10.862047,11.775677,12.693212,13.610746,12.455043,11.295436,10.139732,8.98403,7.824422,7.1060123,6.3915067,5.6730967,4.9546866,4.2362766,4.369026,4.4978714,4.6267166,4.755562,4.8883114,4.5369153,4.181615,3.8302186,3.4788225,3.1235218,2.795552,2.4714866,2.1435168,1.815547,1.4875772,1.4133936,1.33921,1.261122,1.1869383,1.1127546,1.261122,1.4133936,1.5617609,1.7140326,1.8623998,1.7218413,1.5773785,1.43682,1.2923572,1.1517987,2.077142,3.0063896,3.9317331,4.860981,5.786324,6.3602715,6.9342184,7.504261,8.078208,8.648251,0.74964523,0.737932,0.7262188,0.7106012,0.698888,0.6871748,0.6871748,0.6871748,0.6871748,0.6871748,0.6871748,0.698888,0.7106012,0.7262188,0.737932,0.74964523,0.80040246,0.8511597,0.9019169,0.94876975,0.999527,1.0619974,1.1244678,1.1869383,1.2494087,1.3118792,1.3743496,1.43682,1.4992905,1.5617609,1.6242313,1.901444,2.174752,2.4480603,2.7252727,2.998581,3.6857557,4.376835,5.0640097,5.7511845,6.4383593,6.223617,6.012779,5.801942,5.5871997,5.376362,5.6379566,5.899552,6.1611466,6.426646,6.688241,8.074304,9.464272,10.850334,12.236397,13.626364,13.376482,13.1266,12.8767185,12.626837,12.373051,12.537036,12.70102,12.861101,13.025085,13.189071,10.924518,8.663869,6.3993154,4.138666,1.8741131,1.4992905,1.1244678,0.74964523,0.37482262,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.26159495,0.39824903,0.5388075,0.6754616,0.81211567,0.6481308,0.48805028,0.3240654,0.1639849,0.0,0.23816854,0.47633708,0.7106012,0.94876975,1.1869383,1.6008049,2.0107672,2.4246337,2.8385005,3.2484627,3.1118085,2.9751544,2.8385005,2.7018464,2.5612879,3.1508527,3.736513,4.3260775,4.911738,5.5013027,5.950309,6.3993154,6.8483214,7.3012323,7.7502384,7.4495993,7.1489606,6.8483214,6.551587,6.250948,7.4886436,8.726339,9.964035,11.20173,12.439425,12.70102,12.962616,13.224211,13.4858055,13.751305,13.150026,12.548749,11.951375,11.350098,10.748819,9.675109,8.601398,7.523783,6.4500723,5.376362,5.099149,4.825841,4.548629,4.2753205,3.998108,4.025439,4.0488653,4.0761957,4.0996222,4.123049,4.388548,4.650143,4.911738,5.173333,5.4388323,5.036679,4.6384296,4.2362766,3.8380275,3.435874,4.173806,4.911738,5.64967,6.387602,7.125534,6.5633,6.001066,5.4388323,4.8765984,4.3143644,4.4510183,4.5876727,4.7243266,4.860981,5.001539,5.173333,5.349031,5.5247293,5.700427,5.8761253,5.376362,4.8765984,4.376835,3.873167,3.3734035,3.1508527,2.9243972,2.7018464,2.475391,2.2489357,2.1239948,1.999054,1.8741131,1.7491722,1.6242313,1.9482968,2.2762666,2.6003318,2.9243972,3.2484627,2.8619268,2.475391,2.0888553,1.698415,1.3118792,1.5266213,1.737459,1.9482968,2.1630387,2.3738766,2.2255092,2.0732377,1.9248703,1.7765031,1.6242313,1.6359446,1.6515622,1.6632754,1.6749885,1.6867018,1.8858263,2.0888553,2.2879796,2.4871042,2.6862288,2.8619268,3.0376248,3.213323,3.3890212,3.5608149,3.6232853,3.6857557,3.7482262,3.8106966,3.873167,4.2362766,4.5993857,4.9624953,5.3256044,5.688714,6.239235,6.785851,7.336372,7.8868923,8.437413,8.039165,7.6370106,7.238762,6.8366084,6.4383593,5.9268827,5.4115014,4.900025,4.388548,3.873167,4.3260775,4.775084,5.22409,5.6730967,6.126007,6.0244927,5.9268827,5.825368,5.7238536,5.6262436,5.4115014,5.2006636,4.985922,4.775084,4.564246,5.7511845,6.9381227,8.125061,9.311999,10.498938,10.311526,10.124115,9.936704,9.749292,9.561881,13.610746,17.663515,21.712381,25.761246,29.814016,25.085785,20.361458,15.637131,10.912805,6.1884775,7.824422,9.464272,11.100216,12.73616,14.376009,17.800169,21.22433,24.64849,28.076557,31.500717,34.026867,36.54911,39.075256,41.601406,44.12365,40.363712,36.599865,32.83602,29.076084,25.31224,24.976461,24.636778,24.300999,23.961317,23.625538,27.248823,30.876013,34.4993,38.126488,41.749775,39.110397,36.474926,33.83555,31.200079,28.560703,27.674404,26.788103,25.901804,25.0116,24.125301,23.785618,23.44984,23.114061,22.774378,22.4386,22.83685,23.239002,23.63725,24.039404,24.437654,23.137487,21.837322,20.537155,19.23699,17.936825,15.847969,13.763018,11.674163,9.589212,7.5003567,6.13772,4.775084,3.4124475,2.0498111,0.6871748,0.8238289,0.96438736,1.1010414,1.2376955,1.3743496,2.1981785,3.0259118,3.8497405,4.6735697,5.5013027,6.7233806,7.9493628,9.175345,10.401327,11.623405,12.337912,13.048512,13.763018,14.473619,15.188125,13.286681,11.389141,9.487698,7.5862536,5.688714,4.575959,3.4632049,2.35045,1.2376955,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.10151446,0.13665408,0.1756981,0.21083772,0.24988174,0.27330816,0.30063897,0.3240654,0.3513962,0.37482262,0.41386664,0.44900626,0.48805028,0.5231899,0.5622339,0.8238289,1.0893283,1.3509232,1.6125181,1.8741131,2.2879796,2.7018464,3.1118085,3.5256753,3.9356375,3.7013733,3.4632049,3.2250361,2.9868677,2.7486992,2.612045,2.475391,2.338737,2.1981785,2.0615244,2.338737,2.612045,2.8892577,3.1625657,3.435874,3.900498,4.3612175,4.825841,5.2865605,5.7511845,5.735567,5.7238536,5.7121406,5.700427,5.688714,5.9737353,6.262661,6.551587,6.8366084,7.125534,8.164105,9.198771,10.237343,11.275913,12.31058,12.162213,12.013845,11.861574,11.713207,11.560935,14.637604,17.714273,20.787037,23.863707,26.936472,21.564014,16.187653,10.81129,5.4388323,0.062470436,0.5114767,0.96438736,1.4133936,1.8623998,2.3114061,2.260649,2.2137961,2.1630387,2.1122816,2.0615244,2.7486992,3.435874,4.126953,4.814128,5.5013027,6.0752497,6.649197,7.223144,7.800996,8.374943,8.937177,9.499411,10.061645,10.6238785,11.186112,11.162686,11.139259,11.111929,11.088503,11.061172,14.661031,18.26089,21.860748,25.460608,29.064371,26.487465,23.914463,21.337559,18.760653,16.187653,17.27698,18.362404,19.451733,20.537155,21.626484,18.41316,15.199838,11.986515,8.773191,5.563773,4.4510183,3.338264,2.2255092,1.1127546,0.0,0.62470436,1.2494087,1.8741131,2.4988174,3.1235218,3.2016098,3.2757936,3.349977,3.4241607,3.4983444,3.1625657,2.8267872,2.4871042,2.1513257,1.8116426,1.4485333,1.0893283,0.7262188,0.3631094,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.1639849,0.19912452,0.23816854,0.27330816,0.31235218,0.48805028,0.6637484,0.8394465,1.0112402,1.1869383,1.9365835,2.6862288,3.435874,4.185519,4.939069,5.774611,6.6140575,7.4495993,8.289046,9.124588,8.074304,7.0240197,5.9737353,4.9234514,3.873167,4.911738,5.950309,6.98888,8.023546,9.062118,9.725866,10.38571,11.0494585,11.713207,12.373051,10.373997,8.374943,6.375889,4.376835,2.3738766,1.9756275,1.5734742,1.175225,0.77697605,0.37482262,0.78868926,1.1986516,1.6125181,2.0263848,2.436347,2.5612879,2.6862288,2.8111696,2.9361105,3.0610514,3.3734035,3.6857557,3.998108,4.3143644,4.6267166,4.9742084,5.3256044,5.6730967,6.0244927,6.375889,6.5359693,6.699954,6.8639393,7.0240197,7.1880045,7.812709,8.437413,9.062118,9.686822,10.311526,11.350098,12.388668,13.423335,14.461906,15.500477,14.087084,12.67369,11.2642,9.850807,8.437413,7.726812,7.012306,6.3017054,5.5871997,4.8765984,5.024966,5.173333,5.3256044,5.473972,5.6262436,5.212377,4.7985106,4.388548,3.9746814,3.5608149,3.1508527,2.736986,2.3231194,1.9131571,1.4992905,1.43682,1.3743496,1.3118792,1.2494087,1.1869383,1.261122,1.33921,1.4133936,1.4875772,1.5617609,1.43682,1.3118792,1.1869383,1.0619974,0.93705654,1.9248703,2.912684,3.900498,4.8883114,5.8761253,6.4110284,6.949836,7.4886436,8.023546,8.562354,0.737932,0.7262188,0.7106012,0.698888,0.6871748,0.6754616,0.679366,0.679366,0.6832704,0.6832704,0.6871748,0.7027924,0.71841,0.7340276,0.74574083,0.76135844,0.80821127,0.8511597,0.8980125,0.94096094,0.9878138,1.0463798,1.1088502,1.1674163,1.2259823,1.2884527,1.3860629,1.4875772,1.5890918,1.6867018,1.7882162,2.1630387,2.5378613,2.912684,3.2875066,3.6623292,4.173806,4.6813784,5.192855,5.704332,6.211904,6.098676,5.989353,5.8761253,5.7628975,5.64967,5.903456,6.1611466,6.4149327,6.6687193,6.9264097,8.39056,9.854712,11.318862,12.786918,14.251068,13.895767,13.544372,13.192975,12.841579,12.486279,12.96652,13.442857,13.919194,14.399435,14.875772,12.24811,9.6243515,7.000593,4.376835,1.7491722,1.4055848,1.0580931,0.7145056,0.3709182,0.023426414,0.039044023,0.05466163,0.07027924,0.08589685,0.10151446,0.22645533,0.3513962,0.47633708,0.60127795,0.7262188,0.58175594,0.43338865,0.28892577,0.14446288,0.0,0.19131571,0.38653582,0.57785153,0.76916724,0.96438736,1.33921,1.717937,2.096664,2.4714866,2.8502135,3.0024853,3.154757,3.3070288,3.4593005,3.611572,4.3338866,5.0522966,5.7707067,6.493021,7.211431,7.7307167,8.253906,8.773191,9.292478,9.811763,9.526741,9.237816,8.94889,8.663869,8.374943,9.331521,10.284196,11.240774,12.193448,13.150026,13.274967,13.399908,13.524849,13.64979,13.774731,13.2788725,12.786918,12.291059,11.795199,11.29934,10.573121,9.850807,9.124588,8.398369,7.676055,7.191909,6.703859,6.2197127,5.735567,5.251421,5.056201,4.8648853,4.6735697,4.478349,4.2870336,4.6384296,4.985922,5.337318,5.688714,6.036206,5.5989127,5.1616197,4.7243266,4.2870336,3.8497405,4.513489,5.181142,5.84489,6.5086384,7.1762915,6.6257706,6.0752497,5.5247293,4.9742084,4.423688,4.50568,4.591577,4.6735697,4.755562,4.8375545,5.02887,5.2162814,5.407597,5.5989127,5.786324,5.3177958,4.8492675,4.376835,3.9083066,3.435874,3.2445583,3.0532427,2.8619268,2.6667068,2.475391,2.377781,2.280171,2.182561,2.084951,1.9873407,2.3465457,2.7057507,3.06886,3.4280653,3.78727,3.4788225,3.174279,2.8658314,2.5573835,2.2489357,2.2684577,2.2840753,2.3035975,2.3192148,2.338737,2.1435168,1.9522011,1.7608855,1.5656652,1.3743496,1.397776,1.4212024,1.4407244,1.4641509,1.4875772,1.6867018,1.8858263,2.0888553,2.2879796,2.4871042,2.639376,2.7916477,2.9439192,3.096191,3.2484627,3.3265507,3.4007344,3.474918,3.5491016,3.6232853,4.0332475,4.4393053,4.8492675,5.2553253,5.661383,6.1455293,6.6257706,7.1099167,7.5940623,8.074304,7.57454,7.0747766,6.575013,6.0752497,5.575486,5.134289,4.689187,4.2479897,3.8067923,3.3616903,3.767748,4.173806,4.575959,4.9820175,5.388075,5.3724575,5.35684,5.3412223,5.3256044,5.3138914,5.12648,4.939069,4.7516575,4.564246,4.376835,5.520825,6.6648145,7.8088045,8.956698,10.100689,9.882042,9.663396,9.448653,9.230007,9.01136,13.243732,17.4722,21.704573,25.93304,30.161507,25.429373,20.697237,15.965101,11.232965,6.5008297,7.601871,8.706817,9.807858,10.9089,12.013845,14.848442,17.683039,20.517633,23.35223,26.186827,28.623173,31.063425,33.49977,35.93612,38.37637,35.15914,31.941916,28.720783,25.503555,22.286327,21.97788,21.669432,21.35708,21.048632,20.73628,24.578213,28.416239,32.25817,36.0962,39.93813,37.618916,35.303604,32.98439,30.669079,28.349865,27.479183,26.608501,25.741724,24.871042,24.00036,23.855898,23.711435,23.563068,23.418604,23.274141,22.7041,22.134056,21.564014,20.99397,20.423927,19.233086,18.038338,16.847496,15.656653,14.461906,12.771299,11.076789,9.386183,7.6916723,6.001066,4.911738,3.8185053,2.7291772,1.639849,0.5505207,0.98000497,1.4094892,1.8389735,2.2684577,2.7018464,3.1977055,3.6935644,4.193328,4.689187,5.1889505,6.473499,7.7619514,9.050405,10.338858,11.623405,12.291059,12.958711,13.626364,14.294017,14.96167,13.091461,11.217348,9.343235,7.473026,5.5989127,4.5017757,3.4007344,2.2996929,1.1986516,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14836729,0.30063897,0.44900626,0.60127795,0.74964523,0.7418364,0.7301232,0.71841,0.7106012,0.698888,0.74574083,0.78868926,0.8355421,0.8784905,0.92534333,1.1010414,1.2806439,1.456342,1.6359446,1.8116426,1.9092526,2.0029583,2.096664,2.194274,2.2879796,2.5964274,2.9087796,3.2172275,3.5256753,3.8380275,3.7091823,3.5842414,3.455396,3.3265507,3.2016098,3.1586614,3.1196175,3.0805733,3.0415294,2.998581,3.3929255,3.7833657,4.1777105,4.5681505,4.9624953,5.645766,6.3329406,7.016211,7.703386,8.386656,8.234385,8.078208,7.9220324,7.7658563,7.6135845,7.605776,7.601871,7.5979667,7.5940623,7.5862536,8.632633,9.679013,10.721489,11.767868,12.814248,12.845484,12.8767185,12.911859,12.943093,12.974329,15.168603,17.366781,19.561056,21.75533,23.949604,20.080341,16.214983,12.34572,8.480362,4.6110992,4.0605783,3.513962,2.9634414,2.4129205,1.8623998,2.1708477,2.4792955,2.7838387,3.0922866,3.4007344,3.9317331,4.4588275,4.989826,5.520825,6.0518236,6.7975645,7.5433054,8.292951,9.0386915,9.788337,10.510651,11.23687,11.963089,12.689307,13.411622,13.704452,13.993378,14.282304,14.571229,14.864059,18.264793,21.665527,25.070168,28.470901,31.87554,29.564135,27.256632,24.945227,22.63382,20.326319,19.795319,19.26432,18.733322,18.206228,17.675228,15.028045,12.384764,9.741484,7.094299,4.4510183,3.6349986,2.8189783,2.0068626,1.1908426,0.37482262,1.6867018,2.998581,4.3143644,5.6262436,6.9381227,6.356367,5.7707067,5.1889505,4.607195,4.025439,3.5100577,2.9946766,2.4792955,1.9639144,1.4485333,1.43682,1.4212024,1.4055848,1.3899672,1.3743496,1.2142692,1.0541886,0.8941081,0.7340276,0.57394713,0.5583295,0.5466163,0.5309987,0.5153811,0.4997635,0.45681506,0.41386664,0.3709182,0.3318742,0.28892577,0.47633708,0.6637484,0.8511597,1.038571,1.2259823,1.8584955,2.4910088,3.1235218,3.7560349,4.388548,5.087436,5.786324,6.4891167,7.1880045,7.8868923,7.137247,6.387602,5.6379566,4.8883114,4.138666,5.138193,6.141625,7.1450562,8.148487,9.151918,10.198298,11.2446785,12.291059,13.341343,14.387722,12.486279,10.58093,8.679486,6.7780423,4.8765984,4.318269,3.7599394,3.2016098,2.6432803,2.0888553,2.2879796,2.4871042,2.6862288,2.8892577,3.0883822,3.0337205,2.9829633,2.9283018,2.8775444,2.8267872,3.0532427,3.2836022,3.513962,3.7443218,3.9746814,4.263607,4.548629,4.8375545,5.12648,5.4115014,5.5442514,5.6730967,5.801942,5.930787,6.0635366,6.7663293,7.4691215,8.171914,8.870802,9.573594,10.81129,12.0489855,13.286681,14.524376,15.762072,14.254972,12.747873,11.240774,9.733675,8.226576,7.4964523,6.7663293,6.036206,5.3060827,4.575959,4.630621,4.6852827,4.7399445,4.794606,4.8492675,4.560342,4.271416,3.978586,3.68966,3.4007344,3.1157131,2.8345962,2.5534792,2.2684577,1.9873407,1.8819219,1.7725986,1.6632754,1.5578566,1.4485333,1.4680552,1.4914817,1.5110037,1.5305257,1.5500476,1.4133936,1.2767396,1.1361811,0.999527,0.8628729,2.2098918,3.5569105,4.903929,6.250948,7.601871,7.7619514,7.918128,8.078208,8.238289,8.398369,0.7262188,0.7106012,0.698888,0.6871748,0.6754616,0.6637484,0.6676528,0.6715572,0.679366,0.6832704,0.6871748,0.7066968,0.7223144,0.7418364,0.75745404,0.77307165,0.8160201,0.8550641,0.8941081,0.93315214,0.97610056,1.0307622,1.0893283,1.1478943,1.2064602,1.261122,1.4016805,1.5383345,1.6749885,1.8116426,1.9482968,2.4246337,2.900971,3.3734035,3.8497405,4.3260775,4.657952,4.989826,5.3217,5.6535745,5.989353,5.9737353,5.9620223,5.950309,5.938596,5.9268827,6.17286,6.4188375,6.6687193,6.914696,7.1606736,8.706817,10.249056,11.791295,13.333533,14.875772,14.418958,13.966047,13.509232,13.056321,12.599506,13.392099,14.184693,14.977287,15.76988,16.562475,13.575606,10.588739,7.5979667,4.6110992,1.6242313,1.3118792,0.9956226,0.679366,0.3631094,0.05075723,0.05466163,0.058566034,0.06637484,0.07027924,0.07418364,0.18741131,0.30063897,0.41386664,0.5231899,0.63641757,0.5114767,0.38263142,0.25378615,0.12884527,0.0,0.14836729,0.29673457,0.44119745,0.58956474,0.737932,1.0815194,1.4212024,1.7647898,2.1083772,2.4480603,2.893162,3.3343596,3.7794614,4.220659,4.661856,5.5169206,6.36808,7.2192397,8.074304,8.925464,9.515028,10.104593,10.694158,11.283723,11.873287,11.599979,11.326671,11.0494585,10.77615,10.498938,11.174399,11.845957,12.517513,13.189071,13.860628,13.848915,13.837202,13.825488,13.813775,13.798158,13.411622,13.021181,12.630741,12.240301,11.849861,11.475039,11.100216,10.725393,10.350571,9.975748,9.280765,8.58578,7.890797,7.195813,6.5008297,6.0908675,5.6809053,5.270943,4.860981,4.4510183,4.8883114,5.3256044,5.7628975,6.2001905,6.6374836,6.1611466,5.688714,5.212377,4.73604,4.263607,4.853172,5.446641,6.04011,6.6335793,7.223144,6.688241,6.1494336,5.610626,5.0757227,4.5369153,4.564246,4.591577,4.618908,4.646239,4.6735697,4.8805027,5.083532,5.290465,5.493494,5.700427,5.2592297,4.8219366,4.380739,3.9395418,3.4983444,3.338264,3.1781836,3.018103,2.8619268,2.7018464,2.631567,2.5612879,2.4910088,2.4207294,2.35045,2.7447948,3.1391394,3.533484,3.9317331,4.3260775,4.095718,3.8692627,3.6428072,3.416352,3.1859922,3.0102942,2.8306916,2.6549935,2.4792955,2.2996929,2.0654287,1.8311646,1.5969005,1.358732,1.1244678,1.1557031,1.1908426,1.2220778,1.2533131,1.2884527,1.4875772,1.6867018,1.8858263,2.0888553,2.2879796,2.416825,2.5456703,2.67842,2.8072653,2.9361105,3.0259118,3.1118085,3.2016098,3.2875066,3.3734035,3.8263142,4.279225,4.732136,5.185046,5.6379566,6.0518236,6.46569,6.883461,7.297328,7.7111945,7.113821,6.5125427,5.911265,5.3138914,4.7126136,4.3416953,3.9668727,3.5959544,3.2211318,2.8502135,3.2094188,3.5686235,3.9317331,4.290938,4.650143,4.7204223,4.7907014,4.860981,4.93126,5.001539,4.8375545,4.6735697,4.513489,4.349504,4.1894236,5.290465,6.3915067,7.4964523,8.597494,9.698535,9.452558,9.20658,8.956698,8.710721,8.460839,12.872814,17.280884,21.69286,26.10093,30.512903,25.772959,21.033014,16.29307,11.553126,6.813182,7.37932,7.9493628,8.515501,9.081639,9.651682,11.896713,14.141745,16.386776,18.631807,20.876839,23.223385,25.573835,27.924286,30.274734,32.625187,29.95067,27.280058,24.605543,21.934933,19.26432,18.9793,18.698183,18.41316,18.132044,17.850927,21.903696,25.960371,30.017044,34.069813,38.126488,36.127434,34.12838,32.133232,30.134176,28.139027,27.283962,26.432804,25.581644,24.72658,23.87542,23.922272,23.969126,24.015978,24.066736,24.113588,22.57135,21.033014,19.490776,17.952442,16.414106,15.328683,14.243259,13.157836,12.072412,10.986988,9.690726,8.3944645,7.094299,5.7980375,4.5017757,3.6818514,2.8658314,2.0459068,1.2298868,0.41386664,1.1361811,1.8584955,2.5808098,3.3031244,4.025439,4.193328,4.365122,4.5369153,4.704805,4.8765984,6.223617,7.57454,8.925464,10.276386,11.623405,12.24811,12.86891,13.493614,14.114414,14.739119,12.892336,11.0494585,9.202676,7.355894,5.5130157,4.423688,3.338264,2.2489357,1.1635119,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28892577,0.57394713,0.8628729,1.1517987,1.43682,1.3782539,1.3235924,1.2650263,1.2064602,1.1517987,1.2142692,1.2806439,1.3431144,1.4094892,1.475864,1.7921207,2.1083772,2.4285383,2.7447948,3.0610514,2.9907722,2.9165885,2.8463092,2.7721257,2.7018464,2.9087796,3.1157131,3.3226464,3.5295796,3.736513,3.7208953,3.7013733,3.6857557,3.6662338,3.6506162,3.7091823,3.7638438,3.8224099,3.8809757,3.9356375,4.447114,4.958591,5.466163,5.9776397,6.4891167,7.394938,8.300759,9.2104845,10.116306,11.0260315,10.729298,10.4286585,10.131924,9.835189,9.538455,9.24172,8.941081,8.644346,8.347612,8.050878,9.101162,10.155351,11.205634,12.259823,13.314012,13.528754,13.743496,13.958238,14.17298,14.387722,15.7035055,17.019289,18.33117,19.646952,20.962736,18.600573,16.242313,13.884054,11.521891,9.163632,7.6135845,6.0635366,4.513489,2.9634414,1.4133936,2.077142,2.7408905,3.408543,4.0722914,4.73604,5.1108627,5.481781,5.8566036,6.2275214,6.5984397,7.519879,8.441318,9.358852,10.280292,11.20173,12.08803,12.974329,13.860628,14.750832,15.637131,16.242313,16.847496,17.452679,18.057861,18.663042,21.868557,25.074072,28.27568,31.481195,34.68671,32.640804,30.5988,28.552895,26.506987,24.46108,22.31366,20.166237,18.018816,15.871395,13.723974,11.6468315,9.56969,7.492548,5.4154058,3.338264,2.8189783,2.3035975,1.7843118,1.2689307,0.74964523,2.7486992,4.7516575,6.7507114,8.749765,10.748819,9.511124,8.269524,7.0318284,5.7902284,4.548629,3.8575494,3.1664703,2.4714866,1.7804074,1.0893283,1.4212024,1.7530766,2.084951,2.416825,2.7486992,2.4285383,2.1083772,1.7882162,1.4680552,1.1517987,1.0932326,1.038571,0.98390937,0.92924774,0.8745861,0.75354964,0.62860876,0.5075723,0.38653582,0.26159495,0.46071947,0.6637484,0.8628729,1.0619974,1.261122,1.7765031,2.2918842,2.8072653,3.3226464,3.8380275,4.4002614,4.9624953,5.5247293,6.086963,6.649197,6.2001905,5.7511845,5.298274,4.8492675,4.4002614,5.368553,6.336845,7.3012323,8.269524,9.237816,10.670732,12.103647,13.536563,14.965574,16.398489,14.594656,12.790822,10.983084,9.17925,7.375416,6.66091,5.9464045,5.2318993,4.513489,3.7989833,3.78727,3.775557,3.7638438,3.7482262,3.736513,3.506153,3.2757936,3.049338,2.8189783,2.5886188,2.7330816,2.8814487,3.0298162,3.1781836,3.3265507,3.5491016,3.775557,3.998108,4.224563,4.4510183,4.548629,4.646239,4.743849,4.841459,4.939069,5.716045,6.4969254,7.277806,8.058686,8.835662,10.276386,11.713207,13.150026,14.586847,16.023666,14.422862,12.818152,11.217348,9.616543,8.011833,7.266093,6.5164475,5.7707067,5.0210614,4.2753205,4.2362766,4.193328,4.154284,4.11524,4.0761957,3.9083066,3.7404175,3.5725281,3.4046388,3.2367494,3.084478,2.9322062,2.7799344,2.6276627,2.475391,2.3231194,2.1708477,2.018576,1.8663043,1.7140326,1.678893,1.6437533,1.6086137,1.5734742,1.5383345,1.3860629,1.2376955,1.0893283,0.93705654,0.78868926,2.494913,4.2011366,5.911265,7.617489,9.323712,9.108971,8.890324,8.671678,8.456935,8.238289,0.7106012,0.698888,0.6871748,0.6754616,0.6637484,0.6481308,0.6559396,0.6637484,0.6715572,0.679366,0.6871748,0.7066968,0.7262188,0.74574083,0.76916724,0.78868926,0.8238289,0.8589685,0.8941081,0.92924774,0.96438736,1.0190489,1.0737107,1.1283722,1.183034,1.2376955,1.4133936,1.5890918,1.7608855,1.9365835,2.1122816,2.6862288,3.2640803,3.8380275,4.4119744,4.985922,5.142098,5.298274,5.45445,5.606722,5.7628975,5.8487945,5.938596,6.0244927,6.114294,6.2001905,6.4383593,6.6804323,6.918601,7.1606736,7.3988423,9.019169,10.639496,12.259823,13.88015,15.500477,14.942147,14.383818,13.829392,13.271063,12.712734,13.821584,14.92653,16.03538,17.14423,18.249176,14.899199,11.549222,8.1992445,4.8492675,1.4992905,1.2142692,0.92924774,0.6442264,0.359205,0.07418364,0.07027924,0.06637484,0.058566034,0.05466163,0.05075723,0.14836729,0.24988174,0.3513962,0.44900626,0.5505207,0.44119745,0.3318742,0.21864653,0.10932326,0.0,0.10151446,0.20693332,0.30844778,0.40996224,0.5114767,0.8199245,1.1283722,1.43682,1.7413634,2.0498111,2.7838387,3.513962,4.2479897,4.9781127,5.7121406,6.6960497,7.6838636,8.667773,9.651682,10.6355915,11.29934,11.959184,12.619028,13.2788725,13.938716,13.673217,13.411622,13.150026,12.888432,12.626837,13.013372,13.403813,13.794253,14.184693,14.575133,14.426766,14.274494,14.126127,13.973856,13.825488,13.540467,13.2554455,12.970425,12.685403,12.400381,12.373051,12.349625,12.326198,12.298867,12.27544,11.369619,10.4637985,9.561881,8.65606,7.7502384,7.1216297,6.4969254,5.8683167,5.239708,4.6110992,5.138193,5.661383,6.1884775,6.7116675,7.238762,6.7233806,6.211904,5.700427,5.1889505,4.6735697,5.196759,5.716045,6.2353306,6.754616,7.2739015,6.7507114,6.223617,5.700427,5.173333,4.650143,4.6228123,4.5954814,4.5681505,4.5408196,4.513489,4.732136,4.950782,5.173333,5.3919797,5.610626,5.2006636,4.7907014,4.380739,3.970777,3.5608149,3.435874,3.3070288,3.1781836,3.0532427,2.9243972,2.8814487,2.8385005,2.795552,2.7565079,2.7135596,3.1430438,3.5725281,4.0020123,4.4314966,4.860981,4.716518,4.5681505,4.4197836,4.271416,4.123049,3.7521305,3.3812122,3.0063896,2.6354716,2.260649,1.9834363,1.7062237,1.4290112,1.1517987,0.8745861,0.91753453,0.96048295,1.0034313,1.0463798,1.0893283,1.2884527,1.4875772,1.6867018,1.8858263,2.0888553,2.194274,2.3035975,2.4090161,2.5183394,2.6237583,2.7252727,2.8267872,2.9243972,3.0259118,3.1235218,3.6232853,4.1191444,4.618908,5.114767,5.610626,5.958118,6.3056097,6.6531014,7.000593,7.348085,6.649197,5.950309,5.251421,4.548629,3.8497405,3.5491016,3.2445583,2.9439192,2.639376,2.338737,2.6510892,2.9673457,3.2836022,3.5959544,3.912211,4.068387,4.220659,4.376835,4.533011,4.689187,4.548629,4.4119744,4.2753205,4.138666,3.998108,5.0601053,6.1181984,7.180196,8.238289,9.300286,9.023073,8.745861,8.468649,8.191436,7.914223,12.501896,17.093473,21.681147,26.272722,30.8643,26.116547,21.368793,16.62104,11.873287,7.125534,7.1567693,7.191909,7.223144,7.2543793,7.2856145,8.941081,10.596548,12.252014,13.907481,15.562947,17.823597,20.08815,22.348799,24.613352,26.874,24.746101,22.618202,20.494207,18.366308,16.238409,15.980719,15.726933,15.473146,15.21936,14.96167,19.233086,23.500597,27.772013,32.04343,36.31094,34.635952,32.957058,31.278166,29.603178,27.924286,27.088743,26.2532,25.421562,24.586021,23.750479,23.988647,24.23072,24.46889,24.710962,24.949131,22.4386,19.931974,17.421442,14.9109125,12.400381,11.424281,10.444276,9.468176,8.488171,7.5120697,6.610153,5.708236,4.806319,3.9044023,2.998581,2.455869,1.9092526,1.3665408,0.8199245,0.27330816,1.2884527,2.3035975,3.3187418,4.3338866,5.349031,5.192855,5.036679,4.8765984,4.7204223,4.564246,5.9737353,7.387129,8.800523,10.213917,11.623405,12.201257,12.779109,13.35696,13.934812,14.512663,12.693212,10.877665,9.058213,7.2426662,5.423215,4.349504,3.2757936,2.1981785,1.1244678,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.42557985,0.8511597,1.2767396,1.698415,2.1239948,2.018576,1.9131571,1.8116426,1.7062237,1.6008049,1.6867018,1.7686942,1.8545911,1.9404879,2.0263848,2.4831998,2.9400148,3.39683,3.853645,4.3143644,4.0722914,3.8341231,3.59205,3.3538816,3.1118085,3.2172275,3.3226464,3.4280653,3.533484,3.638903,3.7287042,3.8224099,3.9161155,4.0059166,4.0996222,4.2557983,4.40807,4.564246,4.7204223,4.8765984,5.5013027,6.1299114,6.75852,7.3832245,8.011833,9.14411,10.272482,11.400854,12.533132,13.661504,13.224211,12.783013,12.341816,11.900618,11.4633255,10.87376,10.284196,9.690726,9.101162,8.511597,9.573594,10.631687,11.693685,12.751778,13.813775,14.208119,14.606369,15.004618,15.402867,15.801116,16.234505,16.671797,17.105186,17.538574,17.975868,17.120804,16.269644,15.418485,14.56342,13.712261,11.162686,8.6131115,6.0635366,3.513962,0.96438736,1.9834363,3.0063896,4.029343,5.0522966,6.0752497,6.289992,6.504734,6.719476,6.9342184,7.1489606,8.242193,9.335425,10.4286585,11.521891,12.611219,13.661504,14.711788,15.762072,16.812357,17.86264,18.784079,19.701614,20.623053,21.540586,22.462027,25.468416,28.47871,31.4851,34.49149,37.501785,35.721375,33.940968,32.16056,30.380154,28.599747,24.835903,21.07206,17.30431,13.540467,9.776623,8.265619,6.754616,5.2436123,3.736513,2.2255092,2.0068626,1.7843118,1.5656652,1.3431144,1.1244678,3.814601,6.5008297,9.187058,11.873287,14.56342,12.665881,10.768341,8.870802,6.9732623,5.0757227,4.2050414,3.3343596,2.463678,1.5969005,0.7262188,1.4055848,2.084951,2.7643168,3.4436827,4.123049,3.6467118,3.1664703,2.6862288,2.2059872,1.7257458,1.6281357,1.53443,1.4407244,1.3431144,1.2494087,1.0463798,0.8433509,0.6442264,0.44119745,0.23816854,0.44900626,0.6637484,0.8745861,1.0893283,1.3001659,1.698415,2.096664,2.4910088,2.8892577,3.2875066,3.7130866,4.138666,4.564246,4.985922,5.4115014,5.263134,5.1108627,4.9624953,4.814128,4.661856,5.5950084,6.5281606,7.461313,8.39056,9.323712,11.143164,12.958711,14.778163,16.59371,18.41316,16.703033,14.996809,13.2905855,11.584361,9.874233,9.0035515,8.128965,7.2582836,6.3836975,5.5130157,5.2865605,5.0640097,4.8375545,4.6110992,4.388548,3.978586,3.5725281,3.1664703,2.7565079,2.35045,2.416825,2.4792955,2.5456703,2.6081407,2.6745155,2.8385005,2.998581,3.1625657,3.3265507,3.4866312,3.5530062,3.619381,3.6818514,3.7482262,3.8106966,4.6696653,5.5286336,6.3836975,7.2426662,8.101635,9.737579,11.373524,13.013372,14.649317,16.289165,14.590752,12.892336,11.193921,9.499411,7.800996,7.0357327,6.27047,5.505207,4.7399445,3.9746814,3.8419318,3.7052777,3.5686235,3.435874,3.2992198,3.2562714,3.2094188,3.1664703,3.1196175,3.076669,3.0532427,3.0298162,3.0063896,2.9868677,2.9634414,2.7643168,2.5690966,2.3699722,2.1708477,1.9756275,1.8858263,1.796025,1.7062237,1.6164225,1.5266213,1.3626363,1.1986516,1.038571,0.8745861,0.7106012,2.7799344,4.8492675,6.914696,8.98403,11.0494585,10.455989,9.858616,9.265146,8.671678,8.074304,0.698888,0.6871748,0.6754616,0.6637484,0.6481308,0.63641757,0.6481308,0.6559396,0.6676528,0.679366,0.6871748,0.7106012,0.7340276,0.75354964,0.77697605,0.80040246,0.8316377,0.8589685,0.8902037,0.92143893,0.94876975,1.0034313,1.0541886,1.1088502,1.1596074,1.2142692,1.4251068,1.6359446,1.8506867,2.0615244,2.2762666,2.951728,3.6232853,4.298747,4.9742084,5.64967,5.6262436,5.606722,5.5832953,5.559869,5.5364423,5.7238536,5.911265,6.098676,6.2860875,6.473499,6.707763,6.9381227,7.172387,7.406651,7.6370106,9.335425,11.033841,12.728352,14.426766,16.125181,15.465338,14.805493,14.145649,13.4858055,12.825961,14.247164,15.668366,17.093473,18.514675,19.935879,16.226696,12.513609,8.800523,5.087436,1.3743496,1.1205635,0.8667773,0.60908675,0.3553006,0.10151446,0.08589685,0.07027924,0.05466163,0.039044023,0.023426414,0.113227665,0.19912452,0.28892577,0.37482262,0.46071947,0.3709182,0.27721256,0.1835069,0.093705654,0.0,0.058566034,0.113227665,0.1717937,0.23035973,0.28892577,0.5583295,0.8316377,1.1049459,1.3782539,1.6515622,2.6706111,3.6935644,4.716518,5.7394714,6.7624245,7.8790836,8.995743,10.116306,11.232965,12.349625,13.079747,13.809871,14.539994,15.270117,16.00024,15.750359,15.500477,15.250595,15.000713,14.750832,14.856251,14.965574,15.070992,15.180316,15.285735,15.000713,14.711788,14.426766,14.13784,13.848915,13.6693125,13.48971,13.310107,13.130505,12.950902,13.274967,13.599033,13.923099,14.251068,14.575133,13.458474,12.34572,11.229061,10.116306,8.999647,8.156297,7.309041,6.46569,5.618435,4.775084,5.388075,6.001066,6.6140575,7.223144,7.8361354,7.2856145,6.7389984,6.1884775,5.6379566,5.087436,5.5364423,5.9815445,6.4305506,6.8756523,7.3246584,6.813182,6.3017054,5.786324,5.2748475,4.7633705,4.6813784,4.5993857,4.513489,4.4314966,4.349504,4.5837684,4.8219366,5.056201,5.290465,5.5247293,5.1460023,4.7633705,4.3846436,4.0059166,3.6232853,3.5295796,3.435874,3.338264,3.2445583,3.1508527,3.135235,3.1196175,3.1039999,3.0883822,3.076669,3.541293,4.0059166,4.4705405,4.9351645,5.3997884,5.3334136,5.263134,5.196759,5.1303844,5.0640097,4.493967,3.9278288,3.3616903,2.7916477,2.2255092,1.9053483,1.5851873,1.2650263,0.94486535,0.62470436,0.679366,0.7301232,0.78088045,0.8355421,0.8862993,1.0893283,1.2884527,1.4875772,1.6867018,1.8858263,1.9717231,2.05762,2.1435168,2.2294137,2.3114061,2.4246337,2.5378613,2.6510892,2.7643168,2.87364,3.416352,3.959064,4.5017757,5.044488,5.5871997,5.8683167,6.1494336,6.426646,6.707763,6.98888,6.1884775,5.388075,4.5876727,3.78727,2.9868677,2.7565079,2.522244,2.2918842,2.05762,1.8233559,2.096664,2.366068,2.6354716,2.9048753,3.174279,3.416352,3.6545205,3.8965936,4.134762,4.376835,4.263607,4.1503797,4.037152,3.9239242,3.8106966,4.829746,5.8487945,6.8639393,7.882988,8.898132,8.59359,8.285142,7.9766936,7.6682463,7.363703,12.130978,16.902157,21.673336,26.444517,31.211792,26.45623,21.704573,16.94901,12.193448,7.437886,6.9342184,6.434455,5.930787,5.4271193,4.9234514,5.989353,7.055255,8.121157,9.183154,10.249056,12.423808,14.59856,16.773312,18.948065,21.12672,19.541533,17.96025,16.378967,14.79378,13.212498,12.986042,12.755682,12.529227,12.302772,12.076316,16.55857,21.044727,25.530886,30.01314,34.4993,33.140568,31.785738,30.427008,29.068275,27.713448,26.893522,26.077503,25.261482,24.441559,23.625538,24.058928,24.48841,24.921799,25.355188,25.788576,22.305851,18.827028,15.348206,11.8654785,8.386656,7.5159745,6.649197,5.7785153,4.9078336,4.037152,3.5295796,3.0220075,2.514435,2.0068626,1.4992905,1.2259823,0.95657855,0.6832704,0.40996224,0.13665408,1.4446288,2.7526035,4.0605783,5.368553,6.676528,6.1884775,5.704332,5.2201858,4.73604,4.251894,5.7238536,7.1997175,8.675582,10.151445,11.623405,12.158309,12.689307,13.224211,13.755209,14.286208,12.497992,10.705871,8.917655,7.125534,5.337318,4.2753205,3.213323,2.1513257,1.0893283,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5622339,1.1244678,1.6867018,2.2489357,2.8111696,2.6588979,2.5066261,2.3543546,2.2020829,2.0498111,2.15523,2.260649,2.366068,2.4714866,2.5769055,3.174279,3.7716527,4.369026,4.9663997,5.563773,5.153811,4.747753,4.3416953,3.9317331,3.5256753,3.5256753,3.5295796,3.533484,3.533484,3.5373883,3.7404175,3.9434462,4.1464753,4.3455997,4.548629,4.802415,5.056201,5.3060827,5.559869,5.813655,6.559396,7.3012323,8.046973,8.792714,9.538455,10.889378,12.244205,13.595129,14.946052,16.300879,15.719124,15.133463,14.551707,13.969952,13.388195,12.5058,11.623405,10.741011,9.858616,8.976221,10.042123,11.108025,12.177831,13.243732,14.313539,14.89139,15.473146,16.050997,16.632753,17.210606,16.769407,16.324306,15.879204,15.434102,14.989,15.641035,16.296974,16.952915,17.608854,18.26089,14.711788,11.162686,7.6135845,4.0605783,0.5114767,1.893635,3.2718892,4.6540475,6.0323014,7.4144597,7.4691215,7.5276875,7.5862536,7.6409154,7.699481,8.964508,10.229534,11.49456,12.759586,14.024612,15.238882,16.449247,17.663515,18.87388,20.08815,21.321941,22.555733,23.793427,25.027218,26.26101,29.07218,31.883348,34.69452,37.501785,40.312954,38.798046,37.28314,35.76823,34.253323,32.738415,27.354242,21.973976,16.589806,11.205634,5.825368,4.8805027,3.9395418,2.998581,2.0537157,1.1127546,1.1908426,1.2689307,1.3431144,1.4212024,1.4992905,4.8765984,8.250002,11.623405,15.000713,18.374117,15.820638,13.263254,10.709775,8.156297,5.5989127,4.552533,3.506153,2.455869,1.4094892,0.3631094,1.3899672,2.416825,3.4436827,4.474445,5.5013027,4.860981,4.220659,3.5803368,2.9400148,2.2996929,2.1669433,2.0302892,1.893635,1.7608855,1.6242313,1.3431144,1.0580931,0.77697605,0.4958591,0.21083772,0.43729305,0.6637484,0.8862993,1.1127546,1.33921,1.6164225,1.8975395,2.1786566,2.455869,2.736986,3.0259118,3.310933,3.5998588,3.8887846,4.173806,4.3260775,4.474445,4.6267166,4.775084,4.9234514,5.8214636,6.719476,7.617489,8.515501,9.413514,11.615597,13.817679,16.019762,18.221846,20.423927,18.815315,17.206701,15.594183,13.985569,12.376955,11.346193,10.315431,9.284669,8.253906,7.223144,6.785851,6.348558,5.911265,5.473972,5.036679,4.4510183,3.8692627,3.2836022,2.697942,2.1122816,2.096664,2.077142,2.0615244,2.0420024,2.0263848,2.1239948,2.2255092,2.3231194,2.4246337,2.5261483,2.5573835,2.5886188,2.6237583,2.6549935,2.6862288,3.6232853,4.5564375,5.493494,6.426646,7.363703,9.198771,11.037745,12.8767185,14.711788,16.55076,14.75864,12.96652,11.170495,9.378374,7.5862536,6.805373,6.0205884,5.239708,4.4588275,3.6740425,3.4436827,3.213323,2.9868677,2.7565079,2.5261483,2.6042364,2.67842,2.7565079,2.8345962,2.912684,3.018103,3.1274261,3.2367494,3.3421683,3.4514916,3.2094188,2.9634414,2.7213683,2.4792955,2.2372224,2.0927596,1.9482968,1.8038338,1.6593709,1.5110037,1.33921,1.1635119,0.9878138,0.81211567,0.63641757,3.0649557,5.493494,7.9220324,10.346666,12.775204,11.803008,10.8308115,9.858616,8.886419,7.914223,0.6871748,0.6754616,0.6637484,0.6481308,0.63641757,0.62470436,0.63641757,0.6481308,0.6637484,0.6754616,0.6871748,0.7106012,0.737932,0.76135844,0.78868926,0.81211567,0.8394465,0.8628729,0.8862993,0.9136301,0.93705654,0.9878138,1.038571,1.0893283,1.1361811,1.1869383,1.43682,1.6867018,1.9365835,2.1864653,2.436347,3.213323,3.9863946,4.7633705,5.5364423,6.3134184,6.114294,5.911265,5.7121406,5.5130157,5.3138914,5.5989127,5.8878384,6.1767645,6.461786,6.7507114,6.9732623,7.1997175,7.426173,7.648724,7.8751793,9.651682,11.424281,13.200784,14.973383,16.749886,15.988527,15.223265,14.461906,13.700547,12.939189,14.676648,16.414106,18.151566,19.889025,21.626484,17.550287,13.4740925,9.4018,5.3256044,1.2494087,1.0268579,0.80040246,0.57394713,0.3513962,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.30063897,0.5388075,0.77307165,1.0112402,1.2494087,2.5612879,3.873167,5.1889505,6.5008297,7.812709,9.062118,10.311526,11.560935,12.814248,14.063657,14.864059,15.660558,16.46096,17.261362,18.061766,17.823597,17.589333,17.351164,17.112995,16.874826,16.69913,16.52343,16.351637,16.175938,16.00024,15.57466,15.14908,14.723501,14.301826,13.8762455,13.798158,13.723974,13.64979,13.575606,13.501423,14.176885,14.848442,15.523903,16.199366,16.874826,15.551234,14.223738,12.900145,11.576552,10.249056,9.187058,8.125061,7.0630636,6.001066,4.939069,5.6379566,6.336845,7.0357327,7.7385254,8.437413,7.8517528,7.262188,6.676528,6.086963,5.5013027,5.8761253,6.250948,6.6257706,7.000593,7.375416,6.8756523,6.375889,5.8761253,5.376362,4.8765984,4.73604,4.5993857,4.462732,4.3260775,4.1894236,4.4393053,4.689187,4.939069,5.1889505,5.4388323,5.087436,4.73604,4.388548,4.037152,3.6857557,3.6232853,3.5608149,3.4983444,3.435874,3.3734035,3.3890212,3.4007344,3.4124475,3.4241607,3.435874,3.9356375,4.4393053,4.939069,5.4388323,5.938596,5.950309,5.9620223,5.9737353,5.989353,6.001066,5.2358036,4.474445,3.7130866,2.951728,2.1864653,1.8233559,1.4641509,1.1010414,0.737932,0.37482262,0.43729305,0.4997635,0.5622339,0.62470436,0.6871748,0.8862993,1.0893283,1.2884527,1.4875772,1.6867018,1.7491722,1.8116426,1.8741131,1.9365835,1.999054,2.1239948,2.2489357,2.3738766,2.4988174,2.6237583,3.213323,3.7989833,4.388548,4.9742084,5.563773,5.774611,5.989353,6.2001905,6.4110284,6.6257706,5.7238536,4.825841,3.9239242,3.0259118,2.1239948,1.9639144,1.7999294,1.6359446,1.475864,1.3118792,1.5383345,1.7608855,1.9873407,2.2137961,2.436347,2.7643168,3.0883822,3.4124475,3.736513,4.0605783,3.9746814,3.8887846,3.7989833,3.7130866,3.6232853,4.5993857,5.575486,6.551587,7.523783,8.499884,8.164105,7.824422,7.4886436,7.1489606,6.813182,11.763964,16.710842,21.661623,26.612406,31.563189,26.799816,22.036446,17.273075,12.513609,7.7502384,6.7116675,5.6730967,4.6384296,3.5998588,2.5612879,3.0376248,3.513962,3.9863946,4.462732,4.939069,7.0240197,9.112875,11.20173,13.286681,15.375536,14.336966,13.298394,12.263727,11.225157,10.186585,9.987461,9.788337,9.589212,9.386183,9.187058,13.887959,18.58886,23.285854,27.986755,32.687656,31.649084,30.614418,29.575848,28.537275,27.498705,26.698303,25.901804,25.101402,24.300999,23.500597,24.125301,24.750006,25.37471,25.999414,26.624119,22.1731,17.725986,13.274967,8.823949,4.376835,3.611572,2.8502135,2.0888553,1.3235924,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.0,0.0,0.0,0.0,0.0,1.6008049,3.2016098,4.7985106,6.3993154,8.00012,7.1880045,6.375889,5.563773,4.7516575,3.9356375,5.473972,7.012306,8.550641,10.088976,11.623405,12.111456,12.599506,13.087557,13.575606,14.063657,12.298867,10.537982,8.773191,7.012306,5.251421,4.2011366,3.1508527,2.1005683,1.0502841,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.698888,1.4016805,2.1005683,2.7994564,3.4983444,3.2992198,3.1000953,2.900971,2.7018464,2.4988174,2.6237583,2.7486992,2.87364,2.998581,3.1235218,3.8614538,4.5993857,5.337318,6.0752497,6.813182,6.239235,5.661383,5.087436,4.513489,3.9356375,3.8380275,3.736513,3.638903,3.5373883,3.435874,3.7482262,4.0605783,4.376835,4.689187,5.001539,5.349031,5.700427,6.0518236,6.3993154,6.7507114,7.6135845,8.476458,9.339331,10.198298,11.061172,12.63855,14.212025,15.789403,17.362877,18.936352,18.214037,17.487818,16.761599,16.039284,15.313066,14.13784,12.962616,11.787391,10.612165,9.43694,10.510651,11.588266,12.661977,13.735687,14.813302,15.57466,16.33602,17.101282,17.86264,18.623999,17.300406,15.976814,14.649317,13.325725,11.998228,14.161267,16.324306,18.487345,20.650383,22.813423,18.26089,13.712261,9.163632,4.6110992,0.062470436,1.7999294,3.5373883,5.2748475,7.012306,8.749765,8.648251,8.550641,8.449126,8.351517,8.250002,9.686822,11.123642,12.564366,14.001186,15.438006,16.812357,18.186707,19.561056,20.93931,22.31366,23.863707,25.413754,26.963802,28.51385,30.063898,32.67594,35.287987,37.900032,40.512077,43.124123,41.874714,40.625305,39.375896,38.126488,36.873177,29.876486,22.875893,15.875299,8.874706,1.8741131,1.4992905,1.1244678,0.74964523,0.37482262,0.0,0.37482262,0.74964523,1.1244678,1.4992905,1.8741131,5.938596,9.999174,14.063657,18.124235,22.188719,18.975395,15.762072,12.548749,9.339331,6.126007,4.900025,3.6740425,2.4480603,1.2259823,0.0,1.3743496,2.7486992,4.126953,5.5013027,6.8756523,6.0752497,5.2748475,4.474445,3.6740425,2.87364,2.7018464,2.5261483,2.35045,2.174752,1.999054,1.6359446,1.2767396,0.9136301,0.5505207,0.18741131,0.42557985,0.6637484,0.9019169,1.1361811,1.3743496,1.5383345,1.698415,1.8623998,2.0263848,2.1864653,2.338737,2.4871042,2.639376,2.787743,2.9361105,3.3890212,3.8380275,4.2870336,4.73604,5.1889505,6.0518236,6.910792,7.773665,8.636538,9.499411,12.08803,14.676648,17.261362,19.849981,22.4386,20.92369,19.412687,17.901684,16.386776,14.875772,13.688834,12.501896,11.311053,10.124115,8.937177,8.289046,7.6370106,6.98888,6.336845,5.688714,4.9234514,4.1620927,3.4007344,2.639376,1.8741131,1.7765031,1.6749885,1.5734742,1.475864,1.3743496,1.4133936,1.4485333,1.4875772,1.5266213,1.5617609,1.5617609,1.5617609,1.5617609,1.5617609,1.5617609,2.5769055,3.5881457,4.5993857,5.610626,6.6257706,8.663869,10.701966,12.73616,14.774258,16.812357,14.92653,13.036799,11.150972,9.261242,7.375416,6.575013,5.774611,4.9742084,4.173806,3.3734035,3.049338,2.7252727,2.4012074,2.0732377,1.7491722,1.9482968,2.1513257,2.35045,2.5495746,2.7486992,2.9868677,3.2250361,3.4632049,3.7013733,3.9356375,3.6506162,3.3616903,3.076669,2.787743,2.4988174,2.2996929,2.1005683,1.901444,1.698415,1.4992905,1.3118792,1.1244678,0.93705654,0.74964523,0.5622339,3.349977,6.13772,8.925464,11.713207,14.50095,13.150026,11.799104,10.44818,9.101162,7.7502384,0.6754616,0.6676528,0.659844,0.6520352,0.6442264,0.63641757,0.6559396,0.6715572,0.6910792,0.7066968,0.7262188,0.74574083,0.76916724,0.79259366,0.8160201,0.8394465,0.8511597,0.8628729,0.8745861,0.8862993,0.9019169,0.96438736,1.0268579,1.0893283,1.1517987,1.2142692,1.4641509,1.7140326,1.9639144,2.2137961,2.463678,3.0727646,3.6818514,4.290938,4.903929,5.5130157,5.376362,5.2358036,5.099149,4.9624953,4.825841,5.388075,5.9542136,6.520352,7.08649,7.648724,7.9376497,8.226576,8.511597,8.800523,9.089449,10.612165,12.138786,13.661504,15.188125,16.710842,16.136894,15.562947,14.989,14.411149,13.837202,14.582942,15.328683,16.074425,16.816261,17.562002,14.251068,10.936231,7.6252975,4.3143644,0.999527,0.9136301,0.8238289,0.737932,0.6481308,0.5622339,0.698888,0.8394465,0.97610056,1.1127546,1.2494087,1.2650263,1.2806439,1.2962615,1.3118792,1.3235924,1.3157835,1.3040704,1.2962615,1.2845483,1.2767396,1.1439898,1.0151446,0.8862993,0.75354964,0.62470436,0.7301232,0.8355421,0.94096094,1.0463798,1.1517987,2.787743,4.423688,6.0635366,7.699481,9.339331,11.268105,13.200784,15.133463,17.066143,18.998821,19.080814,19.16671,19.248703,19.330696,19.412687,18.787983,18.163279,17.538574,16.91387,16.289165,16.066616,15.844065,15.621513,15.398962,15.176412,14.883581,14.590752,14.297921,14.005091,13.712261,13.6693125,13.622459,13.575606,13.532659,13.4858055,13.911386,14.336966,14.762545,15.188125,15.613705,14.454097,13.2905855,12.130978,10.971371,9.811763,8.94889,8.086017,7.223144,6.364176,5.5013027,6.016684,6.5281606,7.043542,7.558923,8.074304,7.648724,7.223144,6.801469,6.375889,5.950309,6.2860875,6.6257706,6.9615493,7.3012323,7.6370106,7.1606736,6.688241,6.211904,5.735567,5.263134,5.044488,4.825841,4.6110992,4.3924527,4.173806,4.4314966,4.689187,4.9468775,5.2045684,5.462259,5.3021784,5.142098,4.9820175,4.8219366,4.661856,4.5252023,4.388548,4.251894,4.1113358,3.9746814,3.8965936,3.8185053,3.7443218,3.6662338,3.5881457,3.970777,4.357313,4.743849,5.12648,5.5130157,5.5169206,5.520825,5.5286336,5.532538,5.5364423,4.83365,4.1308575,3.4280653,2.7291772,2.0263848,1.7921207,1.5617609,1.3274968,1.0932326,0.8628729,0.98390937,1.1088502,1.2298868,1.3509232,1.475864,1.5149081,1.5539521,1.5969005,1.6359446,1.6749885,1.7647898,1.8545911,1.9443923,2.0341935,2.1239948,2.2567444,2.3855898,2.514435,2.6432803,2.77603,3.416352,4.0605783,4.7009,5.3451266,5.989353,6.1884775,6.3915067,6.5945354,6.7975645,7.000593,6.13772,5.2748475,4.4119744,3.5491016,2.6862288,2.4910088,2.2918842,2.096664,1.8975395,1.698415,1.9443923,2.1903696,2.436347,2.67842,2.9243972,3.1391394,3.3538816,3.5686235,3.7833657,3.998108,3.9044023,3.8067923,3.7091823,3.611572,3.513962,4.3729305,5.2318993,6.0908675,6.9537406,7.812709,7.5159745,7.2192397,6.918601,6.621866,6.3251314,11.053363,15.781594,20.50592,25.234152,29.962383,25.589453,21.212618,16.835783,12.4628525,8.086017,6.98888,5.891743,4.794606,3.697469,2.6003318,2.8814487,3.1586614,3.4397783,3.7208953,3.998108,5.7824197,7.5667315,9.347139,11.131451,12.911859,12.216875,11.521891,10.826907,10.131924,9.43694,9.304191,9.167537,9.030883,8.898132,8.761478,13.013372,17.26917,21.521065,25.772959,30.024853,29.681267,29.333775,28.990187,28.646599,28.299107,27.764204,27.225397,26.68659,26.151686,25.612879,26.706112,27.80325,28.89648,29.993618,31.086851,25.905708,20.728472,15.54733,10.366188,5.1889505,4.376835,3.5686235,2.7565079,1.9482968,1.1361811,1.3782539,1.6164225,1.8584955,2.096664,2.338737,2.3933985,2.4519646,2.5105307,2.5690966,2.6237583,4.134762,5.645766,7.1567693,8.663869,10.174872,9.675109,9.175345,8.675582,8.175818,7.676055,8.636538,9.593117,10.553599,11.514082,12.4745655,12.47847,12.486279,12.490183,12.494087,12.501896,10.838621,9.17925,7.519879,5.860508,4.2011366,3.3616903,2.5183394,1.678893,0.8394465,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.3240654,0.44510186,0.5661383,0.6910792,0.81211567,1.2650263,1.717937,2.1708477,2.6237583,3.076669,2.9165885,2.7565079,2.5964274,2.436347,2.2762666,2.330928,2.3855898,2.4402514,2.494913,2.5495746,3.2211318,3.8965936,4.5681505,5.239708,5.911265,5.4271193,4.942973,4.4588275,3.970777,3.4866312,3.4202564,3.3538816,3.2836022,3.2172275,3.1508527,3.6349986,4.1191444,4.60329,5.0913405,5.575486,5.903456,6.2353306,6.5633,6.8951745,7.223144,8.191436,9.155824,10.120211,11.084598,12.0489855,13.009468,13.966047,14.922626,15.879204,16.835783,16.156416,15.473146,14.789876,14.106606,13.423335,12.544845,11.666354,10.783959,9.905469,9.023073,9.850807,10.67854,11.506273,12.334006,13.16174,13.907481,14.653222,15.398962,16.140799,16.88654,15.926057,14.96167,14.001186,13.036799,12.076316,14.145649,16.214983,18.284315,20.35365,22.426888,19.010534,15.601992,12.185639,8.773191,5.3607445,5.7980375,6.2314262,6.6687193,7.1021075,7.5394006,8.382751,9.226103,10.073358,10.916709,11.763964,12.548749,13.337439,14.126127,14.9109125,15.699601,16.624945,17.550287,18.475632,19.400974,20.326319,23.22729,26.12826,29.033134,31.934107,34.83898,34.819458,34.796032,34.776512,34.75699,34.73747,33.691086,32.648613,31.602232,30.555853,29.513376,23.953508,18.393639,12.83377,7.2739015,1.7140326,1.3704453,1.0268579,0.6832704,0.3435874,0.0,1.0659018,2.135708,3.2016098,4.271416,5.337318,7.968885,10.596548,13.228115,15.855778,18.487345,15.76988,13.052417,10.334952,7.617489,4.900025,4.029343,3.154757,2.2840753,1.4094892,0.5388075,2.069333,3.6037633,5.134289,6.6687193,8.1992445,7.9064145,7.60968,7.3168497,7.0201154,6.7233806,6.0713453,5.4154058,4.759466,4.1035266,3.4514916,3.0141985,2.5769055,2.135708,1.698415,1.261122,1.3509232,1.43682,1.5266213,1.6125181,1.698415,1.8663043,2.0302892,2.194274,2.358259,2.5261483,2.631567,2.7408905,2.8463092,2.9556324,3.0610514,3.3538816,3.6467118,3.9395418,4.2323723,4.5252023,5.3451266,6.165051,6.984976,7.8049,8.624825,10.823003,13.021181,15.21936,17.413633,19.611813,18.475632,17.343355,16.207174,15.070992,13.938716,12.982138,12.029464,11.072885,10.116306,9.163632,8.917655,8.671678,8.4257,8.183627,7.9376497,7.0240197,6.114294,5.2006636,4.2870336,3.3734035,3.3734035,3.3694992,3.3655949,3.3655949,3.3616903,3.1898966,3.018103,2.8463092,2.6706111,2.4988174,2.4207294,2.338737,2.260649,2.1786566,2.1005683,2.8775444,3.6545205,4.4314966,5.2084727,5.989353,7.629202,9.269051,10.9089,12.548749,14.188598,12.825961,11.4633255,10.100689,8.738052,7.375416,6.6531014,5.9346914,5.2162814,4.493967,3.775557,3.4280653,3.084478,2.7408905,2.3933985,2.0498111,2.1239948,2.1981785,2.2762666,2.35045,2.4246337,2.6667068,2.9087796,3.1508527,3.39683,3.638903,3.4046388,3.174279,2.9400148,2.7057507,2.475391,2.4207294,2.366068,2.3114061,2.2567444,2.1981785,1.9248703,1.6515622,1.3743496,1.1010414,0.8238289,3.3460727,5.872221,8.3944645,10.916709,13.438952,12.326198,11.217348,10.108498,8.995743,7.8868923,0.6637484,0.659844,0.6559396,0.6559396,0.6520352,0.6481308,0.6715572,0.6949836,0.71841,0.7418364,0.76135844,0.78088045,0.80430686,0.8238289,0.8433509,0.8628729,0.8628729,0.8628729,0.8628729,0.8628729,0.8628729,0.93705654,1.0112402,1.0893283,1.1635119,1.2376955,1.4875772,1.737459,1.9873407,2.2372224,2.4871042,2.9322062,3.377308,3.8224099,4.267512,4.7126136,4.6384296,4.564246,4.4861584,4.4119744,4.337791,5.181142,6.0205884,6.8639393,7.70729,8.550641,8.898132,9.249529,9.600925,9.948417,10.299813,11.576552,12.849388,14.126127,15.398962,16.675701,16.289165,15.8987255,15.51219,15.125654,14.739119,14.489237,14.243259,13.993378,13.7474,13.501423,10.951848,8.398369,5.8487945,3.2992198,0.74964523,0.80040246,0.8511597,0.9019169,0.94876975,0.999527,1.3001659,1.6008049,1.901444,2.1981785,2.4988174,2.455869,2.4090161,2.366068,2.3192148,2.2762666,2.330928,2.3855898,2.4402514,2.494913,2.5495746,2.2762666,2.0068626,1.7335546,1.4602464,1.1869383,1.1596074,1.1322767,1.1049459,1.077615,1.0502841,3.0141985,4.9742084,6.9381227,8.898132,10.862047,13.477997,16.093946,18.705992,21.321941,23.937891,23.301472,22.668959,22.032541,21.396124,20.76361,19.748466,18.737226,17.725986,16.710842,15.699601,15.430198,15.160794,14.89139,14.618082,14.348679,14.188598,14.028518,13.868437,13.708356,13.548276,13.536563,13.520945,13.505327,13.48971,13.4740925,13.64979,13.825488,14.001186,14.176885,14.348679,13.353056,12.361338,11.365715,10.370092,9.37447,8.710721,8.050878,7.387129,6.7233806,6.0635366,6.3915067,6.7233806,7.0513506,7.3832245,7.7111945,7.4495993,7.1880045,6.9264097,6.66091,6.3993154,6.699954,7.000593,7.3012323,7.601871,7.898606,7.4495993,7.000593,6.551587,6.098676,5.64967,5.3529353,5.056201,4.755562,4.4588275,4.1620927,4.4275923,4.6930914,4.958591,5.22409,5.4856853,5.5169206,5.548156,5.579391,5.606722,5.6379566,5.423215,5.212377,5.001539,4.786797,4.575959,4.40807,4.240181,4.0722914,3.9044023,3.736513,4.0059166,4.279225,4.548629,4.8180323,5.087436,5.083532,5.083532,5.0796275,5.0757227,5.0757227,4.4314966,3.7911747,3.1469483,2.5066261,1.8623998,1.7608855,1.6593709,1.5539521,1.4524376,1.3509232,1.53443,1.7140326,1.8975395,2.0810463,2.260649,2.1435168,2.0224805,1.901444,1.7843118,1.6632754,1.7804074,1.8975395,2.0146716,2.1318035,2.2489357,2.3855898,2.5183394,2.6549935,2.7916477,2.9243972,3.6232853,4.318269,5.017157,5.716045,6.4110284,6.606249,6.7975645,6.98888,7.1841,7.375416,6.551587,5.7238536,4.900025,4.0761957,3.2484627,3.018103,2.7838387,2.5534792,2.3192148,2.0888553,2.3543546,2.6159496,2.8814487,3.1469483,3.4124475,3.5178664,3.6232853,3.7287042,3.8341231,3.9356375,3.8302186,3.7208953,3.6154766,3.506153,3.4007344,4.1464753,4.8883114,5.6340523,6.379793,7.125534,6.8678436,6.610153,6.3524623,6.094772,5.8370814,10.342762,14.848442,19.354122,23.855898,28.361578,24.375183,20.388788,16.398489,12.412095,8.4257,7.266093,6.1103897,4.950782,3.795079,2.639376,2.7213683,2.8072653,2.893162,2.979059,3.0610514,4.5408196,6.016684,7.4964523,8.972317,10.44818,10.096785,9.745388,9.393991,9.0386915,8.687295,8.617016,8.546737,8.476458,8.406178,8.335898,12.142691,15.945579,19.75237,23.559164,27.362051,27.709543,28.057035,28.404526,28.752018,29.09951,28.826202,28.548988,28.27568,27.998468,27.72516,29.290825,30.856491,32.41825,33.983917,35.549583,29.638317,23.730957,17.819693,11.908427,6.001066,5.142098,4.283129,3.4280653,2.5690966,1.7140326,2.3035975,2.8970666,3.4905357,4.084005,4.6735697,4.7907014,4.903929,5.0210614,5.134289,5.251421,6.6687193,8.089922,9.511124,10.928422,12.349625,12.162213,11.974802,11.787391,11.599979,11.412568,11.795199,12.177831,12.560462,12.943093,13.325725,12.849388,12.369146,11.892809,11.416472,10.936231,9.378374,7.824422,6.266566,4.7087092,3.1508527,2.5183394,1.8897307,1.261122,0.62860876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,0.6442264,0.8902037,1.1361811,1.3782539,1.6242313,1.8311646,2.0341935,2.241127,2.4441557,2.6510892,2.5300527,2.4090161,2.2918842,2.1708477,2.0498111,2.0341935,2.018576,2.0068626,1.9912452,1.9756275,2.5808098,3.1898966,3.7989833,4.4041657,5.0132523,4.618908,4.220659,3.8263142,3.4319696,3.0376248,3.0024853,2.9673457,2.9322062,2.8970666,2.8619268,3.521771,4.1777105,4.83365,5.493494,6.1494336,6.461786,6.7702336,7.0786815,7.3910336,7.699481,8.769287,9.835189,10.901091,11.970898,13.036799,13.376482,13.716166,14.055848,14.399435,14.739119,14.098797,13.458474,12.818152,12.177831,11.537509,10.951848,10.366188,9.780528,9.198771,8.6131115,9.190963,9.772718,10.350571,10.932326,11.514082,12.240301,12.96652,13.696643,14.422862,15.14908,14.551707,13.950429,13.349152,12.751778,12.150499,14.126127,16.10566,18.081287,20.06082,22.036446,19.764084,17.487818,15.211552,12.939189,10.662923,9.796145,8.929368,8.058686,7.191909,6.3251314,8.113348,9.905469,11.693685,13.4858055,15.274021,15.410676,15.551234,15.687888,15.824542,15.961197,16.437534,16.91387,17.386303,17.86264,18.338978,22.590872,26.84667,31.102468,35.35827,39.614067,36.959072,34.307983,31.652988,29.0019,26.350811,25.511364,24.668013,23.828568,22.98912,22.149673,18.030529,13.911386,9.788337,5.6691923,1.5500476,1.2415999,0.92924774,0.62079996,0.30844778,0.0,1.7608855,3.521771,5.278752,7.039637,8.800523,9.999174,11.193921,12.392572,13.591225,14.785972,12.564366,10.342762,8.121157,5.8956475,3.6740425,3.154757,2.6354716,2.1161861,1.5969005,1.0737107,2.7643168,4.454923,6.1455293,7.8361354,9.526741,9.733675,9.944512,10.155351,10.366188,10.573121,9.440845,8.304664,7.168483,6.036206,4.900025,4.388548,3.873167,3.3616903,2.8502135,2.338737,2.2762666,2.2137961,2.1513257,2.0888553,2.0263848,2.194274,2.358259,2.5261483,2.6940374,2.8619268,2.9283018,2.9907722,3.057147,3.1235218,3.1859922,3.3226464,3.4593005,3.59205,3.7287042,3.8614538,4.6384296,5.4193106,6.196286,6.9732623,7.7502384,9.557977,11.365715,13.173453,14.981192,16.788929,16.031475,15.274021,14.516567,13.759113,13.001659,12.2793455,11.553126,10.8308115,10.108498,9.386183,9.546264,9.706344,9.866425,10.0265045,10.186585,9.124588,8.062591,7.000593,5.938596,4.8765984,4.970304,5.0640097,5.1616197,5.2553253,5.349031,4.9663997,4.5837684,4.2011366,3.8185053,3.435874,3.2757936,3.1157131,2.9556324,2.7994564,2.639376,3.1781836,3.7208953,4.263607,4.806319,5.349031,6.590631,7.8361354,9.077735,10.319335,11.560935,10.725393,9.885946,9.050405,8.210958,7.375416,6.735094,6.094772,5.45445,4.814128,4.173806,3.8106966,3.4436827,3.0805733,2.7135596,2.35045,2.2996929,2.2489357,2.1981785,2.1513257,2.1005683,2.3465457,2.5964274,2.8424048,3.0883822,3.338264,3.1586614,2.9829633,2.803361,2.6276627,2.4480603,2.541766,2.631567,2.7213683,2.8111696,2.900971,2.5378613,2.174752,1.8116426,1.4485333,1.0893283,3.3460727,5.602817,7.859562,10.116306,12.373051,11.506273,10.6355915,9.76491,8.894228,8.023546,0.6481308,0.6520352,0.6559396,0.6559396,0.659844,0.6637484,0.6910792,0.71841,0.74574083,0.77307165,0.80040246,0.8160201,0.8355421,0.8511597,0.8706817,0.8862993,0.8745861,0.8628729,0.8511597,0.8394465,0.8238289,0.9136301,0.999527,1.0893283,1.175225,1.261122,1.5110037,1.7608855,2.0107672,2.260649,2.514435,2.7916477,3.0727646,3.3538816,3.631094,3.912211,3.900498,3.8887846,3.873167,3.8614538,3.8497405,4.970304,6.0908675,7.211431,8.32809,9.448653,9.86252,10.276386,10.686349,11.100216,11.514082,12.537036,13.563893,14.586847,15.613705,16.636658,16.437534,16.238409,16.039284,15.836256,15.637131,14.399435,13.157836,11.916236,10.67854,9.43694,7.648724,5.8644123,4.0761957,2.2879796,0.4997635,0.6871748,0.8745861,1.0619974,1.2494087,1.43682,1.901444,2.3621633,2.8267872,3.2875066,3.7482262,3.6467118,3.541293,3.435874,3.330455,3.2250361,3.3460727,3.4632049,3.5842414,3.7052777,3.8263142,3.408543,2.9946766,2.5808098,2.1630387,1.7491722,1.5890918,1.4290112,1.2689307,1.1088502,0.94876975,3.2367494,5.5247293,7.812709,10.100689,12.388668,15.683984,18.983204,22.278519,25.57774,28.873055,27.522131,26.171207,24.816381,23.465458,22.11063,20.712854,19.311174,17.913397,16.511717,15.113941,14.79378,14.477524,14.161267,13.841106,13.524849,13.497519,13.470188,13.442857,13.415526,13.388195,13.403813,13.419431,13.431144,13.446761,13.462379,13.388195,13.314012,13.235924,13.16174,13.087557,12.2559185,11.428185,10.596548,9.768814,8.937177,8.476458,8.011833,7.551114,7.08649,6.6257706,6.7702336,6.914696,7.0591593,7.2036223,7.348085,7.250475,7.1489606,7.0513506,6.949836,6.8483214,7.113821,7.375416,7.6370106,7.898606,8.164105,7.7385254,7.3129454,6.8873653,6.461786,6.036206,5.661383,5.282656,4.903929,4.5291066,4.1503797,4.423688,4.6930914,4.9663997,5.239708,5.5130157,5.7316628,5.9542136,6.17286,6.3915067,6.6140575,6.3251314,6.036206,5.7511845,5.462259,5.173333,4.9156423,4.661856,4.4041657,4.1464753,3.8887846,4.041056,4.1972322,4.3534083,4.50568,4.661856,4.6540475,4.6423345,4.630621,4.6228123,4.6110992,4.029343,3.4475873,2.8658314,2.2840753,1.698415,1.7257458,1.7530766,1.7843118,1.8116426,1.8389735,2.0810463,2.3231194,2.5651922,2.8072653,3.049338,2.7682211,2.4910088,2.2098918,1.9287747,1.6515622,1.796025,1.9404879,2.084951,2.2294137,2.3738766,2.514435,2.6549935,2.795552,2.9361105,3.076669,3.8263142,4.579864,5.3334136,6.083059,6.8366084,7.0201154,7.2036223,7.3832245,7.5667315,7.7502384,6.9615493,6.1767645,5.388075,4.5993857,3.8106966,3.5451972,3.2757936,3.0102942,2.7408905,2.475391,2.7604125,3.0454338,3.330455,3.6154766,3.900498,3.8965936,3.8887846,3.8848803,3.8809757,3.873167,3.7560349,3.638903,3.521771,3.4046388,3.2875066,3.9161155,4.548629,5.1772375,5.805846,6.4383593,6.2197127,6.001066,5.786324,5.5676775,5.349031,9.63216,13.91529,18.19842,22.481548,26.760773,23.160913,19.561056,15.961197,12.361338,8.761478,7.5433054,6.329036,5.1108627,3.892689,2.6745155,2.5651922,2.455869,2.3465457,2.233318,2.1239948,3.2992198,4.4705405,5.6418614,6.813182,7.988407,7.9766936,7.968885,7.957172,7.9493628,7.9376497,7.9337454,7.9259367,7.9220324,7.918128,7.914223,11.268105,14.625891,17.983677,21.341463,24.69925,25.741724,26.780294,27.818867,28.861341,29.899912,29.888199,29.876486,29.860868,29.849155,29.837442,31.871635,33.90583,35.943928,37.97812,40.012314,33.370926,26.733442,20.092054,13.450665,6.813182,5.9073606,5.001539,4.095718,3.193801,2.2879796,3.232845,4.1777105,5.1225758,6.067441,7.012306,7.1841,7.355894,7.531592,7.703386,7.8751793,9.20658,10.534078,11.8654785,13.196879,14.524376,14.649317,14.774258,14.899199,15.024139,15.14908,14.95386,14.75864,14.56342,14.3682,14.176885,13.216402,12.2559185,11.295436,10.334952,9.37447,7.918128,6.46569,5.009348,3.5569105,2.1005683,1.678893,1.261122,0.8394465,0.42167544,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12103647,0.23816854,0.359205,0.48024148,0.60127795,0.96829176,1.3353056,1.7023194,2.069333,2.436347,2.3933985,2.3543546,2.3114061,2.2684577,2.2255092,2.1435168,2.0654287,1.9834363,1.9053483,1.8233559,1.7413634,1.6554666,1.5695697,1.4836729,1.4016805,1.9443923,2.4831998,3.0259118,3.5686235,4.1113358,3.8067923,3.5022488,3.1977055,2.893162,2.5886188,2.5847144,2.5808098,2.5808098,2.5769055,2.5769055,3.4046388,4.2362766,5.0640097,5.8956475,6.7233806,7.016211,7.3051367,7.5940623,7.8868923,8.175818,9.343235,10.514555,11.685876,12.853292,14.024612,13.7474,13.470188,13.192975,12.915763,12.63855,12.041177,11.443803,10.84643,10.249056,9.651682,9.358852,9.069926,8.781001,8.488171,8.1992445,8.531119,8.866898,9.198771,9.530646,9.86252,10.573121,11.283723,11.994324,12.70102,13.411622,13.173453,12.939189,12.70102,12.4628525,12.224684,14.11051,15.996336,17.878258,19.764084,21.64991,20.51373,19.373644,18.237463,17.101282,15.961197,13.794253,11.623405,9.452558,7.28171,5.1108627,7.8478484,10.58093,13.317916,16.050997,18.787983,18.276506,17.761126,17.24965,16.738173,16.226696,16.250122,16.273548,16.300879,16.324306,16.351637,21.958359,27.56508,33.171803,38.778522,44.38915,39.10259,33.81603,28.533371,23.24681,17.964155,17.327738,16.69132,16.058807,15.422389,14.785972,12.107552,9.4291315,6.746807,4.068387,1.3860629,1.1088502,0.8316377,0.5544251,0.27721256,0.0,2.4519646,4.903929,7.355894,9.811763,12.263727,12.025558,11.791295,11.557031,11.322766,11.088503,9.358852,7.633106,5.903456,4.1777105,2.4480603,2.2840753,2.1161861,1.9482968,1.7804074,1.6125181,3.4593005,5.3060827,7.1567693,9.0035515,10.850334,11.564839,12.2793455,12.993851,13.708356,14.426766,12.810344,11.193921,9.581403,7.9649806,6.348558,5.7628975,5.173333,4.5876727,3.998108,3.4124475,3.2016098,2.9868677,2.77603,2.5612879,2.35045,2.5183394,2.690133,2.8619268,3.0298162,3.2016098,3.2211318,3.2445583,3.2679846,3.2914112,3.310933,3.2914112,3.2679846,3.2445583,3.2211318,3.2016098,3.9356375,4.6696653,5.4036927,6.141625,6.8756523,8.292951,9.710248,11.127546,12.544845,13.962143,13.583415,13.200784,12.822057,12.44333,12.0606985,11.572648,11.080693,10.592644,10.100689,9.612638,10.178777,10.741011,11.307149,11.873287,12.439425,11.225157,10.010887,8.800523,7.5862536,6.375889,6.5672045,6.75852,6.9537406,7.1450562,7.336372,6.746807,6.153338,5.559869,4.9663997,4.376835,4.134762,3.8965936,3.6545205,3.416352,3.174279,3.4827268,3.7911747,4.095718,4.4041657,4.7126136,5.5559645,6.4032197,7.2465706,8.093826,8.937177,8.624825,8.312472,8.00012,7.687768,7.375416,6.813182,6.2548523,5.6965227,5.134289,4.575959,4.1894236,3.8067923,3.4202564,3.0337205,2.6510892,2.475391,2.2996929,2.1239948,1.9482968,1.7765031,2.0263848,2.280171,2.533957,2.7838387,3.0376248,2.9165885,2.7916477,2.6706111,2.5456703,2.4246337,2.6588979,2.893162,3.1313305,3.3655949,3.5998588,3.1508527,2.7018464,2.2489357,1.7999294,1.3509232,3.3421683,5.3334136,7.328563,9.319808,11.311053,10.682445,10.053836,9.421323,8.792714,8.164105,0.63641757,0.6442264,0.6520352,0.659844,0.6676528,0.6754616,0.7066968,0.7418364,0.77307165,0.80430686,0.8394465,0.8511597,0.8667773,0.8823949,0.8980125,0.9136301,0.8862993,0.8628729,0.8394465,0.81211567,0.78868926,0.8862993,0.9878138,1.0893283,1.1869383,1.2884527,1.5383345,1.7882162,2.0380979,2.2879796,2.5378613,2.6510892,2.7682211,2.8814487,2.998581,3.1118085,3.1625657,3.213323,3.2640803,3.310933,3.3616903,4.759466,6.1572423,7.5550184,8.952794,10.350571,10.826907,11.29934,11.775677,12.24811,12.724447,13.501423,14.274494,15.051471,15.824542,16.601519,16.585901,16.574188,16.562475,16.55076,16.539047,14.30573,12.072412,9.839094,7.605776,5.376362,4.349504,3.3265507,2.2996929,1.2767396,0.24988174,0.57394713,0.9019169,1.2259823,1.5500476,1.8741131,2.4988174,3.1235218,3.7482262,4.376835,5.001539,4.83365,4.6696653,4.50568,4.3416953,4.173806,4.3612175,4.5447245,4.728231,4.9156423,5.099149,4.5408196,3.9863946,3.4280653,2.8697357,2.3114061,2.018576,1.7257458,1.43682,1.1439898,0.8511597,3.4632049,6.0752497,8.687295,11.29934,13.911386,17.893875,21.872461,25.851048,29.833538,33.812122,31.74279,29.673458,27.604124,25.530886,23.461554,21.673336,19.889025,18.10081,16.312593,14.524376,14.161267,13.794253,13.431144,13.06413,12.70102,12.806439,12.911859,13.013372,13.118792,13.224211,13.271063,13.314012,13.360865,13.403813,13.450665,13.1266,12.798631,12.4745655,12.150499,11.826434,11.158782,10.495033,9.8312845,9.163632,8.499884,8.238289,7.9766936,7.7111945,7.4495993,7.1880045,7.1489606,7.1060123,7.066968,7.027924,6.98888,7.0513506,7.113821,7.1762915,7.238762,7.3012323,7.523783,7.7502384,7.9766936,8.1992445,8.4257,8.023546,7.6252975,7.223144,6.824895,6.426646,5.9659266,5.5091114,5.0522966,4.5954814,4.138666,4.415879,4.6969957,4.9781127,5.2592297,5.5364423,5.9464045,6.356367,6.7663293,7.1762915,7.5862536,7.223144,6.8639393,6.5008297,6.13772,5.774611,5.4271193,5.0796275,4.732136,4.3846436,4.037152,4.0761957,4.1191444,4.1581883,4.1972322,4.2362766,4.220659,4.2011366,4.185519,4.165997,4.1503797,3.6271896,3.1039999,2.5808098,2.0615244,1.5383345,1.6945106,1.8506867,2.0107672,2.1669433,2.3231194,2.6276627,2.9283018,3.232845,3.533484,3.8380275,3.39683,2.9556324,2.5183394,2.077142,1.6359446,1.8116426,1.9834363,2.15523,2.3270237,2.4988174,2.6432803,2.7916477,2.9361105,3.0805733,3.2250361,4.0332475,4.841459,5.645766,6.453977,7.262188,7.433982,7.605776,7.7814736,7.9532676,8.125061,7.375416,6.6257706,5.8761253,5.12648,4.376835,4.0722914,3.7716527,3.4671092,3.1664703,2.8619268,3.1664703,3.4710135,3.7794614,4.084005,4.388548,4.271416,4.1581883,4.041056,3.9278288,3.8106966,3.6857557,3.5569105,3.4280653,3.3031244,3.174279,3.68966,4.2050414,4.7204223,5.2358036,5.7511845,5.571582,5.395884,5.2162814,5.040583,4.860981,8.921559,12.982138,17.042715,21.103294,25.163872,21.95055,18.737226,15.523903,12.31058,9.101162,7.824422,6.5437784,5.267039,3.9902992,2.7135596,2.4090161,2.1005683,1.796025,1.4914817,1.1869383,2.0537157,2.9243972,3.7911747,4.657952,5.5247293,5.8566036,6.1884775,6.524256,6.8561306,7.1880045,7.2465706,7.309041,7.367607,7.426173,7.4886436,10.397423,13.306203,16.218887,19.127666,22.036446,23.77,25.503555,27.233206,28.96676,30.700315,30.950197,31.200079,31.44996,31.699842,31.949724,34.45635,36.959072,39.4657,41.96842,44.475044,37.103535,29.735928,22.364416,14.996809,7.6252975,6.6726236,5.7199492,4.7672753,3.814601,2.8619268,4.1581883,5.4583545,6.754616,8.050878,9.351044,9.581403,9.811763,10.0382185,10.268578,10.498938,11.740538,12.978233,14.219833,15.461433,16.69913,17.136421,17.573715,18.011007,18.448301,18.889498,18.116426,17.343355,16.570284,15.797212,15.024139,13.583415,12.138786,10.698062,9.253433,7.812709,6.461786,5.1069584,3.7560349,2.4012074,1.0502841,0.8394465,0.62860876,0.42167544,0.21083772,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16008049,0.32016098,0.48024148,0.64032197,0.80040246,1.2884527,1.7804074,2.2684577,2.7604125,3.2484627,2.959537,2.6706111,2.3816853,2.0888553,1.7999294,1.7608855,1.7218413,1.678893,1.639849,1.6008049,1.4446288,1.2884527,1.1361811,0.98000497,0.8238289,1.3040704,1.7804074,2.2567444,2.7330816,3.213323,2.998581,2.7838387,2.5690966,2.3543546,2.135708,2.1669433,2.1981785,2.2294137,2.2567444,2.2879796,3.2914112,4.290938,5.2943697,6.297801,7.3012323,7.570636,7.8400397,8.109444,8.378847,8.648251,9.921086,11.193921,12.466757,13.739592,15.012426,14.118319,13.224211,12.326198,11.43209,10.537982,9.983557,9.4291315,8.870802,8.316377,7.7619514,7.7658563,7.773665,7.7775693,7.7814736,7.7892823,7.871275,7.957172,8.043069,8.128965,8.210958,8.905942,9.597021,10.2881,10.983084,11.674163,11.799104,11.924045,12.0489855,12.173926,12.298867,14.090988,15.883108,17.679134,19.471254,21.263374,21.263374,21.263374,21.263374,21.263374,21.263374,17.788456,14.317443,10.84643,7.3715115,3.900498,7.578445,11.260296,14.938243,18.620094,22.301945,21.138433,19.974922,18.81141,17.651802,16.48829,16.062712,15.637131,15.211552,14.785972,14.364296,21.321941,28.28349,35.241135,42.202682,49.164234,41.246105,33.327976,25.40985,17.491722,9.573594,9.14411,8.714626,8.285142,7.8556576,7.426173,6.184573,4.9468775,3.7052777,2.463678,1.2259823,0.98000497,0.7340276,0.48805028,0.24597734,0.0,3.1469483,6.289992,9.43694,12.579984,15.726933,14.055848,12.388668,10.721489,9.054309,7.387129,6.153338,4.9234514,3.68966,2.455869,1.2259823,1.4094892,1.5969005,1.7804074,1.9639144,2.1513257,4.154284,6.1611466,8.164105,10.170968,12.173926,13.396004,14.614178,15.836256,17.054428,18.276506,16.179844,14.0831785,11.990419,9.893755,7.800996,7.137247,6.473499,5.813655,5.1499066,4.4861584,4.123049,3.7638438,3.4007344,3.0376248,2.6745155,2.8463092,3.018103,3.193801,3.3655949,3.5373883,3.5178664,3.4983444,3.4788225,3.4593005,3.435874,3.2562714,3.076669,2.8970666,2.717464,2.5378613,3.2289407,3.9239242,4.6150036,5.3060827,6.001066,7.027924,8.054782,9.081639,10.108498,11.139259,11.135355,11.131451,11.131451,11.127546,11.123642,10.865952,10.608261,10.350571,10.096785,9.839094,10.807385,11.775677,12.747873,13.716166,14.688361,13.325725,11.963089,10.600452,9.237816,7.8751793,8.164105,8.456935,8.745861,9.034787,9.323712,8.52331,7.719003,6.918601,6.114294,5.3138914,4.9937305,4.6735697,4.3534083,4.0332475,3.7130866,3.7833657,3.8575494,3.9317331,4.0020123,4.0761957,4.521298,4.970304,5.4193106,5.8644123,6.3134184,6.524256,6.7389984,6.949836,7.1606736,7.375416,6.8951745,6.4149327,5.9346914,5.45445,4.9742084,4.5681505,4.165997,3.7599394,3.3538816,2.951728,2.6510892,2.35045,2.0498111,1.7491722,1.4485333,1.7062237,1.9639144,2.2216048,2.4792955,2.736986,2.6706111,2.6042364,2.533957,2.4675822,2.4012074,2.7799344,3.1586614,3.541293,3.9200199,4.298747,3.7638438,3.2250361,2.6862288,2.1513257,1.6125181,3.338264,5.067914,6.79366,8.52331,10.249056,9.858616,9.468176,9.081639,8.691199,8.300759,0.62470436,0.63641757,0.6481308,0.6637484,0.6754616,0.6871748,0.7262188,0.76135844,0.80040246,0.8394465,0.8745861,0.8862993,0.9019169,0.9136301,0.92534333,0.93705654,0.9019169,0.8628729,0.8238289,0.78868926,0.74964523,0.8628729,0.97610056,1.0893283,1.1986516,1.3118792,1.5617609,1.8116426,2.0615244,2.3114061,2.5612879,2.514435,2.463678,2.4129205,2.3621633,2.3114061,2.4246337,2.5378613,2.6510892,2.7643168,2.87364,4.548629,6.223617,7.898606,9.573594,11.248583,11.787391,12.326198,12.861101,13.399908,13.938716,14.461906,14.989,15.51219,16.039284,16.562475,16.738173,16.91387,17.085665,17.261362,17.437061,14.212025,10.986988,7.7619514,4.5369153,1.3118792,1.0502841,0.78868926,0.5231899,0.26159495,0.0,0.46071947,0.92534333,1.3860629,1.8506867,2.3114061,3.1000953,3.8887846,4.6735697,5.462259,6.250948,6.0244927,5.801942,5.575486,5.349031,5.12648,5.376362,5.6262436,5.8761253,6.126007,6.375889,5.6730967,4.9742084,4.2753205,3.5764325,2.87364,2.4480603,2.0263848,1.6008049,1.175225,0.74964523,3.6857557,6.6257706,9.561881,12.501896,15.438006,20.099863,24.761719,29.423576,34.089336,38.751194,35.963448,33.175705,30.387962,27.60022,24.812477,22.637724,20.462973,18.28822,16.113468,13.938716,13.524849,13.110983,12.70102,12.287154,11.873287,12.111456,12.349625,12.587793,12.825961,13.06413,13.138313,13.212498,13.286681,13.360865,13.438952,12.861101,12.287154,11.713207,11.139259,10.561408,10.061645,9.561881,9.062118,8.562354,8.062591,8.00012,7.9376497,7.8751793,7.812709,7.7502384,7.523783,7.3012323,7.0747766,6.8483214,6.6257706,6.8483214,7.0747766,7.3012323,7.523783,7.7502384,7.9376497,8.125061,8.312472,8.499884,8.687295,8.312472,7.9376497,7.562827,7.1880045,6.813182,6.2743745,5.735567,5.2006636,4.661856,4.123049,4.4119744,4.7009,4.985922,5.2748475,5.563773,6.1611466,6.7624245,7.363703,7.9610763,8.562354,8.125061,7.687768,7.250475,6.813182,6.375889,5.938596,5.5013027,5.0640097,4.6267166,4.1894236,4.1113358,4.037152,3.9629683,3.8887846,3.8106966,3.78727,3.7638438,3.736513,3.7130866,3.6857557,3.2250361,2.7643168,2.2996929,1.8389735,1.3743496,1.6632754,1.9482968,2.2372224,2.5261483,2.8111696,3.174279,3.5373883,3.900498,4.263607,4.6267166,4.025439,3.4241607,2.8267872,2.2255092,1.6242313,1.8233559,2.0263848,2.2255092,2.4246337,2.6237583,2.77603,2.9243972,3.076669,3.2250361,3.3734035,4.2362766,5.099149,5.9620223,6.824895,7.687768,7.8517528,8.011833,8.175818,8.335898,8.499884,7.7892823,7.0747766,6.364176,5.64967,4.939069,4.5993857,4.263607,3.9239242,3.5881457,3.2484627,3.5764325,3.900498,4.224563,4.548629,4.8765984,4.650143,4.423688,4.2011366,3.9746814,3.7482262,3.611572,3.474918,3.338264,3.2016098,3.0610514,3.4632049,3.8614538,4.263607,4.661856,5.0640097,4.9234514,4.786797,4.650143,4.513489,4.376835,8.210958,12.0489855,15.8870125,5052.0,23.563068,20.73628,17.913397,15.086611,12.263727,9.43694,8.101635,6.7624245,5.423215,4.087909,2.7486992,2.2489357,1.7491722,1.2494087,0.74964523,0.24988174,0.81211567,1.3743496,1.9365835,2.4988174,3.0610514,3.736513,4.4119744,5.087436,5.7628975,6.4383593,6.5633,6.688241,6.813182,6.9381227,7.0630636,9.526741,11.986515,14.450192,16.91387,19.373644,21.798277,24.226816,26.65145,29.076084,31.500717,32.012196,32.52367,33.03905,33.55053,34.062004,37.03716,40.012314,42.98747,45.962624,48.93778,40.836143,32.738415,24.636778,16.539047,8.437413,7.437886,6.4383593,5.4388323,4.4393053,3.435874,5.087436,6.7389984,8.386656,10.0382185,11.685876,11.974802,12.263727,12.548749,12.837675,13.1266,14.274494,15.426293,16.574188,17.725986,18.87388,19.623526,20.37317,21.12672,21.876366,22.62601,21.275087,19.924164,18.573242,17.226223,15.875299,13.950429,12.025558,10.100689,8.175818,6.250948,5.001539,3.7482262,2.4988174,1.2494087,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19912452,0.39824903,0.60127795,0.80040246,0.999527,1.6125181,2.2255092,2.8385005,3.4514916,4.0605783,3.5256753,2.9868677,2.4480603,1.9131571,1.3743496,1.3743496,1.3743496,1.3743496,1.3743496,1.3743496,1.1517987,0.92534333,0.698888,0.47633708,0.24988174,0.6637484,1.0737107,1.4875772,1.901444,2.3114061,2.1864653,2.0615244,1.9365835,1.8116426,1.6867018,1.7491722,1.8116426,1.8741131,1.9365835,1.999054,3.174279,4.349504,5.5247293,6.699954,7.8751793,8.125061,8.374943,8.624825,8.874706,9.124588,10.498938,11.873287,13.251541,14.625891,16.00024,14.489237,12.974329,11.4633255,9.948417,8.437413,7.9259367,7.4144597,6.899079,6.387602,5.8761253,6.1767645,6.473499,6.774138,7.0747766,7.375416,7.211431,7.0513506,6.8873653,6.7233806,6.5633,7.238762,7.914223,8.58578,9.261242,9.936704,10.424754,10.912805,11.400854,11.888905,12.373051,14.07537,15.773785,17.476105,19.174519,20.876839,22.01302,23.1492,24.289286,25.425468,26.56165,21.786564,17.01148,12.236397,7.461313,2.6862288,7.3129454,11.935758,16.562475,21.189192,25.812004,24.00036,22.188719,20.37317,18.56153,16.749886,15.875299,15.000713,14.126127,13.251541,12.373051,20.689428,28.997995,37.314373,45.626846,53.939316,43.38572,32.83602,22.286327,11.736633,1.1869383,0.96438736,0.737932,0.5114767,0.28892577,0.062470436,0.26159495,0.46071947,0.6637484,0.8628729,1.0619974,0.8511597,0.63641757,0.42557985,0.21083772,0.0,3.8380275,7.676055,11.514082,15.348206,19.186234,16.086138,12.986042,9.885946,6.785851,3.6857557,2.951728,2.2137961,1.475864,0.737932,0.0,0.5388075,1.0737107,1.6125181,2.1513257,2.6862288,4.8492675,7.012306,9.175345,11.338385,13.501423,15.223265,16.94901,18.674755,20.400501,22.126247,19.549341,16.976341,14.399435,11.826434,9.249529,8.511597,7.773665,7.0357327,6.3017054,5.563773,5.0483923,4.5369153,4.025439,3.513962,2.998581,3.174279,3.349977,3.5256753,3.7013733,3.873167,3.8106966,3.7482262,3.6857557,3.6232853,3.5608149,3.2250361,2.8892577,2.5495746,2.2137961,1.8741131,2.5261483,3.174279,3.8263142,4.474445,5.12648,5.7628975,6.3993154,7.0357327,7.676055,8.312472,8.687295,9.062118,9.43694,9.811763,10.186585,10.163159,10.135828,10.112402,10.088976,10.061645,11.435994,12.814248,14.188598,15.562947,16.937298,15.426293,13.911386,12.400381,10.889378,9.37447,9.761005,10.151445,10.537982,10.924518,11.311053,10.299813,9.288573,8.273428,7.262188,6.250948,5.8487945,5.4505453,5.0483923,4.650143,4.251894,4.087909,3.9239242,3.7638438,3.5998588,3.435874,3.4866312,3.5373883,3.5881457,3.638903,3.6857557,4.423688,5.1616197,5.899552,6.6374836,7.375416,6.9732623,6.575013,6.1767645,5.774611,5.376362,4.950782,4.5252023,4.0996222,3.6740425,3.2484627,2.8267872,2.4012074,1.9756275,1.5500476,1.1244678,1.3860629,1.6515622,1.9131571,2.174752,2.436347,2.4246337,2.4129205,2.4012074,2.3855898,2.3738766,2.900971,3.4241607,3.951255,4.474445,5.001539,4.376835,3.7482262,3.1235218,2.4988174,1.8741131,3.338264,4.7985106,6.262661,7.726812,9.187058,9.0386915,8.886419,8.738052,8.58578,8.437413,0.6637484,0.6715572,0.6832704,0.6910792,0.7027924,0.7106012,0.74964523,0.78868926,0.8238289,0.8628729,0.9019169,0.9058213,0.9136301,0.92143893,0.92924774,0.93705654,0.9058213,0.8784905,0.8472553,0.8160201,0.78868926,0.8784905,0.97219616,1.0659018,1.1557031,1.2494087,1.4524376,1.6554666,1.8584955,2.0615244,2.260649,2.2450314,2.2294137,2.2098918,2.194274,2.174752,2.4714866,2.7643168,3.0610514,3.3538816,3.6506162,5.0718184,6.4891167,7.910319,9.331521,10.748819,11.447707,12.146595,12.841579,13.540467,14.239355,15.008522,15.781594,16.554665,17.327738,18.10081,17.679134,17.253553,16.831879,16.410202,15.988527,13.196879,10.401327,7.60968,4.8180323,2.0263848,1.620327,1.2142692,0.80821127,0.40605783,0.0,0.3709182,0.7418364,1.1088502,1.4797685,1.8506867,2.4792955,3.1118085,3.7404175,4.369026,5.001539,4.8219366,4.6384296,4.4588275,4.279225,4.0996222,4.3065557,4.513489,4.7243266,4.93126,5.138193,4.6110992,4.084005,3.5569105,3.0259118,2.4988174,2.1786566,1.8545911,1.53443,1.2103647,0.8862993,3.240654,5.5989127,7.9532676,10.307622,12.661977,16.32821,19.998348,23.664581,27.330816,31.000954,28.947239,26.893522,24.843712,22.789995,20.73628,19.217468,17.698656,16.175938,14.657126,13.138313,12.681499,12.220779,11.763964,11.307149,10.850334,10.951848,11.053363,11.158782,11.260296,11.361811,11.369619,11.377428,11.385237,11.393045,11.400854,10.971371,10.545791,10.116306,9.690726,9.261242,8.94889,8.632633,8.316377,8.0040245,7.687768,7.6448197,7.601871,7.558923,7.5159745,7.47693,7.266093,7.0591593,6.852226,6.6452928,6.4383593,6.7233806,7.012306,7.3012323,7.5862536,7.8751793,8.101635,8.32809,8.55845,8.784905,9.01136,8.702912,8.39056,8.082112,7.773665,7.461313,6.860035,6.2587566,5.6535745,5.0522966,4.4510183,4.6423345,4.83365,5.02887,5.2201858,5.4115014,5.8956475,6.3836975,6.8678436,7.3519893,7.8361354,7.590158,7.3441806,7.094299,6.8483214,6.5984397,6.297801,5.9932575,5.6926184,5.388075,5.087436,4.8961205,4.7009,4.5095844,4.318269,4.126953,3.9942036,3.8614538,3.7287042,3.5959544,3.4632049,3.1391394,2.8111696,2.4871042,2.1630387,1.8389735,2.1005683,2.3621633,2.6237583,2.8892577,3.1508527,3.5373883,3.9239242,4.3143644,4.7009,5.087436,4.6540475,4.220659,3.7911747,3.357786,2.9243972,2.8619268,2.795552,2.7291772,2.6667068,2.6003318,2.7721257,2.9439192,3.1157131,3.2914112,3.4632049,4.2167544,4.9742084,5.727758,6.481308,7.238762,7.3441806,7.453504,7.558923,7.6682463,7.773665,7.1216297,6.46569,5.8097506,5.153811,4.5017757,4.2440853,3.9863946,3.7287042,3.4710135,3.213323,3.5998588,3.9863946,4.376835,4.7633705,5.1499066,4.884407,4.618908,4.3534083,4.0918136,3.8263142,3.7287042,3.6349986,3.541293,3.4436827,3.349977,3.697469,4.044961,4.3924527,4.7399445,5.087436,4.892216,4.6969957,4.5017757,4.3065557,4.1113358,7.918128,11.728825,15.535617,19.34241,23.1492,20.599627,18.05005,15.500477,12.950902,10.401327,8.929368,7.461313,5.989353,4.521298,3.049338,2.4831998,1.9209659,1.3548276,0.78868926,0.22645533,0.79649806,1.3665408,1.9365835,2.5066261,3.076669,3.959064,4.841459,5.7238536,6.606249,7.4886436,7.562827,7.6370106,7.7111945,7.7892823,7.8634663,9.63216,11.400854,13.173453,14.942147,16.710842,19.518106,22.321468,25.128733,27.932095,30.739359,31.606136,32.47291,33.33969,34.206467,35.073246,36.55692,38.040592,39.524265,41.004032,42.487705,35.596436,28.70907,21.8178,14.92653,8.039165,6.996689,5.958118,4.9156423,3.8770714,2.8385005,4.4432096,6.0518236,7.660437,9.269051,10.87376,11.365715,11.861574,12.353529,12.845484,13.337439,14.2666855,15.192029,16.121277,17.04662,17.975868,18.90121,19.83046,20.755802,21.685051,22.614298,21.368793,20.12329,18.877785,17.63228,16.386776,14.11051,11.834243,9.554072,7.277806,5.001539,4.123049,3.2484627,2.3738766,1.4992905,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.0,0.0,0.0,0.0,0.0,0.0,0.07027924,0.14055848,0.21083772,0.28111696,0.3513962,0.57394713,0.79649806,1.0190489,1.2415999,1.4641509,1.9561055,2.4519646,2.9478238,3.4436827,3.9356375,3.7482262,3.5608149,3.3734035,3.1859922,2.998581,3.0532427,3.1039999,3.1586614,3.2094188,3.2640803,2.77603,2.2918842,1.8077383,1.3235924,0.8394465,1.2064602,1.5773785,1.9482968,2.3192148,2.6862288,2.4246337,2.1630387,1.901444,1.6359446,1.3743496,1.4914817,1.6047094,1.7218413,1.8350691,1.9482968,2.951728,3.951255,4.950782,5.950309,6.949836,7.480835,8.015738,8.546737,9.081639,9.612638,10.38571,11.158782,11.931853,12.70102,13.4740925,12.318389,11.166591,10.010887,8.855185,7.699481,7.4144597,7.1294384,6.844417,6.559396,6.2743745,6.36808,6.461786,6.551587,6.6452928,6.7389984,6.79366,6.8483214,6.902983,6.957645,7.012306,7.676055,8.343708,9.007456,9.671205,10.338858,11.131451,11.927949,12.724447,13.51704,14.313539,15.933866,17.558098,19.178425,20.802654,22.426888,23.110157,23.793427,24.480602,25.163872,25.851048,21.12672,16.406298,11.681972,6.9615493,2.2372224,6.4695945,10.698062,14.92653,19.158901,23.38737,22.469835,21.5523,20.634766,19.717232,18.799696,17.655706,16.511717,15.363823,14.219833,13.075843,21.458595,29.841347,38.2241,46.60685,54.9857,44.21345,33.4373,22.66115,11.888905,1.1127546,0.9136301,0.71841,0.5192855,0.3240654,0.12494087,1.3157835,2.5105307,3.7013733,4.8961205,6.086963,5.5403466,4.9937305,4.4432096,3.8965936,3.349977,7.859562,12.369146,16.87873,21.388315,25.901804,22.969599,20.041296,17.10909,14.180789,11.248583,9.390087,7.531592,5.6691923,3.8106966,1.9482968,2.3075018,2.6667068,3.0220075,3.3812122,3.736513,5.708236,7.676055,9.647778,11.615597,13.58732,15.320874,17.058334,18.791887,20.529346,22.262901,20.006157,17.749413,15.488764,13.232019,10.975275,10.018696,9.058213,8.101635,7.1450562,6.1884775,5.801942,5.4193106,5.0327744,4.646239,4.263607,4.283129,4.3065557,4.3299823,4.3534083,4.376835,4.3260775,4.2753205,4.224563,4.173806,4.126953,3.7833657,3.4397783,3.096191,2.7565079,2.4129205,2.9634414,3.513962,4.0605783,4.6110992,5.1616197,5.958118,6.7507114,7.5472097,8.343708,9.136301,9.491602,9.8429985,10.194394,10.545791,10.901091,10.9089,10.920613,10.928422,10.940135,10.951848,12.0489855,13.150026,14.251068,15.348206,16.449247,15.375536,14.301826,13.224211,12.150499,11.076789,11.354002,11.631214,11.908427,12.185639,12.4628525,11.572648,10.682445,9.792241,8.902037,8.011833,7.6448197,7.277806,6.910792,6.5437784,6.1767645,6.1221027,6.0713453,6.016684,5.9659266,5.911265,6.0635366,6.2158084,6.36808,6.524256,6.676528,6.9810715,7.289519,7.5979667,7.9064145,8.210958,7.648724,7.082586,6.5164475,5.9542136,5.388075,5.0210614,4.657952,4.290938,3.9278288,3.5608149,3.193801,2.822883,2.4519646,2.0810463,1.7140326,1.8194515,1.9209659,2.0263848,2.1318035,2.2372224,2.3192148,2.4012074,2.4831998,2.5690966,2.6510892,3.049338,3.4436827,3.8419318,4.240181,4.6384296,4.087909,3.5373883,2.9868677,2.436347,1.8858263,3.338264,4.786797,6.239235,7.687768,9.136301,9.073831,9.01136,8.94889,8.886419,8.823949,0.698888,0.7066968,0.7145056,0.7223144,0.7301232,0.737932,0.77307165,0.81211567,0.8511597,0.8862993,0.92534333,0.92924774,0.92924774,0.93315214,0.93315214,0.93705654,0.9136301,0.8941081,0.8706817,0.8472553,0.8238289,0.8980125,0.96829176,1.0424755,1.116659,1.1869383,1.3431144,1.4992905,1.6515622,1.8077383,1.9639144,1.9756275,1.9912452,2.0068626,2.0224805,2.0380979,2.514435,2.9907722,3.4710135,3.9473507,4.423688,5.591104,6.754616,7.918128,9.085544,10.249056,11.108025,11.963089,12.822057,13.6810255,14.53609,15.559043,16.578093,17.597141,18.61619,19.639143,18.61619,17.597141,16.578093,15.559043,14.53609,12.177831,9.815667,7.4574084,5.099149,2.736986,2.1903696,1.6437533,1.0932326,0.5466163,0.0,0.27721256,0.5544251,0.8316377,1.1088502,1.3860629,1.8584955,2.330928,2.803361,3.2757936,3.7482262,3.6154766,3.4788225,3.3460727,3.2094188,3.076669,3.240654,3.4046388,3.5686235,3.736513,3.900498,3.5451972,3.1898966,2.8345962,2.4792955,2.1239948,1.9053483,1.6867018,1.4641509,1.2455044,1.0268579,2.795552,4.5681505,6.3407493,8.113348,9.885946,12.560462,15.231073,17.905588,20.5762,23.250715,21.931028,20.615244,19.295555,17.979773,16.663988,15.797212,14.934339,14.067561,13.200784,12.337912,11.834243,11.330575,10.8308115,10.327144,9.823476,9.792241,9.761005,9.725866,9.694631,9.663396,9.600925,9.542359,9.483793,9.421323,9.362757,9.081639,8.804427,8.52331,8.242193,7.9610763,7.832231,7.703386,7.570636,7.4417906,7.3129454,7.289519,7.266093,7.2465706,7.223144,7.1997175,7.008402,6.8209906,6.629675,6.4383593,6.250948,6.5984397,6.949836,7.3012323,7.648724,8.00012,8.265619,8.535024,8.804427,9.069926,9.339331,9.093353,8.847376,8.601398,8.359325,8.113348,7.445695,6.7780423,6.1103897,5.4427366,4.775084,4.872694,4.970304,5.067914,5.165524,5.263134,5.6340523,6.001066,6.3719845,6.7429028,7.113821,7.055255,6.996689,6.9381227,6.883461,6.824895,6.657006,6.4891167,6.321227,6.153338,5.989353,5.677001,5.368553,5.056201,4.747753,4.4393053,4.1972322,3.959064,3.716991,3.4788225,3.2367494,3.049338,2.8619268,2.6745155,2.4871042,2.2996929,2.5378613,2.77603,3.0141985,3.2484627,3.4866312,3.900498,4.3143644,4.7243266,5.138193,5.548156,5.2865605,5.0210614,4.755562,4.4900627,4.224563,3.8965936,3.5647192,3.2367494,2.9048753,2.5769055,2.7682211,2.9634414,3.1586614,3.3538816,3.5491016,4.1972322,4.845363,5.493494,6.141625,6.785851,6.8405128,6.89127,6.9459314,6.996689,7.0513506,6.453977,5.8566036,5.2592297,4.661856,4.0605783,3.8848803,3.7091823,3.5295796,3.3538816,3.174279,3.6232853,4.0761957,4.5252023,4.9742084,5.423215,5.1186714,4.814128,4.5095844,4.2050414,3.900498,3.8458362,3.795079,3.7443218,3.68966,3.638903,3.9317331,4.2284675,4.521298,4.8180323,5.1108627,4.860981,4.607195,4.3534083,4.1035266,3.8497405,7.629202,11.404759,15.18422,18.959778,22.739239,20.462973,18.186707,15.914344,13.638077,11.361811,9.761005,8.156297,6.5554914,4.950782,3.349977,2.7213683,2.0888553,1.4602464,0.8316377,0.19912452,0.77697605,1.3548276,1.9326792,2.5105307,3.0883822,4.1777105,5.267039,6.356367,7.445695,8.538928,8.562354,8.58578,8.6131115,8.636538,8.663869,9.741484,10.819098,11.896713,12.974329,14.048039,17.234032,20.420023,23.606016,26.788103,29.974096,31.196175,32.41825,33.644234,34.866314,36.08839,36.076675,36.068867,36.057156,36.049347,36.037632,30.356728,24.675823,18.998821,13.317916,7.6370106,6.5554914,5.477876,4.396357,3.3187418,2.2372224,3.802888,5.368553,6.9342184,8.495979,10.061645,10.760532,11.45942,12.154405,12.853292,13.548276,14.254972,14.96167,15.664462,16.371159,17.073952,18.178898,19.283842,20.388788,21.493734,22.59868,21.458595,20.31851,19.178425,18.038338,16.898252,14.27059,11.639023,9.01136,6.379793,3.7482262,3.2484627,2.7486992,2.2489357,1.7491722,1.2494087,0.999527,0.74964523,0.4997635,0.24988174,0.0,0.0,0.0,0.0,0.0,0.0,0.14055848,0.28111696,0.42167544,0.5583295,0.698888,0.94486535,1.1908426,1.43682,1.678893,1.9248703,2.3035975,2.67842,3.057147,3.435874,3.8106966,3.9746814,4.138666,4.298747,4.462732,4.6267166,4.728231,4.83365,4.939069,5.044488,5.1499066,4.4041657,3.6584249,2.9165885,2.1708477,1.4251068,1.7530766,2.0810463,2.4090161,2.7330816,3.0610514,2.6628022,2.260649,1.8623998,1.4641509,1.0619974,1.2298868,1.397776,1.5656652,1.7335546,1.901444,2.7252727,3.5491016,4.376835,5.2006636,6.0244927,6.8405128,7.656533,8.468649,9.284669,10.100689,10.268578,10.4403715,10.608261,10.780055,10.951848,10.151445,9.354948,8.55845,7.758047,6.9615493,6.9068875,6.8483214,6.7897553,6.7311897,6.676528,6.559396,6.446168,6.329036,6.2158084,6.098676,6.3719845,6.6452928,6.918601,7.191909,7.461313,8.117252,8.773191,9.4291315,10.081166,10.737106,11.838148,12.943093,14.044135,15.14908,16.250122,17.796265,19.338505,20.884647,22.430792,23.976934,24.207294,24.441559,24.671917,24.906181,25.136541,20.466877,15.797212,11.127546,6.4578815,1.7882162,5.6223392,9.456462,13.29449,17.128613,20.962736,20.93931,20.915882,20.89636,20.872934,20.849508,19.436115,18.018816,16.605423,15.188125,13.774731,22.227762,30.680794,39.133823,47.586853,56.03598,45.03728,34.038578,23.035973,12.037272,1.038571,0.8667773,0.698888,0.5270943,0.359205,0.18741131,2.3738766,4.5564375,6.7429028,8.929368,11.111929,10.229534,9.347139,8.464745,7.5823493,6.699954,11.881096,17.066143,22.247284,27.428427,32.613472,29.85306,27.092648,24.332235,21.571823,18.81141,15.828446,12.849388,9.866425,6.883461,3.900498,4.0761957,4.2557983,4.4314966,4.6110992,4.786797,6.5633,8.343708,10.120211,11.896713,13.673217,15.418485,17.163752,18.90902,20.654287,22.399555,20.459068,18.51858,16.578093,14.641508,12.70102,11.521891,10.346666,9.167537,7.988407,6.813182,6.5554914,6.297801,6.04011,5.7824197,5.5247293,5.395884,5.263134,5.134289,5.0054436,4.8765984,4.8375545,4.7985106,4.7633705,4.7243266,4.689187,4.3416953,3.9942036,3.6467118,3.2992198,2.951728,3.4007344,3.8497405,4.298747,4.7516575,5.2006636,6.153338,7.1060123,8.058686,9.01136,9.964035,10.292005,10.6238785,10.951848,11.283723,11.611692,11.6585455,11.701493,11.748346,11.791295,11.838148,12.661977,13.4858055,14.313539,15.137367,15.961197,15.324779,14.688361,14.048039,13.411622,12.775204,12.943093,13.110983,13.2788725,13.446761,13.610746,12.845484,12.076316,11.311053,10.541886,9.776623,9.440845,9.105066,8.769287,8.433509,8.101635,8.156297,8.214863,8.273428,8.32809,8.386656,8.644346,8.898132,9.151918,9.405705,9.663396,9.538455,9.4174185,9.296382,9.171441,9.050405,8.320281,7.590158,6.860035,6.1299114,5.3997884,5.095245,4.7907014,4.4861584,4.181615,3.873167,3.5608149,3.2445583,2.9283018,2.6159496,2.2996929,2.2489357,2.194274,2.1435168,2.0888553,2.0380979,2.2137961,2.3933985,2.5690966,2.7486992,2.9243972,3.193801,3.4632049,3.736513,4.0059166,4.2753205,3.7989833,3.3265507,2.8502135,2.3738766,1.901444,3.338264,4.775084,6.211904,7.648724,9.089449,9.112875,9.136301,9.163632,9.187058,9.21439,0.737932,0.7418364,0.74574083,0.75354964,0.75745404,0.76135844,0.80040246,0.8394465,0.8745861,0.9136301,0.94876975,0.94876975,0.94486535,0.94096094,0.94096094,0.93705654,0.92143893,0.9058213,0.8941081,0.8784905,0.8628729,0.9136301,0.96829176,1.0190489,1.0737107,1.1244678,1.2337911,1.33921,1.4485333,1.5539521,1.6632754,1.7101282,1.756981,1.8038338,1.8506867,1.901444,2.5612879,3.2211318,3.8809757,4.5408196,5.2006636,6.1103897,7.0201154,7.929841,8.839567,9.749292,10.768341,11.783486,12.802535,13.821584,14.836729,16.10566,17.370686,18.639616,19.908546,21.173573,19.557152,17.94073,16.324306,14.703979,13.087557,11.158782,9.2339115,7.3051367,5.376362,3.4514916,2.7604125,2.069333,1.3782539,0.6910792,0.0,0.1835069,0.3709182,0.5544251,0.7418364,0.92534333,1.2415999,1.5539521,1.8702087,2.1864653,2.4988174,2.4090161,2.3192148,2.2294137,2.1396124,2.0498111,2.1708477,2.2957885,2.416825,2.541766,2.6628022,2.4792955,2.2957885,2.1161861,1.9326792,1.7491722,1.6320401,1.5149081,1.397776,1.2806439,1.1635119,2.3543546,3.541293,4.732136,5.9229784,7.113821,8.78881,10.467703,12.146595,13.821584,15.500477,14.918721,14.336966,13.751305,13.169549,12.587793,12.376955,12.166118,11.959184,11.748346,11.537509,10.990892,10.444276,9.893755,9.347139,8.800523,8.632633,8.464745,8.296855,8.128965,7.9610763,7.8361354,7.70729,7.578445,7.453504,7.3246584,7.191909,7.0591593,6.9264097,6.79366,6.66091,6.715572,6.774138,6.8287997,6.883461,6.9381227,6.9342184,6.9342184,6.930314,6.9264097,6.9264097,6.7507114,6.578918,6.407124,6.2353306,6.0635366,6.473499,6.8873653,7.3012323,7.7111945,8.125061,8.433509,8.738052,9.0465,9.354948,9.663396,9.483793,9.304191,9.120684,8.941081,8.761478,8.031356,7.297328,6.5633,5.833177,5.099149,5.1030536,5.1030536,5.1069584,5.1108627,5.1108627,5.368553,5.6223392,5.8761253,6.133816,6.387602,6.520352,6.6531014,6.785851,6.918601,7.0513506,7.016211,6.984976,6.9537406,6.918601,6.8873653,6.461786,6.0323014,5.606722,5.1772375,4.7516575,4.4041657,4.056674,3.7091823,3.3616903,3.0141985,2.9634414,2.912684,2.8619268,2.8111696,2.7643168,2.9751544,3.1859922,3.4007344,3.611572,3.8263142,4.263607,4.7009,5.138193,5.575486,6.012779,5.9151692,5.8175592,5.7199492,5.6223392,5.5247293,4.93126,4.3338866,3.7404175,3.1430438,2.5495746,2.7682211,2.9868677,3.2016098,3.4202564,3.638903,4.1777105,4.716518,5.2592297,5.7980375,6.336845,6.336845,6.3329406,6.329036,6.329036,6.3251314,5.786324,5.2436123,4.704805,4.165997,3.6232853,3.5256753,3.4280653,3.3343596,3.2367494,3.1391394,3.6506162,4.1620927,4.6735697,5.1889505,5.700427,5.35684,5.009348,4.6657605,4.318269,3.9746814,3.9668727,3.9551594,3.9434462,3.9356375,3.9239242,4.165997,4.40807,4.6540475,4.8961205,5.138193,4.825841,4.5173936,4.2089458,3.8965936,3.5881457,7.336372,11.080693,14.828919,18.577147,22.325373,20.326319,18.32336,16.324306,14.325252,12.326198,10.588739,8.855185,7.1216297,5.3841705,3.6506162,2.9556324,2.260649,1.5656652,0.8706817,0.1756981,0.76135844,1.3431144,1.9287747,2.514435,3.1000953,4.396357,5.6965227,6.9927845,8.289046,9.589212,9.561881,9.538455,9.511124,9.487698,9.464272,9.846903,10.2334385,10.61607,11.002605,11.389141,14.95386,18.51858,22.0833,25.648018,29.212738,30.790115,32.367496,33.944874,35.52225,37.09963,35.596436,34.09324,32.59395,31.090755,29.58756,25.11702,20.646479,16.175938,11.709302,7.238762,6.1181984,4.997635,3.8770714,2.7565079,1.6359446,3.1586614,4.6813784,6.2040954,7.726812,9.249529,10.151445,11.053363,11.959184,12.861101,13.763018,14.243259,14.727406,15.211552,15.6917925,16.175938,17.456583,18.74113,20.021774,21.306324,22.586967,21.5523,20.517633,19.482967,18.448301,17.413633,14.430671,11.447707,8.464745,5.481781,2.4988174,2.3738766,2.2489357,2.1239948,1.999054,1.8741131,1.4992905,1.1244678,0.74964523,0.37482262,0.0,0.0,0.0,0.0,0.0,0.0,0.21083772,0.42167544,0.62860876,0.8394465,1.0502841,1.3157835,1.5851873,1.8506867,2.1200905,2.3855898,2.6471848,2.9087796,3.1664703,3.4280653,3.6857557,4.2011366,4.7126136,5.22409,5.735567,6.250948,6.407124,6.5633,6.7233806,6.8795567,7.0357327,6.0323014,5.02887,4.0215344,3.018103,2.0107672,2.2957885,2.5808098,2.8658314,3.1508527,3.435874,2.900971,2.3621633,1.8233559,1.2884527,0.74964523,0.96829176,1.1908426,1.4094892,1.6281357,1.8506867,2.4988174,3.1508527,3.7989833,4.4510183,5.099149,6.196286,7.2934237,8.3944645,9.491602,10.588739,10.155351,9.721962,9.288573,8.859089,8.4257,7.984503,7.5433054,7.1060123,6.6648145,6.223617,6.395411,6.5633,6.735094,6.9068875,7.0747766,6.7507114,6.4305506,6.1064854,5.786324,5.462259,5.9542136,6.4422636,6.9342184,7.422269,7.914223,8.55845,9.202676,9.846903,10.491129,11.139259,12.548749,13.958238,15.367727,16.777216,18.186707,19.65476,21.122816,22.590872,24.058928,25.523077,25.304432,25.085785,24.863234,24.644587,24.425941,19.807034,15.192029,10.573121,5.9542136,1.33921,4.7789884,8.218767,11.6585455,15.098324,18.538101,19.408783,20.28337,21.15405,22.028637,22.899319,21.216522,19.52982,17.843119,16.16032,14.473619,22.99693,31.520239,40.04355,48.56686,57.086266,45.86111,34.635952,23.410795,12.185639,0.96438736,0.8199245,0.679366,0.5349031,0.39434463,0.24988174,3.4280653,6.606249,9.784432,12.958711,16.136894,14.918721,13.704452,12.486279,11.268105,10.049932,15.906535,21.759233,27.615837,33.468536,39.325138,36.736523,34.143997,31.55538,28.96676,26.374237,22.27071,18.163279,14.059752,9.956225,5.8487945,5.8487945,5.84489,5.840986,5.840986,5.8370814,7.422269,9.007456,10.592644,12.177831,13.763018,15.516094,17.273075,19.026152,20.783133,22.53621,20.915882,19.29165,17.671324,16.047092,14.426766,13.028991,11.631214,10.2334385,8.835662,7.437886,7.309041,7.1762915,7.0474463,6.918601,6.785851,6.504734,6.223617,5.938596,5.657479,5.376362,5.349031,5.3256044,5.298274,5.2748475,5.251421,4.8961205,4.5447245,4.193328,3.8419318,3.4866312,3.8380275,4.1894236,4.5369153,4.8883114,5.2358036,6.348558,7.4574084,8.566258,9.679013,10.787864,11.096312,11.400854,11.709302,12.01775,12.326198,12.404286,12.486279,12.564366,12.6463585,12.724447,13.274967,13.825488,14.376009,14.92653,15.473146,15.274021,15.074897,14.875772,14.676648,14.473619,14.532186,14.590752,14.649317,14.703979,14.762545,14.118319,13.4740925,12.825961,12.181735,11.537509,11.23687,10.932326,10.631687,10.327144,10.0265045,10.194394,10.358379,10.526268,10.694158,10.862047,11.221252,11.576552,11.935758,12.291059,12.650263,12.095839,11.545318,10.990892,10.4403715,9.885946,8.991838,8.097731,7.2036223,6.3056097,5.4115014,5.169429,4.9234514,4.677474,4.4314966,4.1894236,3.9278288,3.6662338,3.408543,3.1469483,2.8892577,2.67842,2.4675822,2.2567444,2.0459068,1.8389735,2.1083772,2.3816853,2.6549935,2.9283018,3.2016098,3.3421683,3.4866312,3.6271896,3.7716527,3.912211,3.513962,3.1118085,2.7135596,2.3114061,1.9131571,3.338264,4.7633705,6.1884775,7.6135845,9.0386915,9.151918,9.261242,9.37447,9.487698,9.600925,0.77307165,0.77697605,0.78088045,0.78088045,0.78478485,0.78868926,0.8238289,0.8628729,0.9019169,0.93705654,0.97610056,0.96829176,0.96048295,0.95267415,0.94486535,0.93705654,0.92924774,0.92143893,0.9136301,0.9058213,0.9019169,0.93315214,0.96438736,0.9956226,1.0307622,1.0619974,1.1205635,1.183034,1.2415999,1.3040704,1.3626363,1.4407244,1.5227169,1.6008049,1.6827974,1.7608855,2.6042364,3.4475873,4.290938,5.134289,5.9737353,6.629675,7.2856145,7.941554,8.59359,9.249529,10.4286585,11.603884,12.783013,13.958238,15.137367,16.652275,18.167183,19.682093,21.197,22.711908,20.498112,18.284315,16.066616,13.852819,11.639023,10.143637,8.648251,7.152865,5.657479,4.1620927,3.330455,2.4988174,1.6632754,0.8316377,0.0,0.093705654,0.1835069,0.27721256,0.3709182,0.46071947,0.62079996,0.77697605,0.93315214,1.0932326,1.2494087,1.2064602,1.1596074,1.116659,1.0698062,1.0268579,1.1049459,1.183034,1.2650263,1.3431144,1.4251068,1.4133936,1.4055848,1.3938715,1.3860629,1.3743496,1.358732,1.3431144,1.3314011,1.3157835,1.3001659,1.9092526,2.514435,3.1235218,3.7287042,4.337791,5.0210614,5.704332,6.3836975,7.066968,7.7502384,7.90251,8.054782,8.207053,8.359325,8.511597,8.956698,9.4018,9.846903,10.292005,10.737106,10.143637,9.554072,8.960603,8.367134,7.773665,7.473026,7.168483,6.8678436,6.5633,6.262661,6.067441,5.872221,5.677001,5.481781,5.2865605,5.3021784,5.3177958,5.3334136,5.349031,5.3607445,5.602817,5.840986,6.083059,6.321227,6.5633,6.578918,6.5984397,6.6140575,6.6335793,6.649197,6.4969254,6.3407493,6.184573,6.028397,5.8761253,6.348558,6.824895,7.3012323,7.773665,8.250002,8.597494,8.944985,9.292478,9.639969,9.987461,9.874233,9.757101,9.643873,9.526741,9.413514,8.6131115,7.816613,7.0201154,6.223617,5.423215,5.3334136,5.239708,5.1460023,5.056201,4.9624953,5.1030536,5.2436123,5.3841705,5.520825,5.661383,5.985449,6.3056097,6.629675,6.9537406,7.2739015,7.37932,7.480835,7.5823493,7.6838636,7.7892823,7.2426662,6.6960497,6.153338,5.606722,5.0640097,4.607195,4.154284,3.697469,3.240654,2.787743,2.87364,2.9634414,3.049338,3.1391394,3.2250361,3.4124475,3.5998588,3.78727,3.9746814,4.1620927,4.6267166,5.087436,5.548156,6.012779,6.473499,6.5437784,6.6140575,6.6843367,6.754616,6.824895,5.9659266,5.1069584,4.2440853,3.3851168,2.5261483,2.7643168,3.0063896,3.2445583,3.4866312,3.7247996,4.1581883,4.591577,5.0210614,5.45445,5.8878384,5.8292727,5.7707067,5.716045,5.657479,5.5989127,5.1186714,4.6345253,4.154284,3.6701381,3.1859922,3.1703746,3.1508527,3.135235,3.1157131,3.1000953,3.6740425,4.251894,4.825841,5.3997884,5.9737353,5.591104,5.2045684,4.8219366,4.435401,4.0488653,4.084005,4.11524,4.1464753,4.181615,4.21285,4.4041657,4.591577,4.7828927,4.9742084,5.1616197,4.794606,4.4275923,4.0605783,3.6935644,3.3265507,7.043542,10.760532,14.477524,18.194515,21.911505,20.18576,18.463919,16.738173,15.012426,13.286681,11.420377,9.554072,7.6838636,5.8175592,3.951255,3.1898966,2.4285383,1.6710842,0.9097257,0.14836729,0.7418364,1.3353056,1.9287747,2.5183394,3.1118085,4.618908,6.1221027,7.629202,9.132397,10.6355915,10.561408,10.487225,10.413041,10.338858,10.260769,9.956225,9.647778,9.339331,9.030883,8.726339,12.6697855,16.613232,20.560583,24.504028,28.45138,30.384058,32.31674,34.249416,36.178192,38.11087,35.116196,32.121517,29.12684,26.132164,23.137487,19.877312,16.617136,13.35696,10.096785,6.8366084,5.677001,4.5173936,3.357786,2.1981785,1.038571,2.5183394,3.998108,5.477876,6.957645,8.437413,9.546264,10.651209,11.760059,12.86891,13.973856,14.235451,14.493141,14.754736,15.016331,15.274021,16.734268,18.194515,19.65476,21.115007,22.575254,21.646006,20.716759,19.783606,18.854359,17.92511,14.590752,11.256392,7.918128,4.5837684,1.2494087,1.4992905,1.7491722,1.999054,2.2489357,2.4988174,1.999054,1.4992905,0.999527,0.4997635,0.0,0.0,0.0,0.0,0.0,0.0,0.28111696,0.5583295,0.8394465,1.1205635,1.4016805,1.6906061,1.979532,2.2684577,2.5612879,2.8502135,2.9907722,3.135235,3.2757936,3.4202564,3.5608149,4.423688,5.2865605,6.1494336,7.012306,7.8751793,8.086017,8.296855,8.503788,8.714626,8.925464,7.660437,6.395411,5.1303844,3.8653584,2.6003318,2.8424048,3.084478,3.3265507,3.5686235,3.8106966,3.1391394,2.463678,1.7882162,1.1127546,0.43729305,0.7106012,0.98390937,1.2533131,1.5266213,1.7999294,2.2762666,2.7486992,3.2250361,3.7013733,4.173806,5.5559645,6.9342184,8.316377,9.694631,11.076789,10.0382185,9.0035515,7.968885,6.9342184,5.899552,5.8175592,5.735567,5.6535745,5.571582,5.4856853,5.883934,6.282183,6.6804323,7.0786815,7.47693,6.9459314,6.4149327,5.883934,5.35684,4.825841,5.532538,6.239235,6.9459314,7.656533,8.36323,8.995743,9.63216,10.268578,10.901091,11.537509,13.2554455,14.973383,16.69132,18.409256,20.12329,21.513256,22.903223,24.29319,25.683159,27.073126,26.401567,25.730011,25.058455,24.386896,23.711435,19.147188,14.582942,10.018696,5.4505453,0.8862993,3.9317331,6.9771667,10.0226,13.068034,16.113468,17.878258,19.646952,21.415646,23.184341,24.949131,22.993025,21.040823,19.084719,17.128613,15.176412,23.766096,32.359688,40.953274,49.546864,58.13655,46.684937,35.237232,23.785618,12.337912,0.8862993,0.77307165,0.6559396,0.5427119,0.42557985,0.31235218,4.482254,8.652155,12.822057,16.991959,21.16186,19.611813,18.057861,16.503908,14.95386,13.399908,19.92807,26.45623,32.98439,39.508648,46.036808,43.616077,41.199253,38.778522,36.357796,33.937065,28.70907,23.481075,18.25308,13.028991,7.800996,7.617489,7.433982,7.2543793,7.0708723,6.8873653,8.281238,9.671205,11.065076,12.458947,13.848915,15.613705,17.378494,19.143284,20.911978,22.67677,21.368793,20.064724,18.760653,17.456583,16.148607,14.532186,12.915763,11.29934,9.679013,8.062591,8.058686,8.058686,8.054782,8.050878,8.050878,7.6135845,7.180196,6.746807,6.309514,5.8761253,5.8644123,5.8487945,5.8370814,5.825368,5.813655,5.45445,5.099149,4.7399445,4.380739,4.025439,4.2753205,4.5252023,4.775084,5.024966,5.2748475,6.5437784,7.8088045,9.077735,10.346666,11.611692,11.896713,12.181735,12.466757,12.751778,13.036799,13.153932,13.2671585,13.384291,13.497519,13.610746,13.887959,14.161267,14.438479,14.711788,14.989,15.223265,15.461433,15.699601,15.93777,16.175938,16.121277,16.07052,16.015858,15.965101,15.914344,15.391153,14.867964,14.344774,13.821584,13.298394,13.028991,12.759586,12.490183,12.220779,11.951375,12.228588,12.5058,12.783013,13.0602255,13.337439,13.798158,14.258877,14.7156925,15.176412,15.637131,14.653222,13.673217,12.689307,11.709302,10.725393,9.663396,8.605303,7.5433054,6.4852123,5.423215,5.239708,5.056201,4.8687897,4.6852827,4.5017757,4.2948427,4.0918136,3.8848803,3.6818514,3.474918,3.1079042,2.7408905,2.3738766,2.0068626,1.6359446,2.0068626,2.3738766,2.7408905,3.1079042,3.474918,3.4905357,3.506153,3.521771,3.533484,3.5491016,3.2250361,2.900971,2.5769055,2.2489357,1.9248703,3.338264,4.7516575,6.1611466,7.57454,8.987934,9.187058,9.386183,9.589212,9.788337,9.987461,0.81211567,0.81211567,0.81211567,0.81211567,0.81211567,0.81211567,0.8511597,0.8862993,0.92534333,0.96438736,0.999527,0.9878138,0.97610056,0.96438736,0.94876975,0.93705654,0.93705654,0.93705654,0.93705654,0.93705654,0.93705654,0.94876975,0.96438736,0.97610056,0.9878138,0.999527,1.0112402,1.0268579,1.038571,1.0502841,1.0619974,1.175225,1.2884527,1.4016805,1.5110037,1.6242313,2.6510892,3.6740425,4.7009,5.7238536,6.7507114,7.1489606,7.551114,7.9493628,8.351517,8.749765,10.088976,11.424281,12.763491,14.098797,15.438006,17.198893,18.963682,20.724567,22.489357,24.250242,21.439074,18.623999,15.812829,13.001659,10.186585,9.124588,8.062591,7.000593,5.938596,4.8765984,3.900498,2.9243972,1.9482968,0.97610056,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.3513962,0.5114767,0.6754616,0.8394465,0.999527,1.0893283,1.175225,1.261122,1.3509232,1.43682,1.4641509,1.4875772,1.5110037,1.5383345,1.5617609,1.2494087,0.93705654,0.62470436,0.31235218,0.0,0.8862993,1.7765031,2.6628022,3.5491016,4.4393053,5.5364423,6.6374836,7.7385254,8.835662,9.936704,9.300286,8.663869,8.023546,7.387129,6.7507114,6.3134184,5.8761253,5.4388323,5.001539,4.564246,4.298747,4.037152,3.775557,3.513962,3.2484627,3.4124475,3.5764325,3.736513,3.900498,4.0605783,4.4861584,4.911738,5.337318,5.7628975,6.1884775,6.223617,6.262661,6.3017054,6.336845,6.375889,6.239235,6.098676,5.9620223,5.825368,5.688714,6.223617,6.7624245,7.3012323,7.8361354,8.374943,8.761478,9.151918,9.538455,9.924991,10.311526,10.260769,10.213917,10.163159,10.112402,10.061645,9.198771,8.335898,7.473026,6.6140575,5.7511845,5.563773,5.376362,5.1889505,5.001539,4.814128,4.8375545,4.860981,4.8883114,4.911738,4.939069,5.4505453,5.9620223,6.473499,6.98888,7.5003567,7.7385254,7.9766936,8.210958,8.449126,8.687295,8.023546,7.363703,6.699954,6.036206,5.376362,4.814128,4.251894,3.6857557,3.1235218,2.5612879,2.787743,3.0141985,3.2367494,3.4632049,3.6857557,3.8497405,4.0137253,4.173806,4.337791,4.5017757,4.985922,5.473972,5.9620223,6.4500723,6.9381227,7.1762915,7.4105554,7.648724,7.8868923,8.125061,7.000593,5.8761253,4.7516575,3.6232853,2.4988174,2.7643168,3.0259118,3.2875066,3.5491016,3.8106966,4.138666,4.462732,4.786797,5.1108627,5.4388323,5.3256044,5.212377,5.099149,4.985922,4.8765984,4.4510183,4.025439,3.5998588,3.174279,2.7486992,2.8111696,2.87364,2.9361105,2.998581,3.0610514,3.7013733,4.337791,4.9742084,5.610626,6.250948,5.825368,5.3997884,4.9742084,4.548629,4.123049,4.2011366,4.2753205,4.349504,4.423688,4.5017757,4.6384296,4.775084,4.911738,5.0483923,5.1889505,4.7633705,4.337791,3.912211,3.4866312,3.0610514,6.7507114,10.436467,14.126127,17.811884,21.501543,20.049105,18.600573,17.148134,15.699601,14.251068,12.24811,10.249056,8.250002,6.250948,4.251894,3.4241607,2.6003318,1.7765031,0.94876975,0.12494087,0.7262188,1.3235924,1.9248703,2.5261483,3.1235218,4.8375545,6.551587,8.261715,9.975748,11.685876,11.560935,11.435994,11.311053,11.186112,11.061172,10.061645,9.062118,8.062591,7.0630636,6.0635366,10.389614,14.711788,19.037865,23.363943,27.686117,29.974096,32.262077,34.550056,36.838036,39.126015,34.635952,30.149794,25.663635,21.173573,16.687416,14.637604,12.587793,10.537982,8.488171,6.4383593,5.2358036,4.037152,2.8385005,1.6359446,0.43729305,1.8741131,3.310933,4.7516575,6.1884775,7.6252975,8.937177,10.249056,11.560935,12.8767185,14.188598,14.223738,14.262781,14.301826,14.336966,14.376009,16.011953,17.651802,19.287746,20.92369,22.563541,21.735807,20.911978,20.08815,19.26432,18.436588,14.750832,11.061172,7.375416,3.6857557,0.0,0.62470436,1.2494087,1.8741131,2.4988174,3.1235218,2.4988174,1.8741131,1.2494087,0.62470436,0.0,0.0,0.0,0.0,0.0,0.0,0.3513962,0.698888,1.0502841,1.4016805,1.7491722,2.0615244,2.3738766,2.6862288,2.998581,3.310933,3.338264,3.3616903,3.3890212,3.4124475,3.435874,4.650143,5.8644123,7.0747766,8.289046,9.499411,9.761005,10.0265045,10.2881,10.549695,10.81129,9.288573,7.7619514,6.239235,4.7126136,3.1859922,3.3890212,3.5881457,3.78727,3.9863946,4.1894236,3.3734035,2.5612879,1.7491722,0.93705654,0.12494087,0.44900626,0.77307165,1.1010414,1.4251068,1.7491722,2.0498111,2.35045,2.6510892,2.951728,3.2484627,4.911738,6.575013,8.238289,9.901564,11.560935,9.924991,8.289046,6.649197,5.0132523,3.3734035,3.6506162,3.9239242,4.2011366,4.474445,4.7516575,5.376362,6.001066,6.6257706,7.250475,7.8751793,7.137247,6.3993154,5.661383,4.9234514,4.1894236,5.1108627,6.036206,6.9615493,7.8868923,8.812236,9.43694,10.061645,10.686349,11.311053,11.935758,13.962143,15.988527,18.011007,20.037392,22.063778,23.375656,24.687536,25.999414,27.311295,28.623173,27.498705,26.374237,25.24977,24.125301,23.000834,18.487345,13.973856,9.464272,4.950782,0.43729305,3.0883822,5.735567,8.386656,11.037745,13.688834,16.351637,19.010534,21.673336,24.33614,26.998941,24.773432,22.551826,20.326319,18.10081,15.875299,24.539167,33.19913,41.863003,50.52687,59.186832,47.512672,35.83851,24.16044,12.486279,0.81211567,0.7262188,0.63641757,0.5505207,0.46071947,0.37482262,5.5364423,10.698062,15.863586,21.025206,26.186827,24.300999,22.411268,20.525442,18.635712,16.749886,23.949604,31.14932,38.349037,45.548756,52.748474,50.49954,48.250603,46.001667,43.74883,41.499893,35.151333,28.79887,22.450314,16.101755,9.749292,9.386183,9.023073,8.663869,8.300759,7.9376497,9.136301,10.338858,11.537509,12.73616,13.938716,15.711315,17.487818,19.26432,21.036919,22.813423,21.82561,20.837795,19.849981,18.862167,17.874353,16.039284,14.200311,12.361338,10.526268,8.687295,8.812236,8.937177,9.062118,9.187058,9.311999,8.726339,8.136774,7.551114,6.9615493,6.375889,6.375889,6.375889,6.375889,6.375889,6.375889,6.012779,5.64967,5.2865605,4.9234514,4.564246,4.7126136,4.860981,5.0132523,5.1616197,5.3138914,6.7389984,8.164105,9.589212,11.014318,12.439425,12.70102,12.962616,13.224211,13.4858055,13.751305,13.899672,14.051944,14.200311,14.348679,14.50095,14.50095,14.50095,14.50095,14.50095,14.50095,15.176412,15.851873,16.52343,17.198893,17.874353,17.714273,17.550287,17.386303,17.226223,17.062239,16.663988,16.261835,15.863586,15.461433,15.063184,14.825015,14.586847,14.348679,14.114414,13.8762455,14.262781,14.649317,15.035853,15.426293,15.812829,16.375063,16.937298,17.49953,18.061766,18.623999,17.210606,15.801116,14.387722,12.974329,11.560935,10.338858,9.112875,7.8868923,6.66091,5.4388323,5.3138914,5.1889505,5.0640097,4.939069,4.814128,4.661856,4.513489,4.3612175,4.21285,4.0605783,3.5373883,3.0141985,2.4871042,1.9639144,1.43682,1.901444,2.3621633,2.8267872,3.2875066,3.7482262,3.638903,3.5256753,3.4124475,3.2992198,3.1859922,2.9361105,2.6862288,2.436347,2.1864653,1.9365835,3.338264,4.73604,6.13772,7.535496,8.937177,9.226103,9.511124,9.80005,10.088976,10.373997,0.78868926,0.78868926,0.79259366,0.79649806,0.79649806,0.80040246,0.8394465,0.8745861,0.9136301,0.94876975,0.9878138,0.98000497,0.97219616,0.96438736,0.95657855,0.94876975,0.95657855,0.96048295,0.96438736,0.96829176,0.97610056,0.97219616,0.96829176,0.96829176,0.96438736,0.96438736,0.9917182,1.0229534,1.0541886,1.0815194,1.1127546,1.1908426,1.2728351,1.3509232,1.4329157,1.5110037,2.3738766,3.232845,4.0918136,4.950782,5.813655,6.356367,6.902983,7.445695,7.9923115,8.538928,10.370092,12.201257,14.036326,15.867491,17.698656,18.335073,18.97149,19.604004,20.240421,20.876839,18.436588,16.00024,13.563893,11.123642,8.687295,7.7658563,6.844417,5.919074,4.997635,4.0761957,3.2640803,2.4519646,1.6359446,0.8238289,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.046852827,0.08199245,0.11713207,0.15227169,0.18741131,0.30844778,0.43338865,0.5544251,0.679366,0.80040246,0.8706817,0.94096094,1.0112402,1.0815194,1.1517987,1.1713207,1.1908426,1.2103647,1.2298868,1.2494087,1.2103647,1.1713207,1.1283722,1.0893283,1.0502841,1.9482968,2.8502135,3.7482262,4.650143,5.548156,6.3836975,7.2192397,8.054782,8.890324,9.725866,9.081639,8.441318,7.7970915,7.1567693,6.5125427,6.211904,5.911265,5.610626,5.3138914,5.0132523,5.009348,5.009348,5.0054436,5.001539,5.001539,5.134289,5.270943,5.4036927,5.5403466,5.6730967,5.8761253,6.0752497,6.2743745,6.473499,6.676528,6.66091,6.649197,6.6374836,6.6257706,6.6140575,6.4305506,6.2470436,6.0635366,5.883934,5.700427,6.2353306,6.7702336,7.3051367,7.8400397,8.374943,8.609207,8.839567,9.073831,9.304191,9.538455,9.554072,9.573594,9.589212,9.608734,9.6243515,8.913751,8.203149,7.4964523,6.785851,6.0752497,6.036206,5.9932575,5.9542136,5.9151692,5.8761253,5.891743,5.903456,5.919074,5.9346914,5.950309,6.387602,6.824895,7.262188,7.699481,8.136774,8.148487,8.164105,8.175818,8.187531,8.1992445,7.621393,7.043542,6.46569,5.891743,5.3138914,4.8883114,4.466636,4.044961,3.6232853,3.2016098,3.3070288,3.416352,3.521771,3.631094,3.736513,3.8887846,4.041056,4.193328,4.3455997,4.5017757,4.9546866,5.4115014,5.8644123,6.321227,6.774138,7.1489606,7.523783,7.898606,8.273428,8.648251,7.531592,6.4149327,5.298274,4.181615,3.0610514,3.3655949,3.6740425,3.978586,4.283129,4.5876727,4.7985106,5.009348,5.2162814,5.4271193,5.6379566,5.4388323,5.2358036,5.036679,4.8375545,4.6384296,4.396357,4.1581883,3.9161155,3.677947,3.435874,3.3929255,3.3460727,3.3031244,3.2562714,3.213323,3.7560349,4.298747,4.841459,5.3841705,5.9268827,5.6340523,5.3412223,5.0483923,4.755562,4.462732,4.5681505,4.677474,4.786797,4.892216,5.001539,4.939069,4.8805027,4.8219366,4.759466,4.7009,4.447114,4.193328,3.9434462,3.68966,3.435874,6.8483214,10.256865,13.6693125,17.077856,20.486399,19.799223,19.11205,18.424873,17.7377,17.050524,14.543899,12.033368,9.526741,7.0201154,4.513489,3.631094,2.7526035,1.8741131,0.9917182,0.113227665,0.7027924,1.2923572,1.8819219,2.4714866,3.0610514,4.415879,5.7668023,7.1216297,8.472553,9.823476,9.901564,9.979652,10.05774,10.135828,10.213917,10.081166,9.952321,9.823476,9.690726,9.561881,13.739592,17.917301,22.095013,26.272722,30.450434,31.114182,31.781834,32.445583,33.10933,33.77308,30.196648,26.620214,23.043781,19.463446,15.8870125,14.0831785,12.2793455,10.471607,8.667773,6.8639393,5.708236,4.552533,3.39683,2.241127,1.0893283,2.4519646,3.8106966,5.173333,6.5359693,7.898606,8.956698,10.0147915,11.072885,12.130978,13.189071,13.337439,13.4858055,13.638077,13.786445,13.938716,15.266212,16.59371,17.921206,19.248703,20.5762,19.842173,19.108145,18.378021,17.643993,16.91387,13.544372,10.178777,6.8092775,3.4436827,0.07418364,0.59737355,1.1205635,1.6437533,2.1669433,2.6862288,2.3465457,2.0029583,1.6593709,1.3157835,0.97610056,1.3470187,1.7218413,2.0927596,2.463678,2.8385005,2.6081407,2.3816853,2.15523,1.9287747,1.698415,2.135708,2.5769055,3.0141985,3.4514916,3.8887846,4.0527697,4.2167544,4.380739,4.548629,4.7126136,5.6535745,6.5984397,7.5394006,8.484266,9.425227,10.081166,10.741011,11.39695,12.056794,12.712734,11.584361,10.455989,9.331521,8.203149,7.0747766,7.113821,7.1489606,7.1880045,7.223144,7.262188,6.852226,6.4422636,6.0323014,5.6223392,5.212377,5.196759,5.181142,5.169429,5.153811,5.138193,5.376362,5.610626,5.8487945,6.086963,6.3251314,7.570636,8.8200445,10.069453,11.314958,12.564366,10.881569,9.202676,7.523783,5.840986,4.1620927,4.5993857,5.036679,5.473972,5.911265,6.348558,6.883461,7.4144597,7.9493628,8.480362,9.01136,8.890324,8.769287,8.644346,8.52331,8.398369,9.909373,11.420377,12.93138,14.438479,15.949483,15.726933,15.500477,15.274021,15.051471,14.825015,16.898252,18.97149,21.040823,23.114061,25.1873,26.585075,27.982851,29.380627,30.778402,32.176178,31.820879,31.469482,31.118086,30.76669,30.411388,25.53479,20.658192,15.781594,10.901091,6.0244927,8.281238,10.541886,12.798631,15.055375,17.31212,19.318983,21.321941,23.328804,25.331762,27.338625,27.338625,27.34253,27.346434,27.346434,27.350338,33.944874,40.53941,47.133945,53.72848,60.32692,48.60981,36.896603,25.179491,13.466284,1.7491722,1.8702087,1.9912452,2.1083772,2.2294137,2.35045,7.039637,11.72492,16.414106,21.09939,25.788576,23.625538,21.466404,19.30727,17.148134,14.989,23.656773,32.32064,40.988415,49.65619,58.32396,54.96227,51.60058,48.23889,44.873295,41.511604,35.04201,28.572416,22.102821,15.633226,9.163632,9.0386915,8.913751,8.78881,8.663869,8.538928,9.538455,10.537982,11.537509,12.537036,13.536563,15.832351,18.12814,20.423927,22.715813,25.0116,23.891037,22.76657,21.646006,20.521538,19.400974,17.351164,15.305257,13.25935,11.209538,9.163632,9.358852,9.554072,9.749292,9.940608,10.135828,9.386183,8.636538,7.8868923,7.137247,6.387602,6.461786,6.5359693,6.6140575,6.688241,6.7624245,6.688241,6.617962,6.5437784,6.473499,6.3993154,6.735094,7.0708723,7.406651,7.7385254,8.074304,9.468176,10.858143,12.252014,13.645885,15.035853,14.949956,14.864059,14.774258,14.688361,14.59856,14.559516,14.520472,14.481428,14.438479,14.399435,14.30573,14.215929,14.122223,14.028518,13.938716,14.6805525,15.422389,16.164225,16.906061,17.651802,17.581524,17.515148,17.448774,17.378494,17.31212,16.75379,16.191557,15.633226,15.070992,14.512663,14.243259,13.97776,13.708356,13.442857,13.173453,13.567798,13.958238,14.352583,14.743023,15.137367,15.629322,16.121277,16.613232,17.10909,17.601046,16.55076,15.504381,14.458001,13.411622,12.361338,11.424281,10.48332,9.542359,8.601398,7.6643414,7.172387,6.6843367,6.192382,5.704332,5.212377,5.0601053,4.9078336,4.755562,4.60329,4.4510183,4.0215344,3.5959544,3.1664703,2.7408905,2.3114061,2.6588979,3.0024853,3.3460727,3.6935644,4.037152,3.9395418,3.8419318,3.7443218,3.6467118,3.5491016,3.2757936,3.0063896,2.7330816,2.4597735,2.1864653,3.5686235,4.9468775,6.329036,7.70729,9.089449,9.280765,9.47208,9.663396,9.858616,10.049932,0.76135844,0.76916724,0.77307165,0.77697605,0.78088045,0.78868926,0.8238289,0.8628729,0.9019169,0.93705654,0.97610056,0.97219616,0.96829176,0.96829176,0.96438736,0.96438736,0.97219616,0.98390937,0.9917182,1.0034313,1.0112402,0.9956226,0.97610056,0.96048295,0.94096094,0.92534333,0.97219616,1.0190489,1.0659018,1.116659,1.1635119,1.2103647,1.2572175,1.3040704,1.3509232,1.4016805,2.096664,2.7916477,3.4866312,4.181615,4.8765984,5.563773,6.2548523,6.9459314,7.633106,8.324185,10.651209,12.978233,15.309161,17.636185,19.96321,19.471254,18.9793,18.48344,17.991486,17.49953,15.438006,13.376482,11.311053,9.249529,7.1880045,6.4032197,5.6223392,4.841459,4.056674,3.2757936,2.6237583,1.9756275,1.3235924,0.6754616,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.058566034,0.08980125,0.12103647,0.15617609,0.18741131,0.26940376,0.3513962,0.43338865,0.5192855,0.60127795,0.6520352,0.7066968,0.75745404,0.80821127,0.8628729,0.8784905,0.8941081,0.9058213,0.92143893,0.93705654,1.1713207,1.4016805,1.6359446,1.8663043,2.1005683,3.0141985,3.9239242,4.8375545,5.7511845,6.66091,7.230953,7.800996,8.371038,8.941081,9.511124,8.866898,8.218767,7.570636,6.9225054,6.2743745,6.114294,5.950309,5.786324,5.6262436,5.462259,5.7199492,5.9776397,6.2353306,6.493021,6.7507114,6.8561306,6.9654536,7.0708723,7.180196,7.2856145,7.262188,7.238762,7.211431,7.1880045,7.1606736,7.098203,7.0357327,6.9732623,6.910792,6.8483214,6.621866,6.395411,6.168956,5.938596,5.7121406,6.2431393,6.7780423,7.309041,7.843944,8.374943,8.453031,8.531119,8.609207,8.683391,8.761478,8.847376,8.933272,9.019169,9.101162,9.187058,8.628729,8.074304,7.5159745,6.957645,6.3993154,6.5086384,6.6140575,6.7233806,6.8287997,6.9381227,6.942027,6.9459314,6.9537406,6.957645,6.9615493,7.3246584,7.687768,8.050878,8.413987,8.773191,8.562354,8.351517,8.136774,7.9259367,7.7111945,7.2192397,6.727285,6.2353306,5.743376,5.251421,4.9663997,4.6852827,4.4041657,4.1191444,3.8380275,3.8263142,3.8185053,3.8067923,3.7989833,3.78727,3.9317331,4.0722914,4.2167544,4.357313,4.5017757,4.9234514,5.3451266,5.7668023,6.1884775,6.6140575,7.125534,7.6370106,8.148487,8.663869,9.175345,8.066495,6.9537406,5.84489,4.73604,3.6232853,3.970777,4.318269,4.6657605,5.0132523,5.3607445,5.4583545,5.55206,5.645766,5.743376,5.8370814,5.548156,5.263134,4.9742084,4.689187,4.4002614,4.3455997,4.290938,4.2362766,4.181615,4.126953,3.970777,3.8185053,3.6662338,3.513962,3.3616903,3.8106966,4.2557983,4.704805,5.153811,5.5989127,5.4388323,5.278752,5.1186714,4.958591,4.7985106,4.939069,5.0796275,5.2201858,5.3607445,5.5013027,5.2436123,4.985922,4.728231,4.4705405,4.21285,4.1308575,4.0527697,3.970777,3.892689,3.8106966,6.9459314,10.077262,13.208592,16.343828,19.475159,19.549341,19.623526,19.701614,19.775797,19.849981,16.835783,13.821584,10.803481,7.7892823,4.775084,3.8419318,2.9048753,1.9717231,1.0346665,0.10151446,0.679366,1.261122,1.8389735,2.4207294,2.998581,3.9942036,4.985922,5.9776397,6.969358,7.9610763,8.242193,8.52331,8.804427,9.081639,9.362757,10.100689,10.8425255,11.584361,12.322293,13.06413,17.093473,21.122816,25.152159,29.181503,33.210846,32.25427,31.297688,30.34111,29.380627,28.42405,25.757341,23.090635,20.423927,17.753317,15.086611,13.528754,11.966993,10.409137,8.847376,7.2856145,6.1767645,5.067914,3.959064,2.8463092,1.737459,3.0259118,4.3143644,5.5989127,6.8873653,8.175818,8.976221,9.780528,10.58093,11.385237,12.185639,12.4511385,12.712734,12.974329,13.235924,13.501423,14.516567,15.535617,16.55076,17.56981,18.58886,17.948538,17.308216,16.667892,16.02757,15.387249,12.337912,9.292478,6.2431393,3.1977055,0.14836729,0.5700427,0.9917182,1.4094892,1.8311646,2.2489357,2.1903696,2.1318035,2.069333,2.0107672,1.9482968,2.6940374,3.4397783,4.185519,4.93126,5.6730967,4.8687897,4.0644827,3.260176,2.455869,1.6515622,2.2137961,2.77603,3.338264,3.900498,4.462732,4.7672753,5.0718184,5.376362,5.6809053,5.989353,6.66091,7.3324676,8.0040245,8.675582,9.351044,10.401327,11.455516,12.5058,13.559989,14.614178,13.884054,13.153932,12.423808,11.693685,10.963562,10.838621,10.71368,10.588739,10.4637985,10.338858,10.331048,10.323239,10.315431,10.307622,10.299813,9.944512,9.589212,9.2339115,8.878611,8.52331,8.699008,8.874706,9.050405,9.226103,9.4018,10.2334385,11.065076,11.896713,12.728352,13.563893,11.838148,10.116306,8.3944645,6.6726236,4.950782,5.548156,6.1494336,6.7507114,7.348085,7.9493628,8.39056,8.831758,9.269051,9.710248,10.151445,10.6434,11.135355,11.62731,12.119265,12.611219,14.707883,16.800642,18.897306,20.99397,23.086731,22.01302,20.93931,19.861694,18.787983,17.714273,19.834364,21.95055,24.07064,26.190731,28.310822,29.794493,31.278166,32.76184,34.241608,35.72528,36.146957,36.564728,36.986404,37.404175,37.825848,32.582237,27.338625,22.098917,16.855305,11.611692,13.477997,15.344301,17.206701,19.073006,20.93931,22.286327,23.633347,24.980366,26.327385,27.674404,29.903816,32.133232,34.36655,36.595963,38.825375,43.354485,47.879684,52.40879,56.933994,61.4631,49.706944,37.954693,26.19854,14.442384,2.6862288,3.0141985,3.3421683,3.6701381,3.998108,4.3260775,8.538928,12.751778,16.960724,21.173573,25.386423,22.953981,20.521538,18.089096,15.656653,13.224211,23.360039,33.49587,43.631695,53.76362,63.89945,59.425003,54.950558,50.476112,46.001667,41.52332,34.932686,28.34596,21.75533,15.164699,8.574067,8.687295,8.800523,8.913751,9.023073,9.136301,9.936704,10.737106,11.537509,12.337912,13.138313,15.953387,18.768461,21.583536,24.39861,27.213684,25.956467,24.69925,23.438128,22.18091,20.92369,18.666946,16.410202,14.153459,11.896713,9.636065,9.901564,10.167064,10.432563,10.698062,10.963562,10.049932,9.136301,8.226576,7.3129454,6.3993154,6.551587,6.699954,6.8483214,7.000593,7.1489606,7.367607,7.5862536,7.800996,8.019642,8.238289,8.757574,9.276859,9.796145,10.319335,10.838621,12.197352,13.556085,14.918721,16.277452,17.636185,17.198893,16.761599,16.324306,15.8870125,15.449719,15.21936,14.989,14.75864,14.528281,14.301826,14.114414,13.930907,13.743496,13.559989,13.376482,14.184693,14.996809,15.80502,16.613232,17.425346,17.452679,17.48001,17.50734,17.53467,17.562002,16.843592,16.121277,15.402867,14.684457,13.962143,13.665408,13.368673,13.0719385,12.771299,12.4745655,12.872814,13.271063,13.6693125,14.063657,14.461906,14.883581,15.309161,15.730837,16.152512,16.574188,15.890917,15.211552,14.528281,13.845011,13.16174,12.5058,11.8537655,11.197825,10.541886,9.885946,9.030883,8.175818,7.320754,6.46569,5.610626,5.4583545,5.3021784,5.1460023,4.9937305,4.8375545,4.50568,4.1777105,3.8458362,3.5178664,3.1859922,3.416352,3.6428072,3.8692627,4.095718,4.3260775,4.2440853,4.1581883,4.0761957,3.9942036,3.912211,3.619381,3.3226464,3.0259118,2.7330816,2.436347,3.7989833,5.1577153,6.5164475,7.8790836,9.237816,9.335425,9.433036,9.530646,9.628256,9.725866,0.737932,0.74574083,0.75354964,0.76135844,0.76916724,0.77307165,0.81211567,0.8511597,0.8862993,0.92534333,0.96438736,0.96438736,0.96829176,0.96829176,0.97219616,0.97610056,0.9917182,1.0034313,1.0190489,1.0346665,1.0502841,1.0190489,0.98390937,0.95267415,0.92143893,0.8862993,0.95267415,1.0190489,1.0815194,1.1478943,1.2142692,1.2259823,1.2415999,1.2572175,1.2728351,1.2884527,1.815547,2.3465457,2.8775444,3.408543,3.9356375,4.7711797,5.606722,6.4422636,7.277806,8.113348,10.936231,13.759113,16.581997,19.400974,22.223858,20.60353,18.983204,17.366781,15.746454,14.126127,12.439425,10.748819,9.062118,7.375416,5.688714,5.044488,4.4041657,3.7599394,3.1157131,2.475391,1.9873407,1.4992905,1.0112402,0.5231899,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.06637484,0.09761006,0.12884527,0.15617609,0.18741131,0.23035973,0.27330816,0.31625658,0.359205,0.39824903,0.43338865,0.46852827,0.5036679,0.5388075,0.57394713,0.58566034,0.59346914,0.60518235,0.61689556,0.62470436,1.1283722,1.6359446,2.1396124,2.6432803,3.1508527,4.0761957,5.001539,5.9268827,6.8483214,7.773665,8.078208,8.386656,8.691199,8.995743,9.300286,8.648251,7.996216,7.3441806,6.688241,6.036206,6.012779,5.989353,5.9620223,5.938596,5.911265,6.4305506,6.9459314,7.465217,7.9805984,8.499884,8.581876,8.659965,8.738052,8.8200445,8.898132,8.648251,8.398369,8.148487,7.898606,7.648724,7.5394006,7.426173,7.3129454,7.1997175,7.08649,6.813182,6.5437784,6.27047,5.997162,5.7238536,6.2548523,6.785851,7.3168497,7.843944,8.374943,8.296855,8.218767,8.140678,8.066495,7.988407,8.140678,8.292951,8.445222,8.597494,8.749765,8.343708,7.941554,7.535496,7.1294384,6.7233806,6.9810715,7.2348576,7.4886436,7.746334,8.00012,7.996216,7.988407,7.984503,7.9805984,7.9766936,8.261715,8.550641,8.835662,9.124588,9.413514,8.976221,8.538928,8.101635,7.6643414,7.223144,6.817086,6.4110284,6.001066,5.5950084,5.1889505,5.044488,4.903929,4.759466,4.618908,4.474445,4.3455997,4.220659,4.0918136,3.9668727,3.8380275,3.970777,4.1035266,4.2362766,4.369026,4.5017757,4.8883114,5.278752,5.6691923,6.0596323,6.4500723,7.098203,7.7502384,8.398369,9.050405,9.698535,8.597494,7.4964523,6.3915067,5.290465,4.1894236,4.575959,4.9663997,5.35684,5.74728,6.13772,6.1181984,6.098676,6.0791545,6.055728,6.036206,5.661383,5.2865605,4.911738,4.5369153,4.1620927,4.290938,4.423688,4.552533,4.6813784,4.814128,4.552533,4.290938,4.0332475,3.7716527,3.513962,3.8653584,4.2167544,4.5681505,4.9234514,5.2748475,5.2475166,5.2201858,5.192855,5.165524,5.138193,5.309987,5.481781,5.6535745,5.8292727,6.001066,5.5442514,5.0913405,4.6345253,4.181615,3.7247996,3.8185053,3.9083066,4.0020123,4.095718,4.1894236,7.043542,9.897659,12.751778,15.605896,18.463919,19.29946,20.138906,20.97445,21.813896,22.649437,19.127666,15.605896,12.084125,8.55845,5.036679,4.0488653,3.057147,2.069333,1.077615,0.08589685,0.6559396,1.2259823,1.796025,2.366068,2.9361105,3.5686235,4.2011366,4.83365,5.466163,6.098676,6.5828223,7.0630636,7.5472097,8.031356,8.511597,10.124115,11.732729,13.341343,14.95386,16.562475,20.44345,24.328331,28.209307,32.094185,35.975163,33.394352,30.813543,28.236637,25.655827,23.075018,21.318037,19.561056,17.804073,16.043188,14.286208,12.974329,11.6585455,10.342762,9.026978,7.7111945,6.649197,5.5832953,4.5173936,3.4514916,2.3855898,3.5998588,4.814128,6.0244927,7.238762,8.449126,8.995743,9.546264,10.09288,10.639496,11.186112,11.560935,11.935758,12.31058,12.689307,13.06413,13.770826,14.477524,15.18422,15.890917,16.601519,16.050997,15.504381,14.957765,14.411149,13.860628,11.135355,8.406178,5.6809053,2.951728,0.22645533,0.5427119,0.8589685,1.1791295,1.4953861,1.8116426,2.0341935,2.2567444,2.4792955,2.7018464,2.9243972,4.041056,5.1616197,6.278279,7.394938,8.511597,7.1294384,5.74728,4.365122,2.9829633,1.6008049,2.2879796,2.9751544,3.6623292,4.349504,5.036679,5.481781,5.9268827,6.3719845,6.817086,7.262188,7.6643414,8.066495,8.468649,8.870802,9.276859,10.721489,12.170022,13.618555,15.063184,16.511717,16.179844,15.847969,15.516094,15.18422,14.848442,14.56342,14.274494,13.985569,13.700547,13.411622,13.805966,14.204215,14.59856,14.992905,15.387249,14.6922655,13.997282,13.302299,12.607315,11.912332,12.025558,12.138786,12.24811,12.361338,12.4745655,12.892336,13.310107,13.727879,14.145649,14.56342,12.798631,11.033841,9.269051,7.504261,5.735567,6.5008297,7.262188,8.023546,8.78881,9.550168,9.897659,10.2451515,10.592644,10.940135,11.287627,12.396477,13.501423,14.610273,15.719124,16.82407,19.506393,22.184814,24.863234,27.545557,30.223978,28.299107,26.374237,24.449368,22.524496,20.599627,22.76657,24.933514,27.10436,29.271303,31.438248,33.003914,34.573483,36.13915,37.708717,39.274384,40.469128,41.659973,42.850815,44.045563,45.236404,39.629684,34.02296,28.416239,22.805614,17.198893,18.67085,20.146715,21.618675,23.090635,24.562595,25.253674,25.94085,26.631927,27.323008,28.014086,32.46901,36.927837,41.386665,45.841587,50.300415,52.76019,55.21996,57.679733,60.139507,62.59928,50.80408,39.008884,27.213684,15.418485,3.6232853,4.1581883,4.6930914,5.2318993,5.7668023,6.3017054,10.0382185,13.774731,17.511244,21.251661,24.988174,22.282423,19.576674,16.870922,14.169076,11.4633255,23.06721,34.667187,46.271072,57.87105,69.47494,63.887733,58.300533,52.713333,47.126137,41.538937,34.827267,28.119505,21.407837,14.69617,7.988407,8.335898,8.687295,9.0386915,9.386183,9.737579,10.338858,10.936231,11.537509,12.138786,12.73616,16.074425,19.408783,22.743143,26.077503,29.411861,28.01799,26.628023,25.234152,23.844185,22.450314,19.98273,17.515148,15.047566,12.579984,10.112402,10.44818,10.783959,11.115833,11.4516115,11.787391,10.71368,9.636065,8.562354,7.4886436,6.4110284,6.6374836,6.8639393,7.08649,7.3129454,7.5394006,8.046973,8.550641,9.058213,9.565785,10.073358,10.780055,11.486752,12.189544,12.89624,13.599033,14.92653,16.254026,17.581524,18.90902,20.236517,19.451733,18.663042,17.874353,17.085665,16.300879,15.879204,15.461433,15.039758,14.618082,14.200311,13.923099,13.645885,13.368673,13.091461,12.814248,13.688834,14.567325,15.445815,16.324306,17.198893,17.323833,17.44487,17.565907,17.690847,17.811884,16.933393,16.050997,15.172507,14.294017,13.411622,13.083652,12.755682,12.431617,12.103647,11.775677,12.177831,12.579984,12.982138,13.384291,13.786445,14.141745,14.493141,14.844538,15.195933,15.551234,15.231073,14.914817,14.59856,14.278399,13.962143,13.591225,13.224211,12.853292,12.482374,12.111456,10.893282,9.671205,8.453031,7.230953,6.012779,5.8566036,5.6965227,5.5403466,5.3841705,5.22409,4.9937305,4.759466,4.5291066,4.2948427,4.0605783,4.173806,4.283129,4.3924527,4.5017757,4.6110992,4.5447245,4.478349,4.40807,4.3416953,4.2753205,3.959064,3.638903,3.3226464,3.0063896,2.6862288,4.029343,5.368553,6.707763,8.046973,9.386183,9.390087,9.393991,9.393991,9.397896,9.4018,0.7106012,0.7223144,0.7340276,0.7418364,0.75354964,0.76135844,0.80040246,0.8394465,0.8745861,0.9136301,0.94876975,0.95657855,0.96438736,0.97219616,0.98000497,0.9878138,1.0073358,1.0268579,1.0463798,1.0659018,1.0893283,1.038571,0.9917182,0.94486535,0.8980125,0.8511597,0.93315214,1.0151446,1.097137,1.1791295,1.261122,1.2455044,1.2259823,1.2103647,1.1908426,1.175225,1.5383345,1.9053483,2.2684577,2.6354716,2.998581,3.978586,4.958591,5.938596,6.918601,7.898606,11.217348,14.53609,17.850927,21.169668,24.48841,21.739712,18.991013,16.246218,13.497519,10.748819,9.43694,8.125061,6.813182,5.5013027,4.1894236,3.6857557,3.182088,2.67842,2.1786566,1.6749885,1.3509232,1.0268579,0.698888,0.37482262,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.078088045,0.10541886,0.13274968,0.16008049,0.18741131,0.19131571,0.19131571,0.19522011,0.19912452,0.19912452,0.21864653,0.23426414,0.25378615,0.26940376,0.28892577,0.29283017,0.29673457,0.30063897,0.30844778,0.31235218,1.0893283,1.8663043,2.6432803,3.4241607,4.2011366,5.138193,6.0752497,7.012306,7.9493628,8.886419,8.929368,8.968412,9.007456,9.0465,9.089449,8.429605,7.773665,7.113821,6.4578815,5.801942,5.911265,6.0244927,6.13772,6.250948,6.364176,7.141152,7.918128,8.695104,9.47208,10.249056,10.303718,10.354475,10.409137,10.459893,10.510651,10.0382185,9.561881,9.089449,8.6131115,8.136774,7.9766936,7.812709,7.648724,7.4886436,7.3246584,7.008402,6.688241,6.3719845,6.055728,5.735567,6.266566,6.79366,7.320754,7.8478484,8.374943,8.140678,7.910319,7.676055,7.445695,7.211431,7.433982,7.6526284,7.871275,8.093826,8.312472,8.058686,7.8088045,7.5550184,7.3012323,7.0513506,7.453504,7.8556576,8.257811,8.659965,9.062118,9.0465,9.030883,9.019169,9.0035515,8.987934,9.198771,9.413514,9.6243515,9.839094,10.049932,9.386183,8.726339,8.062591,7.3988423,6.7389984,6.4149327,6.0908675,5.7707067,5.446641,5.12648,5.1225758,5.1186714,5.1186714,5.114767,5.1108627,4.8687897,4.6228123,4.376835,4.1308575,3.8887846,4.009821,4.1308575,4.2557983,4.376835,4.5017757,4.8570766,5.2162814,5.571582,5.930787,6.2860875,7.0747766,7.8634663,8.648251,9.43694,10.22563,9.128492,8.03526,6.9381227,5.84489,4.7516575,5.181142,5.6145306,6.0479193,6.481308,6.910792,6.7780423,6.6413884,6.5086384,6.3719845,6.239235,5.774611,5.3138914,4.8492675,4.388548,3.9239242,4.240181,4.5564375,4.8687897,5.185046,5.5013027,5.134289,4.7633705,4.396357,4.029343,3.6623292,3.9200199,4.1777105,4.435401,4.6930914,4.950782,5.056201,5.1616197,5.263134,5.368553,5.473972,5.6809053,5.883934,6.0908675,6.2938967,6.5008297,5.8487945,5.196759,4.5408196,3.8887846,3.2367494,3.5022488,3.767748,4.0332475,4.298747,4.564246,7.141152,9.718058,12.294963,14.871868,17.448774,19.049578,20.650383,22.251188,23.851994,25.448895,21.41955,17.390207,13.360865,9.331521,5.298274,4.2557983,3.2094188,2.1630387,1.1205635,0.07418364,0.63641757,1.1947471,1.7530766,2.3153105,2.87364,3.1469483,3.4202564,3.6935644,3.9668727,4.2362766,4.9234514,5.606722,6.2938967,6.9771667,7.6643414,10.143637,12.622932,15.102228,17.581524,20.06082,23.79733,27.533844,31.266453,35.002968,38.73948,34.53444,30.333302,26.12826,21.927124,17.725986,16.87873,16.031475,15.18422,14.33306,13.4858055,12.415999,11.346193,10.276386,9.20658,8.136774,7.1177254,6.098676,5.0757227,4.056674,3.0376248,4.173806,5.3138914,6.4500723,7.5862536,8.726339,9.019169,9.308095,9.600925,9.893755,10.186585,10.674636,11.162686,11.650736,12.138786,12.626837,13.021181,13.419431,13.817679,14.215929,14.614178,14.157363,13.700547,13.247637,12.790822,12.337912,9.928895,7.523783,5.114767,2.7057507,0.30063897,0.5153811,0.7301232,0.94486535,1.1596074,1.3743496,1.8819219,2.3855898,2.8892577,3.39683,3.900498,5.3919797,6.8795567,8.371038,9.858616,11.350098,9.390087,7.4300776,5.4700675,3.5100577,1.5500476,2.3621633,3.174279,3.9863946,4.7985106,5.610626,6.196286,6.7819467,7.367607,7.9532676,8.538928,8.671678,8.804427,8.933272,9.066022,9.198771,11.04165,12.884527,14.727406,16.570284,18.41316,18.475632,18.542006,18.608381,18.67085,18.737226,18.28822,17.839214,17.386303,16.937298,16.48829,17.284788,18.081287,18.88169,19.678188,20.474686,19.44002,18.405352,17.370686,16.33602,15.3013525,15.348206,15.398962,15.449719,15.500477,15.551234,15.551234,15.555139,15.559043,15.559043,15.562947,13.755209,11.947471,10.139732,8.331994,6.524256,7.4495993,8.374943,9.300286,10.22563,11.150972,11.404759,11.6585455,11.916236,12.170022,12.423808,14.149553,15.871395,17.593237,19.315079,21.036919,24.300999,27.568985,30.833065,34.097145,37.361225,34.5891,31.81307,29.037039,26.26101,23.488884,25.70268,27.916475,30.134176,32.347973,34.561768,36.21333,37.868797,39.52036,41.17192,42.823483,44.7913,46.75522,48.71913,50.68695,52.650864,46.677128,40.703392,34.733562,28.759827,22.78609,23.86761,24.949131,26.026745,27.108265,28.18588,28.22102,28.252254,28.28349,28.31863,28.349865,35.034203,41.718536,48.40678,55.091114,61.77545,62.165894,62.560238,62.950676,63.345024,63.73937,51.90122,40.066975,28.232733,16.398489,4.564246,5.3060827,6.0479193,6.7897553,7.531592,8.273428,11.537509,14.801589,18.061766,21.325846,24.586021,21.610867,18.631807,15.656653,12.677594,9.698535,22.770473,35.83851,48.910446,61.97848,75.05042,68.350464,61.650513,54.950558,48.250603,41.550648,34.717945,27.889145,21.060347,14.231546,7.3988423,7.988407,8.574067,9.163632,9.749292,10.338858,10.737106,11.139259,11.537509,11.935758,12.337912,16.191557,20.049105,23.90275,27.756395,31.613945,30.08342,28.556799,27.030176,25.503555,23.976934,21.298513,18.620094,15.941674,13.263254,10.588739,10.990892,11.39695,11.803008,12.209065,12.611219,11.373524,10.135828,8.898132,7.6643414,6.426646,6.7233806,7.0240197,7.3246584,7.6252975,7.9259367,8.722435,9.518932,10.319335,11.115833,11.912332,12.802535,13.692739,14.582942,15.473146,16.36335,17.655706,18.95197,20.24823,21.540586,22.83685,21.700668,20.564487,19.4244,18.28822,17.148134,16.539047,15.929961,15.320874,14.711788,14.098797,13.731783,13.360865,12.989946,12.619028,12.24811,13.196879,14.141745,15.086611,16.031475,16.976341,17.191084,17.409729,17.628376,17.843119,18.061766,17.023193,15.980719,14.942147,13.903577,12.861101,12.5058,12.146595,11.791295,11.43209,11.076789,11.482847,11.888905,12.298867,12.704925,13.110983,13.396004,13.677121,13.958238,14.243259,14.524376,14.571229,14.618082,14.668839,14.7156925,14.762545,14.676648,14.590752,14.508759,14.422862,14.336966,12.751778,11.166591,9.581403,7.996216,6.4110284,6.250948,6.0908675,5.930787,5.7707067,5.610626,5.477876,5.3412223,5.2084727,5.0718184,4.939069,4.93126,4.9234514,4.9156423,4.9078336,4.900025,4.8492675,4.794606,4.743849,4.689187,4.6384296,4.298747,3.959064,3.619381,3.2757936,2.9361105,4.2557983,5.579391,6.899079,8.218767,9.538455,9.444749,9.351044,9.261242,9.167537,9.073831,0.6871748,0.698888,0.7106012,0.7262188,0.737932,0.74964523,0.78868926,0.8238289,0.8628729,0.9019169,0.93705654,0.94876975,0.96438736,0.97610056,0.9878138,0.999527,1.0268579,1.0502841,1.0737107,1.1010414,1.1244678,1.0619974,0.999527,0.93705654,0.8745861,0.81211567,0.9136301,1.0112402,1.1127546,1.2142692,1.3118792,1.261122,1.2142692,1.1635119,1.1127546,1.0619974,1.261122,1.4641509,1.6632754,1.8623998,2.0615244,3.1859922,4.3143644,5.4388323,6.5633,7.687768,11.498465,15.313066,19.123762,22.938364,26.74906,22.875893,18.998821,15.125654,11.248583,7.375416,6.4383593,5.5013027,4.564246,3.6232853,2.6862288,2.3231194,1.9639144,1.6008049,1.2376955,0.8745861,0.7106012,0.5505207,0.38653582,0.22645533,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0502841,2.1005683,3.1508527,4.2011366,5.251421,6.2001905,7.1489606,8.101635,9.050405,9.999174,9.776623,9.550168,9.323712,9.101162,8.874706,8.210958,7.551114,6.8873653,6.223617,5.563773,5.813655,6.0635366,6.3134184,6.5633,6.813182,7.8517528,8.886419,9.924991,10.963562,11.998228,12.025558,12.0489855,12.076316,12.099743,12.123169,11.424281,10.725393,10.0265045,9.323712,8.624825,8.413987,8.1992445,7.988407,7.773665,7.562827,7.1997175,6.8366084,6.473499,6.114294,5.7511845,6.2743745,6.801469,7.3246584,7.8517528,8.374943,7.988407,7.601871,7.211431,6.824895,6.4383593,6.7233806,7.012306,7.3012323,7.5862536,7.8751793,7.773665,7.676055,7.57454,7.47693,7.375416,7.9259367,8.476458,9.023073,9.573594,10.124115,10.100689,10.073358,10.049932,10.0265045,9.999174,10.135828,10.276386,10.413041,10.549695,10.686349,9.80005,8.913751,8.023546,7.137247,6.250948,6.012779,5.774611,5.5364423,5.298274,5.0640097,5.2006636,5.337318,5.473972,5.610626,5.7511845,5.388075,5.024966,4.661856,4.298747,3.9356375,4.0488653,4.1620927,4.2753205,4.388548,4.5017757,4.825841,5.1499066,5.473972,5.801942,6.126007,7.0513506,7.9766936,8.898132,9.823476,10.748819,9.663396,8.574067,7.4886436,6.3993154,5.3138914,5.786324,6.262661,6.7389984,7.211431,7.687768,7.437886,7.1880045,6.9381227,6.688241,6.4383593,5.8878384,5.337318,4.786797,4.2362766,3.6857557,4.1894236,4.689187,5.1889505,5.688714,6.1884775,5.7121406,5.2358036,4.7633705,4.2870336,3.8106966,3.9746814,4.138666,4.298747,4.462732,4.6267166,4.860981,5.099149,5.337318,5.575486,5.813655,6.0518236,6.2860875,6.524256,6.7624245,7.000593,6.1494336,5.298274,4.4510183,3.5998588,2.7486992,3.1859922,3.6232853,4.0605783,4.5017757,4.939069,7.238762,9.538455,11.838148,14.13784,16.437534,18.799696,21.16186,23.524023,25.886187,28.24835,23.711435,19.174519,14.637604,10.100689,5.563773,4.462732,3.3616903,2.260649,1.1635119,0.062470436,0.61299115,1.1635119,1.7140326,2.260649,2.8111696,2.7252727,2.639376,2.5495746,2.463678,2.3738766,3.2640803,4.1503797,5.036679,5.9268827,6.813182,10.163159,13.513136,16.863113,20.21309,23.563068,27.151213,30.735455,34.3236,37.911747,41.499893,35.674522,29.849155,24.023787,18.19842,12.373051,12.439425,12.501896,12.564366,12.626837,12.689307,11.861574,11.037745,10.213917,9.386183,8.562354,7.5862536,6.6140575,5.6379566,4.661856,3.6857557,4.7516575,5.813655,6.8756523,7.9376497,8.999647,9.0386915,9.073831,9.112875,9.151918,9.187058,9.788337,10.38571,10.986988,11.588266,12.185639,12.27544,12.361338,12.4511385,12.537036,12.626837,12.263727,11.900618,11.537509,11.174399,10.81129,8.726339,6.6374836,4.548629,2.463678,0.37482262,0.48805028,0.60127795,0.7106012,0.8238289,0.93705654,1.7257458,2.5105307,3.2992198,4.087909,4.8765984,6.7389984,8.601398,10.4637985,12.326198,14.188598,11.650736,9.112875,6.575013,4.037152,1.4992905,2.436347,3.3734035,4.3143644,5.251421,6.1884775,6.910792,7.6370106,8.36323,9.089449,9.811763,9.675109,9.538455,9.4018,9.261242,9.124588,11.361811,13.599033,15.836256,18.073479,20.310701,20.775324,21.236044,21.700668,22.161386,22.62601,22.01302,21.400028,20.787037,20.174046,19.561056,20.76361,21.962263,23.160913,24.36347,25.562122,24.187773,22.813423,21.439074,20.06082,18.68647,18.674755,18.663042,18.651329,18.635712,18.623999,18.214037,17.800169,17.386303,16.976341,16.562475,14.711788,12.861101,11.014318,9.163632,7.3129454,8.398369,9.487698,10.573121,11.66245,12.751778,12.911859,13.075843,13.235924,13.399908,13.563893,15.8987255,18.237463,20.5762,22.911032,25.24977,29.09951,32.94925,36.798992,40.64873,44.498474,40.875187,37.251904,33.624714,30.001427,26.374237,28.63879,30.899439,33.163994,35.42464,37.689194,39.426655,41.164112,42.901573,44.63903,46.37649,49.113476,51.850464,54.58745,57.324432,60.06142,53.724575,47.38773,41.050884,34.71404,28.373291,29.064371,29.751545,30.43872,31.125895,31.81307,31.188366,30.563662,29.938957,29.314253,28.685644,37.599392,46.513145,55.426895,64.33674,73.25049,71.5755,69.90051,68.225525,66.55054,64.87555,52.998356,41.12507,29.247877,17.37459,5.5013027,6.4500723,7.3988423,8.351517,9.300286,10.249056,13.036799,15.824542,18.612286,21.400028,24.187773,20.935406,17.686943,14.438479,11.186112,7.9376497,22.477644,37.013733,51.549824,66.085915,80.62591,72.813194,65.00049,57.18778,49.375072,41.562363,34.612526,27.66269,20.712854,13.763018,6.813182,7.6370106,8.460839,9.288573,10.112402,10.936231,11.139259,11.338385,11.537509,11.736633,11.935758,16.312593,20.685524,25.062359,29.439194,33.812122,32.14885,30.489477,28.826202,27.162926,25.499651,22.610394,5052.0,16.835783,13.950429,11.061172,11.537509,12.013845,12.486279,12.962616,13.438952,12.037272,10.6355915,9.237816,7.8361354,6.4383593,6.813182,7.1880045,7.562827,7.9376497,8.312472,9.4018,10.487225,11.576552,12.661977,13.751305,14.825015,15.8987255,16.976341,18.05005,19.123762,20.388788,21.64991,22.911032,24.17606,25.437181,23.949604,22.462027,20.97445,19.486872,17.999294,17.198893,16.398489,15.598087,14.801589,14.001186,13.536563,13.075843,12.611219,12.150499,11.685876,12.70102,13.712261,14.723501,15.738646,16.749886,17.062239,17.37459,17.686943,17.999294,18.311647,17.112995,15.914344,14.711788,13.513136,12.31058,11.924045,11.537509,11.150972,10.764437,10.373997,10.787864,11.20173,11.611692,12.025558,12.439425,12.650263,12.861101,13.075843,13.286681,13.501423,13.911386,14.325252,14.739119,15.14908,15.562947,15.762072,15.961197,16.164225,16.36335,16.562475,14.614178,12.661977,10.71368,8.761478,6.813182,6.649197,6.4891167,6.3251314,6.1611466,6.001066,5.9620223,5.9268827,5.8878384,5.8487945,5.813655,5.688714,5.563773,5.4388323,5.3138914,5.1889505,5.1499066,5.1108627,5.0757227,5.036679,5.001539,4.6384296,4.2753205,3.912211,3.5491016,3.1859922,4.4861584,5.786324,7.08649,8.386656,9.686822,9.499411,9.311999,9.124588,8.937177,8.749765,0.698888,0.7145056,0.7301232,0.74574083,0.76135844,0.77307165,0.80430686,0.8355421,0.8667773,0.8941081,0.92534333,0.93705654,0.94876975,0.96438736,0.97610056,0.9878138,1.0073358,1.0268579,1.0463798,1.0659018,1.0893283,1.0463798,1.0034313,0.96048295,0.91753453,0.8745861,0.96048295,1.0463798,1.1283722,1.2142692,1.3001659,1.2767396,1.2494087,1.2259823,1.1986516,1.175225,1.4016805,1.6242313,1.8506867,2.0732377,2.2996929,3.2679846,4.2362766,5.2006636,6.168956,7.137247,10.975275,14.813302,18.651329,22.489357,26.32348,22.555733,18.791887,15.024139,11.256392,7.4886436,6.446168,5.407597,4.369026,3.3265507,2.2879796,2.0107672,1.737459,1.4641509,1.1869383,0.9136301,0.75354964,0.59737355,0.44119745,0.28111696,0.12494087,0.113227665,0.10541886,0.093705654,0.08589685,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.07027924,0.08980125,0.10932326,0.12884527,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.1835069,0.24597734,0.30454338,0.3631094,0.42557985,1.397776,2.3699722,3.3421683,4.3143644,5.2865605,6.153338,7.016211,7.882988,8.745861,9.612638,9.483793,9.358852,9.230007,9.101162,8.976221,8.550641,8.128965,7.70729,7.2856145,6.8639393,7.4886436,8.113348,8.738052,9.362757,9.987461,10.608261,11.232965,11.8537655,12.47847,13.09927,12.954806,12.810344,12.665881,12.521418,12.373051,11.533605,10.694158,9.854712,9.0152645,8.175818,7.9064145,7.633106,7.363703,7.094299,6.824895,6.66091,6.4969254,6.329036,6.165051,6.001066,6.5125427,7.0240197,7.5394006,8.050878,8.562354,8.187531,7.812709,7.437886,7.0630636,6.688241,6.8483214,7.012306,7.1762915,7.336372,7.5003567,7.4300776,7.3597984,7.289519,7.2192397,7.1489606,7.793187,8.441318,9.085544,9.729771,10.373997,10.120211,9.866425,9.608734,9.354948,9.101162,9.20658,9.308095,9.413514,9.518932,9.6243515,8.894228,8.160201,7.426173,6.6960497,5.9620223,5.8566036,5.74728,5.6418614,5.532538,5.423215,5.563773,5.700427,5.8370814,5.9737353,6.114294,5.8214636,5.532538,5.2436123,4.950782,4.661856,4.9156423,5.173333,5.4271193,5.6809053,5.938596,5.9932575,6.0518236,6.1103897,6.168956,6.223617,7.375416,8.52331,9.675109,10.826907,11.974802,10.4286585,8.886419,7.3402762,5.794133,4.251894,4.8961205,5.5442514,6.192382,6.8405128,7.4886436,7.4886436,7.4886436,7.4886436,7.4886436,7.4886436,6.9225054,6.356367,5.794133,5.2279944,4.661856,5.024966,5.388075,5.7511845,6.114294,6.473499,6.055728,5.6340523,5.2162814,4.794606,4.376835,4.482254,4.591577,4.6969957,4.806319,4.911738,5.1108627,5.3138914,5.5130157,5.7121406,5.911265,6.2040954,6.493021,6.7819467,7.0708723,7.363703,6.6687193,5.9776397,5.2865605,4.591577,3.900498,4.482254,5.0640097,5.645766,6.2314262,6.813182,9.108971,11.408664,13.704452,16.004145,18.299932,20.435642,22.575254,24.710962,26.850574,28.986282,24.13311,19.276033,14.422862,9.565785,4.7126136,3.7794614,2.8463092,1.9131571,0.98390937,0.05075723,0.5036679,0.95657855,1.4055848,1.8584955,2.3114061,2.5690966,2.8267872,3.084478,3.3421683,3.5998588,4.939069,6.2743745,7.6135845,8.94889,10.2881,13.583415,16.87873,20.174046,23.469362,26.760773,28.646599,30.532425,32.41825,34.304077,36.186,31.161034,26.132164,21.103294,16.07833,11.0494585,11.330575,11.615597,11.896713,12.181735,12.4628525,11.6585455,10.858143,10.053836,9.253433,8.449126,7.531592,6.6140575,5.6965227,4.7789884,3.8614538,4.73604,5.610626,6.4891167,7.363703,8.238289,8.406178,8.577971,8.745861,8.917655,9.089449,9.671205,10.256865,10.8425255,11.428185,12.013845,12.212971,12.412095,12.611219,12.814248,13.013372,12.201257,11.389141,10.573121,9.761005,8.94889,7.230953,5.5169206,3.7989833,2.0810463,0.3631094,0.6442264,0.92143893,1.2025559,1.4836729,1.7608855,2.2137961,2.6628022,3.1118085,3.5608149,4.0137253,5.481781,6.9459314,8.413987,9.882042,11.350098,9.378374,7.4105554,5.4388323,3.4710135,1.4992905,2.2059872,2.9087796,3.6154766,4.318269,5.024966,5.6145306,6.2040954,6.79366,7.3832245,7.9766936,7.8947015,7.816613,7.734621,7.656533,7.57454,9.612638,11.650736,13.688834,15.726933,17.761126,18.374117,18.987108,19.6001,20.21309,20.826082,20.24823,19.670378,19.092527,18.514675,17.936825,19.186234,20.435642,21.688955,22.938364,24.187773,22.98912,21.794373,20.595722,19.39707,18.19842,17.999294,17.796265,17.593237,17.390207,17.18718,16.968533,16.745981,16.527334,16.30869,16.086138,14.481428,12.872814,11.2642,9.655587,8.050878,8.886419,9.718058,10.553599,11.389141,12.224684,12.685403,13.146122,13.606842,14.063657,14.524376,16.683512,18.84655,21.005684,23.164818,25.323954,28.849628,32.375305,35.900978,39.426655,42.948425,39.96546,36.978592,33.995632,31.008762,28.025799,29.74764,31.469482,33.191322,34.913166,36.638912,38.69653,40.758057,42.815674,44.8772,46.938725,48.98073,51.026634,53.07254,55.118446,57.164352,51.62401,46.087563,40.55112,35.010777,29.474333,30.485573,31.496813,32.50415,33.51539,34.52663,35.651096,36.77947,37.90784,39.036213,40.160683,44.84206,49.51563,54.197006,58.87448,63.54805,61.338158,59.124363,56.91057,54.700676,52.48688,45.00214,37.517403,30.032661,22.547922,15.063184,14.56342,14.063657,13.563893,13.06413,12.564366,15.641035,18.72161,21.802181,24.882755,27.96333,27.330816,26.698303,26.06579,25.433277,24.800762,34.725754,44.650745,54.575733,64.500725,74.42571,66.53101,58.640217,50.745518,42.85472,34.96392,29.579752,24.199486,18.815315,13.431144,8.050878,9.304191,10.561408,11.814721,13.0719385,14.325252,14.247164,14.169076,14.090988,14.016804,13.938716,18.194515,22.454218,26.710016,30.965815,35.225517,33.121044,31.016571,28.908194,26.803722,24.69925,22.278519,19.861694,17.440966,15.020235,12.599506,12.849388,13.09927,13.349152,13.599033,13.848915,12.747873,11.6468315,10.541886,9.440845,8.335898,8.683391,9.030883,9.378374,9.725866,10.073358,10.955752,11.838148,12.724447,13.606842,14.489237,15.152986,15.816733,16.484386,17.148134,17.811884,18.760653,19.713327,20.662096,21.610867,22.563541,21.349272,20.131098,18.916828,17.70256,16.48829,15.926057,15.367727,14.809398,14.247164,13.688834,13.411622,13.134409,12.853292,12.576079,12.298867,13.2554455,14.208119,15.164699,16.121277,17.073952,17.593237,18.116426,18.635712,19.154997,19.674282,18.506866,17.335546,16.164225,14.996809,13.825488,13.528754,13.235924,12.939189,12.6463585,12.349625,12.70102,13.056321,13.407718,13.759113,14.114414,14.364296,14.614178,14.864059,15.113941,15.363823,15.656653,15.953387,16.246218,16.542952,16.835783,16.812357,16.788929,16.761599,16.738173,16.710842,15.168603,13.622459,12.076316,10.534078,8.987934,8.55845,8.13287,7.703386,7.277806,6.8483214,7.1450562,7.4417906,7.734621,8.031356,8.324185,8.011833,7.699481,7.387129,7.0747766,6.7624245,6.3836975,6.001066,5.6223392,5.2436123,4.860981,4.50568,4.1464753,3.7911747,3.4319696,3.076669,4.3143644,5.5559645,6.79366,8.03526,9.276859,9.413514,9.550168,9.686822,9.823476,9.964035,0.7106012,0.7301232,0.74574083,0.76526284,0.78088045,0.80040246,0.8238289,0.8433509,0.8667773,0.8902037,0.9136301,0.92534333,0.93705654,0.94876975,0.96438736,0.97610056,0.9917182,1.0034313,1.0190489,1.0346665,1.0502841,1.0268579,1.0034313,0.98390937,0.96048295,0.93705654,1.0073358,1.077615,1.1478943,1.2181735,1.2884527,1.2884527,1.2884527,1.2884527,1.2884527,1.2884527,1.5383345,1.7882162,2.0380979,2.2879796,2.5378613,3.3460727,4.1581883,4.9663997,5.7785153,6.5867267,10.44818,14.313539,18.174992,22.036446,25.901804,22.239475,18.58105,14.918721,11.260296,7.601871,6.4578815,5.3138914,4.173806,3.0298162,1.8858263,1.698415,1.5110037,1.3235924,1.1361811,0.94876975,0.79649806,0.6442264,0.49195468,0.339683,0.18741131,0.1796025,0.1717937,0.1639849,0.15617609,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.05075723,0.06637484,0.08199245,0.09761006,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.3709182,0.48805028,0.60908675,0.7301232,0.8511597,1.7452679,2.639376,3.533484,4.4314966,5.3256044,6.1064854,6.883461,7.6643414,8.445222,9.226103,9.194867,9.163632,9.136301,9.105066,9.073831,8.894228,8.710721,8.527214,8.343708,8.164105,9.163632,10.163159,11.162686,12.162213,13.16174,13.368673,13.575606,13.786445,13.993378,14.200311,13.884054,13.571702,13.2554455,12.939189,12.626837,11.6468315,10.666827,9.686822,8.706817,7.726812,7.3988423,7.0708723,6.7429028,6.4149327,6.086963,6.1181984,6.153338,6.184573,6.2158084,6.250948,6.7507114,7.250475,7.7502384,8.250002,8.749765,8.386656,8.023546,7.6643414,7.3012323,6.9381227,6.9732623,7.012306,7.0513506,7.08649,7.125534,7.08649,7.043542,7.0044975,6.9654536,6.9264097,7.6643414,8.406178,9.14411,9.885946,10.6238785,10.139732,9.655587,9.171441,8.683391,8.1992445,8.273428,8.343708,8.4178915,8.488171,8.562354,7.984503,7.406651,6.8287997,6.250948,5.6730967,5.6965227,5.7199492,5.743376,5.7668023,5.786324,5.9268827,6.0635366,6.2001905,6.336845,6.473499,6.2587566,6.04011,5.8214636,5.606722,5.388075,5.786324,6.180669,6.578918,6.9771667,7.375416,7.164578,6.9537406,6.746807,6.5359693,6.3251314,7.699481,9.073831,10.44818,11.826434,13.200784,11.197825,9.194867,7.191909,5.1889505,3.1859922,4.0059166,4.825841,5.645766,6.46569,7.2856145,7.5394006,7.7892823,8.039165,8.289046,8.538928,7.957172,7.37932,6.7975645,6.2158084,5.6379566,5.8644123,6.086963,6.3134184,6.5359693,6.7624245,6.3993154,6.0323014,5.6691923,5.3021784,4.939069,4.989826,5.040583,5.095245,5.1460023,5.2006636,5.3607445,5.5247293,5.688714,5.8487945,6.012779,6.356367,6.6960497,7.039637,7.3832245,7.726812,7.191909,6.6531014,6.1181984,5.5832953,5.0483923,5.7785153,6.504734,7.230953,7.9610763,8.687295,10.983084,13.2788725,15.570756,17.866545,20.162333,22.07549,23.988647,25.901804,27.811058,29.724215,24.55088,19.381453,14.208119,9.034787,3.8614538,3.096191,2.330928,1.5656652,0.80430686,0.039044023,0.39434463,0.74574083,1.1010414,1.456342,1.8116426,2.416825,3.018103,3.619381,4.220659,4.825841,6.6140575,8.398369,10.186585,11.974802,13.763018,17.003672,20.244326,23.481075,26.72173,29.962383,30.14589,30.329397,30.508999,30.692507,30.876013,26.64364,22.415173,18.186707,13.954333,9.725866,10.22563,10.729298,11.232965,11.736633,12.236397,11.455516,10.67854,9.897659,9.116779,8.335898,7.47693,6.617962,5.758993,4.8961205,4.037152,4.7243266,5.4115014,6.098676,6.785851,7.47693,7.7775693,8.078208,8.382751,8.683391,8.987934,9.557977,10.128019,10.698062,11.268105,11.838148,12.150499,12.4628525,12.775204,13.087557,13.399908,12.138786,10.87376,9.612638,8.351517,7.08649,5.7394714,4.3924527,3.0454338,1.698415,0.3513962,0.79649806,1.2455044,1.6906061,2.1396124,2.5886188,2.7018464,2.8111696,2.9243972,3.0376248,3.1508527,4.220659,5.2943697,6.36808,7.4417906,8.511597,7.1099167,5.708236,4.3065557,2.900971,1.4992905,1.9717231,2.4441557,2.9165885,3.3890212,3.8614538,4.318269,4.7711797,5.2279944,5.6809053,6.13772,6.114294,6.0908675,6.0713453,6.0479193,6.0244927,7.8634663,9.698535,11.537509,13.376482,15.211552,15.976814,16.738173,17.49953,18.26089,19.026152,18.48344,17.94073,17.398016,16.855305,16.312593,17.612759,18.912924,20.21309,21.513256,22.813423,21.794373,20.77142,19.75237,18.733322,17.714273,17.31993,16.925583,16.535143,16.140799,15.750359,15.723028,15.695697,15.668366,15.641035,15.613705,14.247164,12.880623,11.517986,10.151445,8.78881,9.370565,9.952321,10.534078,11.115833,11.701493,12.458947,13.216402,13.973856,14.73131,15.488764,17.468296,19.451733,21.43517,23.418604,25.398136,28.599747,31.801357,34.99906,38.200672,41.398376,39.055737,36.70919,34.36655,32.020004,29.673458,30.856491,32.039524,33.222557,34.405594,35.588627,37.97031,40.351997,42.733685,45.119274,47.500957,48.851883,50.206707,51.557632,52.908554,54.263382,49.523438,44.7874,40.051357,35.311413,30.575375,31.906775,33.23818,34.573483,35.904884,37.236286,40.117733,42.999184,45.876728,48.758175,51.63572,52.080822,52.52202,52.963215,53.408318,53.849518,51.100815,48.348213,45.599514,42.850815,40.09821,37.005924,33.909733,30.813543,27.721256,24.625065,22.67677,20.724567,18.77627,16.82407,14.875772,18.249176,21.618675,24.992079,28.365482,31.738886,33.72232,35.705757,37.6931,39.676537,41.663876,46.97386,52.287754,57.601646,62.911633,68.225525,60.252735,52.279945,44.307156,36.334366,28.361578,24.546976,20.732376,16.917774,13.103174,9.288573,10.971371,12.658072,14.34087,16.02757,17.714273,17.358973,17.003672,16.64837,16.29307,15.93777,20.076437,24.219007,28.357674,32.49634,36.638912,34.089336,31.543665,28.994091,26.448421,23.898846,21.946646,19.994444,18.042242,16.090042,14.13784,14.161267,14.188598,14.212025,14.239355,14.262781,13.458474,12.654168,11.845957,11.04165,10.237343,10.557504,10.877665,11.197825,11.517986,11.838148,12.513609,13.192975,13.868437,14.547803,15.223265,15.480955,15.734741,15.988527,16.246218,16.500004,17.136421,17.776743,18.41316,19.049578,19.685997,18.745035,17.804073,16.85921,15.918248,14.973383,14.653222,14.33306,14.016804,13.696643,13.376482,13.282777,13.189071,13.09927,13.005564,12.911859,13.809871,14.707883,15.605896,16.503908,17.40192,18.12814,18.854359,19.584482,20.310701,21.036919,19.896833,18.756748,17.616663,16.476578,15.336493,15.133463,14.934339,14.73131,14.528281,14.325252,14.618082,14.9109125,15.203742,15.4965725,15.789403,16.074425,16.36335,16.64837,16.937298,17.226223,17.40192,17.581524,17.757221,17.936825,18.112522,17.86264,17.612759,17.362877,17.112995,16.863113,15.723028,14.582942,13.442857,12.302772,11.162686,10.471607,9.776623,9.085544,8.3944645,7.699481,8.32809,8.956698,9.581403,10.2100115,10.838621,10.338858,9.839094,9.339331,8.835662,8.335898,7.6135845,6.89127,6.168956,5.446641,4.7243266,4.3729305,4.0215344,3.6662338,3.3148375,2.9634414,4.142571,5.3217,6.5008297,7.6838636,8.862993,9.323712,9.788337,10.249056,10.71368,11.174399,0.7262188,0.74574083,0.76526284,0.78478485,0.80430686,0.8238289,0.8394465,0.8550641,0.8706817,0.8862993,0.9019169,0.9136301,0.92534333,0.93705654,0.94876975,0.96438736,0.97219616,0.98390937,0.9917182,1.0034313,1.0112402,1.0112402,1.0073358,1.0034313,1.0034313,0.999527,1.0541886,1.1088502,1.1635119,1.2181735,1.2767396,1.3001659,1.3235924,1.3509232,1.3743496,1.4016805,1.6749885,1.9482968,2.2255092,2.4988174,2.77603,3.4280653,4.0801005,4.732136,5.3841705,6.036206,9.924991,13.813775,17.698656,21.58744,25.476225,21.923218,18.370213,14.817206,11.2642,7.7111945,6.46569,5.22409,3.978586,2.7330816,1.4875772,1.3860629,1.2884527,1.1869383,1.0893283,0.9878138,0.8394465,0.6910792,0.5466163,0.39824903,0.24988174,0.24597734,0.23816854,0.23426414,0.23035973,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.03513962,0.046852827,0.05466163,0.06637484,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.5544251,0.7340276,0.9136301,1.0932326,1.2767396,2.0927596,2.9087796,3.7287042,4.5447245,5.3607445,6.055728,6.7507114,7.445695,8.140678,8.835662,8.905942,8.972317,9.0386915,9.108971,9.175345,9.2339115,9.288573,9.347139,9.405705,9.464272,10.838621,12.212971,13.58732,14.96167,16.33602,16.129086,15.9221525,15.7152195,15.5082855,15.3013525,14.813302,14.329156,13.845011,13.360865,12.8767185,11.756155,10.6355915,9.515028,8.3944645,7.2739015,6.89127,6.504734,6.1181984,5.735567,5.349031,5.579391,5.8097506,6.04011,6.27047,6.5008297,6.98888,7.47693,7.9610763,8.449126,8.937177,8.58578,8.238289,7.8868923,7.5394006,7.1880045,7.098203,7.012306,6.9264097,6.8366084,6.7507114,6.7389984,6.7311897,6.719476,6.7116675,6.699954,7.535496,8.371038,9.20658,10.0382185,10.87376,10.159255,9.444749,8.730244,8.015738,7.3012323,7.3402762,7.37932,7.4183645,7.461313,7.5003567,7.0786815,6.6531014,6.2314262,5.8097506,5.388075,5.5403466,5.6926184,5.84489,5.997162,6.1494336,6.2860875,6.426646,6.5633,6.699954,6.8366084,6.6921453,6.547683,6.4032197,6.2587566,6.114294,6.6531014,7.191909,7.7307167,8.273428,8.812236,8.335898,7.8556576,7.37932,6.902983,6.426646,8.023546,9.6243515,11.225157,12.825961,14.426766,11.963089,9.503315,7.043542,4.5837684,2.1239948,3.1157131,4.1113358,5.1030536,6.094772,7.08649,7.5862536,8.086017,8.58578,9.089449,9.589212,8.991838,8.398369,7.800996,7.2075267,6.6140575,6.699954,6.785851,6.8756523,6.9615493,7.0513506,6.7389984,6.4305506,6.1181984,5.8097506,5.5013027,5.4973984,5.493494,5.493494,5.4895897,5.4856853,5.610626,5.735567,5.8644123,5.989353,6.114294,6.5086384,6.902983,7.297328,7.6916723,8.086017,7.7111945,7.3324676,6.9537406,6.578918,6.2001905,7.0708723,7.9454584,8.81614,9.690726,10.561408,12.853292,15.14908,17.440966,19.73285,22.024733,23.711435,25.398136,27.088743,28.775444,30.462147,24.972557,19.482967,13.993378,8.503788,3.0141985,2.416825,1.8194515,1.2181735,0.62079996,0.023426414,0.28111696,0.5388075,0.79649806,1.0541886,1.3118792,2.260649,3.2094188,4.154284,5.1030536,6.0518236,8.289046,10.526268,12.763491,15.000713,17.237936,20.423927,23.606016,26.792007,29.978,33.163994,31.641275,30.122463,28.603651,27.080935,25.562122,22.130152,18.698183,15.266212,11.834243,8.398369,9.120684,9.846903,10.569217,11.291532,12.013845,11.256392,10.498938,9.741484,8.98403,8.226576,7.422269,6.621866,5.8175592,5.0132523,4.21285,4.7126136,5.212377,5.7121406,6.211904,6.7116675,7.1489606,7.5823493,8.015738,8.453031,8.886419,9.440845,9.999174,10.553599,11.108025,11.66245,12.08803,12.513609,12.939189,13.360865,13.786445,12.076316,10.362284,8.648251,6.9381227,5.22409,4.2479897,3.2718892,2.2918842,1.3157835,0.3357786,0.95267415,1.5656652,2.182561,2.7994564,3.4124475,3.1859922,2.9634414,2.736986,2.514435,2.2879796,2.9634414,3.6428072,4.318269,4.997635,5.6730967,4.841459,4.0059166,3.1703746,2.3348327,1.4992905,1.7413634,1.979532,2.2216048,2.4597735,2.7018464,3.018103,3.338264,3.6584249,3.978586,4.298747,4.3338866,4.369026,4.4041657,4.4393053,4.474445,6.114294,7.7502384,9.386183,11.0260315,12.661977,13.575606,14.489237,15.398962,16.312593,17.226223,16.71865,16.211079,15.7035055,15.195933,14.688361,16.039284,17.386303,18.737226,20.08815,21.439074,20.595722,19.75237,18.90902,18.06567,17.226223,16.640562,16.058807,15.477051,14.895294,14.313539,14.477524,14.641508,14.809398,14.973383,15.137367,14.016804,12.892336,11.771772,10.647305,9.526741,9.854712,10.186585,10.514555,10.84643,11.174399,12.228588,13.286681,14.34087,15.395058,16.449247,18.256985,20.06082,21.864653,23.668486,25.476225,28.349865,31.223505,34.101048,36.97469,39.848328,38.14601,36.439785,34.733562,33.031242,31.32502,31.969246,32.609566,33.253796,33.894115,34.53834,37.244095,39.94594,42.65169,45.35744,48.06319,48.723034,49.38288,50.042725,50.702568,51.36241,47.42287,43.487232,39.551594,35.612053,31.676416,33.331882,34.983444,36.638912,38.294376,39.949844,44.58437,49.21499,53.849518,58.480137,63.11076,59.319584,55.528408,51.73333,47.942154,44.15098,40.863476,37.575966,34.28846,31.000954,27.713448,29.005804,30.302067,31.598328,32.890686,34.186947,30.786211,27.389381,23.988647,20.587914,17.18718,20.853413,24.515741,28.181976,31.84821,35.51054,40.11383,44.717117,49.320408,53.9237,58.523087,59.22588,59.924767,60.623653,61.326447,62.025333,53.97055,45.919674,37.868797,29.814016,21.763138,19.514202,17.26917,15.020235,12.771299,10.526268,12.63855,14.754736,16.870922,18.983204,21.09939,20.466877,19.834364,19.20185,18.569338,17.936825,21.958359,25.983797,30.005331,34.026867,38.0484,35.06153,32.07076,29.079988,26.089216,23.098444,21.61477,20.131098,18.64352,17.159847,15.676175,15.473146,15.274021,15.074897,14.875772,14.676648,14.169076,13.661504,13.153932,12.6463585,12.138786,12.431617,12.720543,13.013372,13.306203,13.599033,14.0714655,14.543899,15.016331,15.488764,15.961197,15.808925,15.652749,15.4965725,15.344301,15.188125,15.51219,15.836256,16.164225,16.48829,16.812357,16.140799,15.473146,14.801589,14.133936,13.462379,13.384291,13.302299,13.224211,13.142218,13.06413,13.153932,13.247637,13.341343,13.431144,13.524849,14.364296,15.203742,16.043188,16.88654,17.725986,18.659138,19.596195,20.529346,21.466404,22.399555,21.290705,20.181856,19.069101,17.96025,16.8514,16.738173,16.628849,16.519526,16.410202,16.300879,16.531239,16.765503,16.995863,17.230127,17.464392,17.788456,18.112522,18.436588,18.760653,19.088623,19.147188,19.205755,19.268225,19.326792,19.389261,18.912924,18.436588,17.964155,17.487818,17.01148,16.277452,15.543426,14.809398,14.0714655,13.337439,12.380859,11.424281,10.4637985,9.507219,8.550641,9.511124,10.471607,11.428185,12.388668,13.349152,12.661977,11.974802,11.287627,10.600452,9.913278,8.847376,7.7814736,6.715572,5.6535745,4.5876727,4.240181,3.892689,3.5451972,3.1977055,2.8502135,3.970777,5.0913405,6.211904,7.328563,8.449126,9.237816,10.0265045,10.81129,11.599979,12.388668,0.737932,0.76135844,0.78088045,0.80430686,0.8277333,0.8511597,0.8589685,0.8667773,0.8706817,0.8784905,0.8862993,0.9019169,0.9136301,0.92534333,0.93705654,0.94876975,0.95657855,0.96048295,0.96438736,0.96829176,0.97610056,0.9917182,1.0112402,1.0268579,1.0463798,1.0619974,1.1010414,1.1439898,1.183034,1.2220778,1.261122,1.3118792,1.3626363,1.4133936,1.4641509,1.5110037,1.8116426,2.1122816,2.4129205,2.7135596,3.0141985,3.506153,4.0020123,4.4978714,4.9937305,5.4856853,9.4018,13.314012,17.226223,21.138433,25.050644,21.606962,18.159374,14.7156925,11.268105,7.824422,6.477403,5.1303844,3.7833657,2.436347,1.0893283,1.0737107,1.0619974,1.0502841,1.038571,1.0268579,0.8823949,0.7418364,0.59737355,0.45681506,0.31235218,0.30844778,0.30844778,0.30454338,0.30063897,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.015617609,0.023426414,0.027330816,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.7418364,0.98000497,1.2181735,1.4602464,1.698415,2.4402514,3.1781836,3.9200199,4.661856,5.3997884,6.008875,6.621866,7.230953,7.8400397,8.449126,8.6131115,8.781001,8.944985,9.108971,9.276859,9.573594,9.870329,10.167064,10.4637985,10.764437,12.513609,14.262781,16.011953,17.761126,19.514202,18.889498,18.268698,17.643993,17.023193,16.398489,15.746454,15.090515,14.434575,13.778636,13.1266,11.8654785,10.604357,9.343235,8.086017,6.824895,6.3836975,5.938596,5.4973984,5.056201,4.6110992,5.040583,5.466163,5.8956475,6.321227,6.7507114,7.223144,7.699481,8.175818,8.648251,9.124588,8.78881,8.449126,8.113348,7.773665,7.437886,7.223144,7.012306,6.801469,6.5867267,6.375889,6.395411,6.4149327,6.434455,6.453977,6.473499,7.406651,8.335898,9.265146,10.194394,11.123642,10.178777,9.2339115,8.289046,7.3441806,6.3993154,6.407124,6.4149327,6.422742,6.4305506,6.4383593,6.168956,5.903456,5.6340523,5.368553,5.099149,5.3841705,5.6652875,5.9464045,6.2314262,6.5125427,6.649197,6.785851,6.9264097,7.0630636,7.1997175,7.1294384,7.055255,6.9810715,6.910792,6.8366084,7.519879,8.203149,8.886419,9.565785,10.249056,9.503315,8.761478,8.015738,7.269997,6.524256,8.351517,10.174872,11.998228,13.825488,15.648844,12.732256,9.815667,6.899079,3.978586,1.0619974,2.2294137,3.3929255,4.5564375,5.7238536,6.8873653,7.6370106,8.386656,9.136301,9.885946,10.6355915,10.0265045,9.4174185,8.8083315,8.1992445,7.5862536,7.5394006,7.4886436,7.437886,7.387129,7.336372,7.082586,6.8287997,6.571109,6.3173227,6.0635366,6.0049706,5.9464045,5.891743,5.833177,5.774611,5.8644123,5.950309,6.036206,6.126007,6.211904,6.66091,7.1060123,7.5550184,8.0040245,8.449126,8.23048,8.011833,7.7892823,7.570636,7.348085,8.367134,9.386183,10.401327,11.420377,12.439425,14.727406,17.019289,19.30727,21.599154,23.887133,25.351284,26.811531,28.27568,29.735928,31.200079,25.394232,19.584482,13.778636,7.968885,2.1630387,1.7335546,1.3040704,0.8706817,0.44119745,0.011713207,0.1717937,0.3318742,0.49195468,0.6520352,0.81211567,2.1044729,3.39683,4.689187,5.9815445,7.2739015,9.964035,12.650263,15.336493,18.026625,20.712854,23.844185,26.971611,30.102942,33.234272,36.3617,33.140568,29.919434,26.694399,23.473267,20.24823,17.616663,14.981192,12.34572,9.710248,7.0747766,8.015738,8.960603,9.901564,10.84643,11.787391,11.053363,10.319335,9.581403,8.847376,8.113348,7.367607,6.621866,5.8761253,5.134289,4.388548,4.7009,5.0132523,5.3256044,5.6379566,5.950309,6.5164475,7.08649,7.6526284,8.218767,8.78881,9.327617,9.866425,10.409137,10.947944,11.486752,12.025558,12.564366,13.09927,13.638077,14.176885,12.013845,9.850807,7.687768,5.5247293,3.3616903,2.7565079,2.1474214,1.5383345,0.93315214,0.3240654,1.1088502,1.8897307,2.6706111,3.455396,4.2362766,3.6740425,3.1118085,2.5495746,1.9873407,1.4251068,1.7062237,1.9912452,2.2723622,2.5534792,2.8385005,2.5690966,2.3035975,2.0341935,1.7686942,1.4992905,1.5070993,1.5149081,1.5227169,1.5305257,1.5383345,1.7218413,1.9092526,2.0927596,2.2762666,2.463678,2.5534792,2.6471848,2.7408905,2.8306916,2.9243972,4.3612175,5.7980375,7.238762,8.675582,10.112402,11.174399,12.236397,13.298394,14.364296,15.426293,14.95386,14.481428,14.008995,13.536563,13.06413,14.461906,15.863586,17.261362,18.663042,20.06082,19.39707,18.733322,18.06567,17.40192,16.738173,15.965101,15.192029,14.418958,13.645885,12.8767185,13.232019,13.591225,13.946525,14.30573,14.661031,13.78254,12.90405,12.021654,11.143164,10.260769,10.338858,10.416945,10.495033,10.573121,10.651209,12.002132,13.353056,14.707883,16.058807,17.413633,19.041769,20.666,22.294136,23.922272,25.550407,28.099983,30.649557,33.19913,35.748707,38.298283,37.236286,36.170383,35.10448,34.038578,32.97658,33.078094,33.17961,33.281124,33.386543,33.48806,36.51397,39.543785,42.5697,45.595608,48.625427,48.59419,48.55905,48.527817,48.496582,48.46144,45.326206,42.187065,39.05183,35.912693,32.773552,34.753086,36.72871,38.708244,40.683872,42.663403,49.0471,55.430798,61.8184,68.202095,74.58579,66.55834,58.530895,50.503445,42.47599,34.44854,30.626131,26.799816,22.973503,19.151093,15.324779,21.009588,26.694399,32.379208,38.06402,43.74883,38.89956,34.050293,29.201025,24.351757,19.498585,23.45765,27.416712,31.371872,35.330936,39.286095,46.50924,53.72848,60.94772,68.16696,75.3862,71.47399,67.561775,63.649567,59.737354,55.82514,47.692272,39.559402,31.426535,23.293663,15.160794,14.481428,13.802062,13.122696,12.44333,11.763964,14.30573,16.8514,19.39707,21.942741,24.48841,23.578686,22.668959,21.759233,20.845604,19.935879,23.844185,27.748587,31.652988,35.557392,39.461792,36.029823,32.597855,29.165884,25.733915,22.29804,21.282896,20.263847,19.248703,18.229654,17.210606,16.788929,16.36335,15.93777,15.51219,15.086611,14.875772,14.668839,14.458001,14.247164,14.036326,14.301826,14.567325,14.832824,15.098324,15.363823,15.629322,15.8987255,16.164225,16.43363,16.69913,16.136894,15.570756,15.004618,14.438479,13.8762455,13.887959,13.899672,13.911386,13.923099,13.938716,13.540467,13.142218,12.743969,12.34572,11.951375,12.111456,12.271536,12.431617,12.591698,12.751778,13.028991,13.306203,13.583415,13.860628,14.13784,14.918721,15.7035055,16.484386,17.26917,18.05005,19.194042,20.334127,21.478117,22.618202,23.762192,22.680674,21.603058,20.521538,19.443924,18.362404,18.346786,18.327265,18.311647,18.292124,18.276506,18.448301,18.620094,18.791887,18.963682,19.13938,19.498585,19.861694,20.224804,20.587914,20.951023,20.892456,20.83389,20.779228,20.720663,20.662096,19.96321,19.26432,18.56153,17.86264,17.163752,16.831879,16.503908,16.172033,15.844065,15.51219,14.2901125,13.068034,11.845957,10.6238785,9.4018,10.694158,11.986515,13.2788725,14.571229,15.863586,14.989,14.11051,13.235924,12.361338,11.486752,10.081166,8.671678,7.266093,5.8566036,4.4510183,4.1074314,3.7638438,3.4241607,3.0805733,2.736986,3.7989833,4.8570766,5.919074,6.9771667,8.039165,9.151918,10.260769,11.373524,12.486279,13.599033,0.74964523,0.77307165,0.80040246,0.8238289,0.8511597,0.8745861,0.8745861,0.8745861,0.8745861,0.8745861,0.8745861,0.8862993,0.9019169,0.9136301,0.92534333,0.93705654,0.93705654,0.93705654,0.93705654,0.93705654,0.93705654,0.97610056,1.0112402,1.0502841,1.0893283,1.1244678,1.1517987,1.175225,1.1986516,1.2259823,1.2494087,1.3235924,1.4016805,1.475864,1.5500476,1.6242313,1.9482968,2.2762666,2.6003318,2.9243972,3.2484627,3.5881457,3.9239242,4.263607,4.5993857,4.939069,8.874706,12.814248,16.749886,20.689428,24.625065,21.2868,17.948538,14.614178,11.275913,7.9376497,6.4891167,5.036679,3.5881457,2.135708,0.6871748,0.76135844,0.8394465,0.9136301,0.9878138,1.0619974,0.92534333,0.78868926,0.6481308,0.5114767,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,0.92534333,1.2259823,1.5266213,1.8233559,2.1239948,2.787743,3.4514916,4.1113358,4.775084,5.4388323,5.9620223,6.4891167,7.012306,7.5394006,8.062591,8.324185,8.58578,8.85128,9.112875,9.37447,9.913278,10.44818,10.986988,11.525795,12.0606985,14.188598,16.312593,18.436588,20.560583,22.688482,21.64991,20.61134,19.576674,18.538101,17.49953,16.675701,15.851873,15.024139,14.200311,13.376482,11.974802,10.573121,9.175345,7.773665,6.375889,5.8761253,5.376362,4.8765984,4.376835,3.873167,4.5017757,5.12648,5.7511845,6.375889,7.000593,7.461313,7.9259367,8.386656,8.85128,9.311999,8.987934,8.663869,8.335898,8.011833,7.687768,7.348085,7.012306,6.676528,6.336845,6.001066,6.0518236,6.098676,6.1494336,6.2001905,6.250948,7.2739015,8.300759,9.323712,10.350571,11.373524,10.198298,9.026978,7.8517528,6.676528,5.5013027,5.473972,5.4505453,5.423215,5.3997884,5.376362,5.263134,5.1499066,5.036679,4.9234514,4.814128,5.22409,5.6379566,6.0518236,6.461786,6.8756523,7.012306,7.1489606,7.2856145,7.426173,7.562827,7.562827,7.562827,7.562827,7.562827,7.562827,8.386656,9.21439,10.0382185,10.862047,11.685876,10.674636,9.663396,8.648251,7.6370106,6.6257706,8.675582,10.725393,12.775204,14.825015,16.874826,13.501423,10.124115,6.7507114,3.3734035,0.0,1.33921,2.6745155,4.0137253,5.349031,6.688241,7.687768,8.687295,9.686822,10.686349,11.685876,11.061172,10.436467,9.811763,9.187058,8.562354,8.374943,8.187531,8.00012,7.812709,7.6252975,7.426173,7.223144,7.0240197,6.824895,6.6257706,6.5125427,6.3993154,6.2860875,6.1767645,6.0635366,6.114294,6.1611466,6.211904,6.262661,6.3134184,6.813182,7.3129454,7.812709,8.312472,8.812236,8.749765,8.687295,8.624825,8.562354,8.499884,9.663396,10.826907,11.986515,13.150026,14.313539,16.601519,18.885593,21.173573,23.461554,25.749533,26.987228,28.224924,29.46262,30.700315,31.938011,25.812004,19.685997,13.563893,7.437886,1.3118792,1.0502841,0.78868926,0.5231899,0.26159495,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,1.9482968,3.5881457,5.22409,6.8639393,8.499884,11.639023,14.774258,17.913397,21.048632,24.187773,27.260536,30.337206,33.413876,36.48664,39.56331,34.635952,29.712502,24.78905,19.861694,14.938243,13.09927,11.2642,9.425227,7.5862536,5.7511845,6.910792,8.074304,9.237816,10.401327,11.560935,10.850334,10.135828,9.425227,8.710721,8.00012,7.3129454,6.6257706,5.938596,5.251421,4.564246,4.689187,4.814128,4.939069,5.0640097,5.1889505,5.8878384,6.5867267,7.2856145,7.988407,8.687295,9.21439,9.737579,10.260769,10.787864,11.311053,11.963089,12.611219,13.263254,13.911386,14.56342,11.951375,9.339331,6.7233806,4.1113358,1.4992905,1.261122,1.0268579,0.78868926,0.5505207,0.31235218,1.261122,2.2137961,3.1625657,4.1113358,5.0640097,4.1620927,3.2640803,2.3621633,1.4641509,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.30063897,0.60127795,0.9019169,1.1986516,1.4992905,1.2767396,1.0502841,0.8238289,0.60127795,0.37482262,0.42557985,0.47633708,0.5231899,0.57394713,0.62470436,0.77307165,0.92534333,1.0737107,1.2259823,1.3743496,2.612045,3.8497405,5.087436,6.3251314,7.562827,8.773191,9.987461,11.20173,12.412095,13.626364,13.189071,12.751778,12.31058,11.873287,11.435994,12.888432,14.336966,15.789403,17.237936,18.68647,18.19842,17.714273,17.226223,16.738173,16.250122,15.285735,14.325252,13.360865,12.400381,11.435994,11.986515,12.537036,13.087557,13.638077,14.188598,13.548276,12.911859,12.27544,11.639023,10.998701,10.826907,10.651209,10.475512,10.299813,10.124115,11.775677,13.423335,15.074897,16.72646,18.374117,19.826555,21.275087,22.723621,24.17606,25.624592,27.850101,30.075611,32.30112,34.52663,36.748234,36.326557,35.900978,35.4754,35.04982,34.62424,34.186947,33.749653,33.31236,32.87507,32.437775,35.78775,39.13773,42.487705,45.83768,49.18766,48.46144,47.73913,47.01291,46.28669,45.564373,43.225636,40.8869,38.548164,36.21333,33.874596,36.174286,38.47398,40.773674,43.073364,45.37306,53.513737,61.650513,69.787285,77.92406,86.06084,73.80101,61.537285,49.273556,37.013733,24.750006,20.388788,16.023666,11.66245,7.3012323,2.9361105,13.013372,23.086731,33.163994,43.23735,53.310707,47.01291,40.7112,34.413403,28.111696,21.813896,26.061886,30.31378,34.561768,38.813663,43.061653,52.900745,62.735935,72.57503,82.41412,92.24931,83.726006,75.198784,66.675476,58.148262,49.624954,41.41009,33.19913,24.988174,16.773312,8.562354,9.448653,10.338858,11.225157,12.111456,13.001659,15.976814,18.948065,21.923218,24.898373,27.873528,26.68659,25.499651,24.312714,23.125774,21.938837,25.726107,29.513376,33.300648,37.087917,40.875187,36.998116,33.12495,29.251781,25.37471,21.501543,20.951023,20.400501,19.849981,19.29946,18.74894,18.10081,17.448774,16.800642,16.148607,15.500477,15.586374,15.676175,15.762072,15.851873,15.93777,16.175938,16.414106,16.64837,16.88654,17.124708,17.18718,17.24965,17.31212,17.37459,17.437061,16.46096,15.488764,14.512663,13.536563,12.564366,12.263727,11.963089,11.66245,11.361811,11.061172,10.936231,10.81129,10.686349,10.561408,10.436467,10.838621,11.23687,11.639023,12.037272,12.439425,12.900145,13.360865,13.825488,14.286208,14.750832,15.473146,16.199366,16.925583,17.651802,18.374117,5052.0,21.075964,22.426888,23.773905,25.124828,24.074545,23.02426,21.973976,20.92369,19.873407,19.951496,20.025679,20.099863,20.174046,20.24823,20.361458,20.474686,20.587914,20.701141,20.81437,21.212618,21.610867,22.01302,22.411268,22.813423,22.637724,22.462027,22.286327,22.11063,21.938837,21.013493,20.08815,19.162806,18.237463,17.31212,17.386303,17.464392,17.538574,17.612759,17.686943,16.199366,14.711788,13.224211,11.736633,10.249056,11.873287,13.501423,15.125654,16.749886,18.374117,17.31212,16.250122,15.188125,14.126127,13.06413,11.311053,9.561881,7.812709,6.0635366,4.3143644,3.9746814,3.638903,3.2992198,2.9634414,2.6237583,3.6232853,4.6267166,5.6262436,6.6257706,7.6252975,9.062118,10.498938,11.935758,13.376482,14.813302,0.78868926,0.81211567,0.8394465,0.8628729,0.8862993,0.9136301,0.9136301,0.9136301,0.9136301,0.9136301,0.9136301,0.92534333,0.93705654,0.94876975,0.96438736,0.97610056,0.9878138,0.999527,1.0112402,1.0268579,1.038571,1.0619974,1.0893283,1.1127546,1.1361811,1.1635119,1.1869383,1.2142692,1.2376955,1.261122,1.2884527,1.3470187,1.4055848,1.4680552,1.5266213,1.5890918,1.8389735,2.0927596,2.3465457,2.5964274,2.8502135,3.4593005,4.0644827,4.6735697,5.278752,5.8878384,9.4174185,12.946998,16.476578,20.006157,23.535736,20.24823,16.95682,13.6693125,10.377901,7.08649,5.813655,4.5408196,3.2718892,1.999054,0.7262188,0.77307165,0.8238289,0.8745861,0.92534333,0.97610056,0.8472553,0.71841,0.59346914,0.46462387,0.3357786,0.3357786,0.3318742,0.3318742,0.3279698,0.3240654,0.26159495,0.19522011,0.12884527,0.06637484,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.20693332,0.30844778,0.40996224,0.5114767,0.8823949,1.2533131,1.6242313,1.9912452,2.3621633,2.9946766,3.6271896,4.2597027,4.892216,5.5247293,6.0635366,6.5984397,7.137247,7.676055,8.210958,8.581876,8.952794,9.323712,9.690726,10.061645,10.346666,10.627783,10.9089,11.193921,11.475039,13.431144,15.391153,17.34726,19.303364,21.263374,20.28337,19.303364,18.32336,17.343355,16.36335,15.457528,14.551707,13.645885,12.743969,11.838148,10.674636,9.511124,8.351517,7.1880045,6.0244927,5.7707067,5.520825,5.267039,5.0132523,4.7633705,5.3295093,5.8956475,6.46569,7.0318284,7.601871,7.793187,7.984503,8.175818,8.371038,8.562354,8.273428,7.988407,7.699481,7.4105554,7.125534,6.9732623,6.824895,6.676528,6.524256,6.375889,6.321227,6.27047,6.2158084,6.165051,6.114294,6.8287997,7.5433054,8.257811,8.972317,9.686822,8.769287,7.8517528,6.9342184,6.016684,5.099149,5.0796275,5.0601053,5.040583,5.0210614,5.001539,4.9663997,4.9351645,4.903929,4.8687897,4.8375545,5.2592297,5.6809053,6.1064854,6.5281606,6.949836,7.137247,7.3246584,7.5120697,7.699481,7.8868923,7.8556576,7.824422,7.7892823,7.758047,7.726812,8.374943,9.023073,9.675109,10.323239,10.975275,10.112402,9.249529,8.386656,7.523783,6.66091,8.468649,10.276386,12.084125,13.891863,15.699601,12.661977,9.6243515,6.5867267,3.5491016,0.5114767,1.8311646,3.1508527,4.474445,5.794133,7.113821,8.113348,9.112875,10.112402,11.111929,12.111456,11.818625,11.521891,11.229061,10.932326,10.6355915,10.213917,9.788337,9.362757,8.937177,8.511597,8.234385,7.957172,7.6799593,7.4027467,7.125534,7.0708723,7.0201154,6.969358,6.914696,6.8639393,6.832704,6.801469,6.774138,6.7429028,6.7116675,7.211431,7.70729,8.203149,8.702912,9.198771,9.167537,9.136301,9.101162,9.069926,9.0386915,10.272482,11.506273,12.743969,13.97776,15.211552,17.698656,20.181856,22.668959,25.152159,27.639263,27.935999,28.232733,28.529467,28.826202,29.12684,23.574781,18.026625,12.4745655,6.9264097,1.3743496,1.1010414,0.8238289,0.5505207,0.27330816,0.0,0.12884527,0.26159495,0.39044023,0.5192855,0.6481308,2.366068,4.084005,5.801942,7.519879,9.237816,12.0489855,14.856251,17.66742,20.47859,23.285854,25.67535,28.06094,30.450434,32.83602,35.225517,30.708124,26.194635,21.681147,17.163752,12.650263,11.549222,10.44818,9.351044,8.250002,7.1489606,7.9337454,8.714626,9.499411,10.280292,11.061172,10.61607,10.170968,9.725866,9.280765,8.835662,8.121157,7.406651,6.6921453,5.9776397,5.263134,5.3021784,5.3412223,5.3841705,5.423215,5.462259,6.0908675,6.715572,7.3441806,7.9727893,8.601398,9.14411,9.690726,10.2334385,10.780055,11.326671,11.736633,12.146595,12.556558,12.96652,13.376482,11.240774,9.108971,6.9771667,4.845363,2.7135596,2.6276627,2.541766,2.455869,2.3738766,2.2879796,2.6588979,3.0259118,3.39683,3.767748,4.138666,3.416352,2.6940374,1.9717231,1.2494087,0.5231899,0.42167544,0.31625658,0.21083772,0.10541886,0.0,0.23816854,0.48024148,0.71841,0.96048295,1.1986516,1.0190489,0.8394465,0.659844,0.48024148,0.30063897,0.3474918,0.39434463,0.44119745,0.48805028,0.5388075,0.7340276,0.92924774,1.1205635,1.3157835,1.5110037,2.5261483,3.541293,4.5564375,5.571582,6.5867267,7.605776,8.62092,9.639969,10.6590185,11.674163,11.256392,10.834716,10.413041,9.99527,9.573594,10.768341,11.963089,13.16174,14.356487,15.551234,15.125654,14.703979,14.282304,13.860628,13.438952,12.919667,12.404286,11.885,11.365715,10.850334,11.205634,11.564839,11.924045,12.2793455,12.63855,12.029464,11.424281,10.815194,10.206107,9.600925,9.593117,9.589212,9.585307,9.581403,9.573594,11.123642,12.6697855,14.215929,15.765976,17.31212,18.678661,20.049105,21.415646,22.782187,24.148727,25.86276,27.576794,29.28692,31.000954,32.711082,32.543194,32.3714,32.20351,32.031715,31.863827,31.606136,31.35235,31.098564,30.840874,30.587088,33.105427,35.623768,38.138203,40.65654,43.17488,42.905476,42.636074,42.36667,42.09336,41.823956,40.785385,39.746815,38.704338,37.665768,36.623295,38.716053,40.80881,42.901573,44.99433,47.08709,53.248238,59.40548,65.56663,71.727776,77.88892,66.89022,55.891518,44.89282,33.89802,22.899319,19.23699,15.57466,11.912332,8.250002,4.5876727,13.884054,23.176533,32.47291,41.769295,51.06177,46.20079,41.335907,36.474926,31.613945,26.74906,31.293783,35.834602,40.37933,44.920147,49.460968,55.93837,62.41187,68.889275,75.36277,81.83627,74.06261,66.29285,58.51918,50.745518,42.975754,37.423695,31.871635,26.315672,20.76361,15.211552,16.500004,17.788456,19.07691,20.361458,21.64991,22.965694,24.281477,25.593357,26.90914,28.224924,27.287867,26.350811,25.413754,24.476698,23.535736,26.573362,29.607082,32.640804,35.67843,38.712147,35.409023,32.1059,28.80668,25.503555,22.200432,22.258997,22.321468,22.380033,22.4386,22.50107,21.360985,20.2209,19.080814,17.94073,16.800642,16.976341,17.155943,17.331642,17.511244,17.686943,18.011007,18.33117,18.655233,18.9793,19.29946,18.799696,18.299932,17.800169,17.300406,16.800642,16.113468,15.430198,14.746927,14.059752,13.376482,13.286681,13.200784,13.110983,13.025085,12.939189,12.755682,12.572175,12.388668,12.209065,12.025558,12.0489855,12.076316,12.099743,12.123169,12.150499,12.572175,12.993851,13.419431,13.841106,14.262781,14.770353,15.277926,15.785499,16.29307,16.800642,17.847023,18.893402,19.943687,20.990067,22.036446,21.501543,20.96664,20.431738,19.896833,19.36193,19.646952,19.931974,20.216995,20.502016,20.787037,20.80656,20.822178,20.8417,20.857317,20.876839,21.142338,21.411741,21.677242,21.946646,22.212145,22.20824,22.204336,22.196527,22.192623,22.188719,21.353176,20.521538,19.689901,18.858263,18.026625,17.99539,17.964155,17.936825,17.905588,17.874353,16.574188,15.270117,13.966047,12.665881,11.361811,12.70102,14.044135,15.383345,16.722555,18.061766,17.054428,16.047092,15.039758,14.032422,13.025085,11.6351185,10.2451515,8.855185,7.465217,6.0752497,5.520825,4.9663997,4.40807,3.853645,3.2992198,4.2479897,5.196759,6.141625,7.0903945,8.039165,9.308095,10.577025,11.845957,13.118792,14.387722,0.8238289,0.8511597,0.8745861,0.9019169,0.92534333,0.94876975,0.94876975,0.94876975,0.94876975,0.94876975,0.94876975,0.96438736,0.97610056,0.9878138,0.999527,1.0112402,1.038571,1.0619974,1.0893283,1.1127546,1.1361811,1.1517987,1.1635119,1.175225,1.1869383,1.1986516,1.2259823,1.2494087,1.2767396,1.3001659,1.3235924,1.3704453,1.4133936,1.4602464,1.5031948,1.5500476,1.7296503,1.9092526,2.0888553,2.2684577,2.4480603,3.3265507,4.2050414,5.083532,5.958118,6.8366084,9.96013,13.083652,16.20327,19.326792,22.450314,19.205755,15.965101,12.720543,9.479889,6.239235,5.142098,4.0488653,2.951728,1.8584955,0.76135844,0.78868926,0.81211567,0.8394465,0.8628729,0.8862993,0.76916724,0.6520352,0.5349031,0.41777104,0.30063897,0.29673457,0.28892577,0.28502136,0.28111696,0.27330816,0.21864653,0.1639849,0.10932326,0.05466163,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,0.8394465,1.2806439,1.7218413,2.1591344,2.6003318,3.2016098,3.8067923,4.40807,5.009348,5.610626,6.1611466,6.7116675,7.262188,7.812709,8.36323,8.839567,9.315904,9.796145,10.272482,10.748819,10.77615,10.803481,10.8308115,10.858143,10.889378,12.677594,14.465811,16.25793,18.046146,19.838268,18.916828,17.991486,17.070047,16.148607,15.223265,14.239355,13.2554455,12.271536,11.283723,10.299813,9.37447,8.449126,7.523783,6.5984397,5.6730967,5.6691923,5.6652875,5.661383,5.6535745,5.64967,6.1611466,6.6687193,7.180196,7.6916723,8.1992445,8.121157,8.043069,7.968885,7.890797,7.812709,7.562827,7.3129454,7.0630636,6.813182,6.5633,6.5984397,6.6374836,6.676528,6.7116675,6.7507114,6.5945354,6.4383593,6.2860875,6.1299114,5.9737353,6.379793,6.785851,7.191909,7.5940623,8.00012,7.3402762,6.6804323,6.0205884,5.3607445,4.7009,4.6852827,4.6696653,4.6540475,4.6384296,4.6267166,4.6735697,4.7204223,4.7672753,4.814128,4.860981,5.2943697,5.727758,6.1611466,6.590631,7.0240197,7.262188,7.5003567,7.7385254,7.9766936,8.210958,8.148487,8.082112,8.015738,7.9532676,7.8868923,8.36323,8.835662,9.311999,9.788337,10.260769,9.550168,8.835662,8.125061,7.4105554,6.699954,8.265619,9.8312845,11.39695,12.958711,14.524376,11.826434,9.124588,6.426646,3.7247996,1.0268579,2.3270237,3.631094,4.93126,6.2353306,7.5394006,8.538928,9.538455,10.537982,11.537509,12.537036,12.572175,12.607315,12.642454,12.677594,12.712734,12.0489855,11.389141,10.725393,10.061645,9.4018,9.0465,8.691199,8.335898,7.9805984,7.6252975,7.633106,7.6409154,7.648724,7.656533,7.6643414,7.551114,7.4417906,7.3324676,7.223144,7.113821,7.605776,8.101635,8.597494,9.093353,9.589212,9.585307,9.581403,9.581403,9.577498,9.573594,10.881569,12.189544,13.497519,14.805493,16.113468,18.795792,21.478117,24.16044,26.842766,29.52509,28.880863,28.240541,27.596315,26.955994,26.311768,21.337559,16.36335,11.389141,6.4110284,1.43682,1.1517987,0.8628729,0.57394713,0.28892577,0.0,0.19912452,0.39434463,0.59346914,0.78868926,0.9878138,2.7838387,4.5837684,6.379793,8.175818,9.975748,12.458947,14.938243,17.421442,19.904642,22.387842,24.086258,25.788576,27.486992,29.189312,30.887726,26.780294,22.67677,18.573242,14.465811,10.362284,9.999174,9.636065,9.276859,8.913751,8.550641,8.952794,9.354948,9.757101,10.159255,10.561408,10.38571,10.206107,10.03041,9.850807,9.675109,8.933272,8.191436,7.445695,6.703859,5.9620223,5.919074,5.872221,5.8292727,5.7824197,5.735567,6.2938967,6.8483214,7.4027467,7.957172,8.511597,9.077735,9.643873,10.206107,10.772245,11.338385,11.506273,11.678067,11.845957,12.01775,12.185639,10.534078,8.882515,7.230953,5.579391,3.9239242,3.9942036,4.0605783,4.126953,4.193328,4.263607,4.0527697,3.8419318,3.631094,3.4241607,3.213323,2.6667068,2.1239948,1.5773785,1.0307622,0.48805028,0.39044023,0.29283017,0.19522011,0.09761006,0.0,0.1796025,0.359205,0.5388075,0.71841,0.9019169,0.76526284,0.62860876,0.4958591,0.359205,0.22645533,0.26940376,0.31625658,0.359205,0.40605783,0.44900626,0.6910792,0.92924774,1.1713207,1.4094892,1.6515622,2.4441557,3.2367494,4.029343,4.8219366,5.610626,6.434455,7.2582836,8.078208,8.902037,9.725866,9.323712,8.921559,8.519405,8.113348,7.7111945,8.652155,9.593117,10.534078,11.471134,12.412095,12.056794,11.697589,11.338385,10.983084,10.6238785,10.553599,10.479416,10.409137,10.334952,10.260769,10.4286585,10.592644,10.756628,10.920613,11.088503,10.510651,9.932799,9.354948,8.777096,8.1992445,8.36323,8.531119,8.695104,8.859089,9.023073,10.471607,11.916236,13.360865,14.805493,16.250122,17.53467,18.81922,20.103767,21.388315,22.67677,23.87542,25.074072,26.276627,27.475279,28.673931,28.759827,28.845724,28.931622,29.013613,29.09951,29.02923,28.955048,28.880863,28.810585,28.7364,30.423103,32.1059,33.792603,35.4793,37.1621,37.345608,37.53302,37.716526,37.90394,38.087444,38.345135,38.602825,38.860516,39.118206,39.375896,41.261723,43.143646,45.029472,46.9153,48.801125,52.98274,57.164352,61.34597,65.53149,69.713104,59.979427,50.249657,40.515984,30.782307,21.048632,18.089096,15.125654,12.162213,9.198771,6.239235,14.754736,23.266333,31.781834,40.297337,48.812836,45.388676,41.964516,38.53645,35.11229,31.68813,36.52178,41.359333,46.19298,51.026634,55.86419,58.975998,62.087803,65.199615,68.311424,71.42323,64.403114,57.386906,50.362885,43.346672,36.326557,33.433395,30.540234,27.647072,24.75391,21.860748,23.551353,25.238056,26.924759,28.61146,30.29816,29.954575,29.610987,29.263494,28.919907,28.57632,27.889145,27.201971,26.510891,25.823717,25.136541,27.420616,29.700788,31.984863,34.26894,36.54911,33.81993,31.090755,28.361578,25.628496,22.899319,23.570877,24.23853,24.910086,25.581644,26.249296,24.62116,22.98912,21.360985,19.728945,18.10081,18.366308,18.635712,18.90121,19.170614,19.436115,19.846077,20.252134,20.658192,21.068155,21.474213,20.412214,19.350218,18.28822,17.226223,16.164225,15.765976,15.371632,14.977287,14.582942,14.188598,14.313539,14.438479,14.56342,14.688361,14.813302,14.571229,14.33306,14.090988,13.852819,13.610746,13.263254,12.911859,12.564366,12.212971,11.861574,12.244205,12.626837,13.009468,13.392099,13.774731,14.063657,14.356487,14.645412,14.934339,15.223265,15.969006,16.714746,17.460487,18.206228,18.948065,18.928543,18.90902,18.889498,18.869976,18.850454,19.346313,19.838268,20.334127,20.829987,21.325846,21.247757,21.169668,21.091581,21.013493,20.93931,21.07206,21.208714,21.341463,21.478117,21.610867,21.778755,21.942741,22.106726,22.27071,22.4386,21.696764,20.958832,20.216995,19.479063,18.737226,18.600573,18.467823,18.33117,18.19842,18.061766,16.945107,15.828446,14.711788,13.591225,12.4745655,13.528754,14.586847,15.641035,16.695225,17.749413,16.796738,15.844065,14.89139,13.938716,12.986042,11.959184,10.928422,9.897659,8.866898,7.8361354,7.0630636,6.2938967,5.520825,4.747753,3.9746814,4.8687897,5.7668023,6.66091,7.5550184,8.449126,9.554072,10.655114,11.756155,12.861101,13.962143,0.8628729,0.8862993,0.9136301,0.93705654,0.96438736,0.9878138,0.9878138,0.9878138,0.9878138,0.9878138,0.9878138,0.999527,1.0112402,1.0268579,1.038571,1.0502841,1.0893283,1.1244678,1.1635119,1.1986516,1.2376955,1.2376955,1.2376955,1.2376955,1.2376955,1.2376955,1.261122,1.2884527,1.3118792,1.33921,1.3626363,1.3938715,1.4212024,1.4524376,1.4836729,1.5110037,1.620327,1.7257458,1.8350691,1.9443923,2.0498111,3.1977055,4.3455997,5.493494,6.6413884,7.7892823,10.502842,13.216402,15.933866,18.647425,21.360985,18.167183,14.973383,11.775677,8.581876,5.388075,4.4705405,3.5530062,2.6354716,1.717937,0.80040246,0.80040246,0.80040246,0.80040246,0.80040246,0.80040246,0.6910792,0.58566034,0.47633708,0.3709182,0.26159495,0.25378615,0.24597734,0.23816854,0.23426414,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.113227665,0.1717937,0.23035973,0.28892577,0.79649806,1.3079748,1.8194515,2.3270237,2.8385005,3.408543,3.9824903,4.5564375,5.12648,5.700427,6.262661,6.824895,7.387129,7.9493628,8.511597,9.097258,9.682918,10.268578,10.8542385,11.435994,11.209538,10.983084,10.756628,10.526268,10.299813,11.924045,13.544372,15.168603,16.788929,18.41316,17.546383,16.683512,15.816733,14.95386,14.087084,13.021181,11.959184,10.893282,9.82738,8.761478,8.074304,7.387129,6.699954,6.012779,5.3256044,5.5676775,5.8097506,6.0518236,6.2938967,6.5359693,6.98888,7.4417906,7.8947015,8.347612,8.800523,8.453031,8.105539,7.758047,7.4105554,7.0630636,6.8483214,6.6374836,6.426646,6.211904,6.001066,6.223617,6.4500723,6.676528,6.899079,7.125534,6.8678436,6.610153,6.3524623,6.094772,5.8370814,5.930787,6.028397,6.1221027,6.2158084,6.3134184,5.911265,5.5091114,5.1030536,4.7009,4.298747,4.290938,4.279225,4.271416,4.2597027,4.251894,4.376835,4.50568,4.630621,4.759466,4.8883114,5.3295093,5.7707067,6.2158084,6.657006,7.098203,7.387129,7.676055,7.9610763,8.250002,8.538928,8.441318,8.343708,8.246098,8.148487,8.050878,8.351517,8.648251,8.94889,9.249529,9.550168,8.987934,8.4257,7.8634663,7.3012323,6.7389984,8.058686,9.382278,10.705871,12.029464,13.349152,10.986988,8.624825,6.262661,3.900498,1.5383345,2.822883,4.1074314,5.3919797,6.676528,7.9610763,8.960603,9.964035,10.963562,11.963089,12.962616,13.325725,13.692739,14.055848,14.422862,14.785972,13.887959,12.986042,12.08803,11.186112,10.2881,9.854712,9.421323,8.991838,8.55845,8.125061,8.191436,8.261715,8.32809,8.3944645,8.460839,8.273428,8.082112,7.890797,7.703386,7.5120697,8.0040245,8.495979,8.991838,9.483793,9.975748,10.003078,10.03041,10.05774,10.085071,10.112402,11.490656,12.872814,14.251068,15.633226,17.01148,19.89293,22.770473,25.651922,28.533371,31.410915,29.829634,28.24835,26.663162,25.08188,23.500597,19.100336,14.700074,10.299813,5.899552,1.4992905,1.1986516,0.9019169,0.60127795,0.30063897,0.0,0.26549935,0.5309987,0.79649806,1.0580931,1.3235924,3.2016098,5.0796275,6.957645,8.835662,10.71368,12.86891,15.024139,17.17937,19.330696,21.485926,22.50107,23.51231,24.52355,25.538694,26.549934,22.85637,19.158901,15.465338,11.771772,8.074304,8.449126,8.823949,9.198771,9.573594,9.948417,9.971844,9.99527,10.018696,10.0382185,10.061645,10.151445,10.241247,10.331048,10.42085,10.510651,9.741484,8.972317,8.203149,7.433982,6.66091,6.532065,6.4032197,6.2743745,6.141625,6.012779,6.4969254,6.9771667,7.461313,7.941554,8.4257,9.01136,9.593117,10.178777,10.764437,11.350098,11.279819,11.209538,11.139259,11.06898,10.998701,9.82738,8.65606,7.480835,6.309514,5.138193,5.35684,5.579391,5.7980375,6.016684,6.239235,5.446641,4.657952,3.8692627,3.076669,2.2879796,1.9209659,1.5539521,1.1869383,0.8160201,0.44900626,0.359205,0.26940376,0.1796025,0.08980125,0.0,0.12103647,0.23816854,0.359205,0.48024148,0.60127795,0.5114767,0.42167544,0.3318742,0.23816854,0.14836729,0.19131571,0.23426414,0.27721256,0.32016098,0.3631094,0.6481308,0.93315214,1.2181735,1.5031948,1.7882162,2.358259,2.9283018,3.4983444,4.068387,4.6384296,5.263134,5.891743,6.520352,7.1489606,7.773665,7.3910336,7.0044975,6.621866,6.2353306,5.8487945,6.5359693,7.2192397,7.9064145,8.589685,9.276859,8.98403,8.691199,8.398369,8.105539,7.812709,8.183627,8.55845,8.929368,9.304191,9.675109,9.647778,9.620447,9.593117,9.565785,9.538455,8.991838,8.441318,7.8947015,7.348085,6.801469,7.1333427,7.4691215,7.8049,8.140678,8.476458,9.815667,11.158782,12.501896,13.845011,15.188125,16.39068,17.593237,18.795792,19.998348,21.200905,21.888079,22.575254,23.262428,23.949604,24.636778,24.976461,25.316145,25.655827,25.999414,26.339098,26.448421,26.557745,26.667067,26.77639,26.885714,27.740778,28.591938,29.447002,30.29816,31.14932,31.789642,32.429966,33.070286,33.71061,34.35093,35.904884,37.458836,39.016693,40.570644,42.124596,43.80349,45.478477,47.15737,48.83626,50.511253,52.71724,54.923225,57.129215,59.331295,61.537285,53.068634,44.60389,36.135242,27.666594,19.20185,16.937298,14.676648,12.412095,10.151445,7.8868923,15.621513,23.356134,31.09466,38.82928,46.5639,44.57656,42.58922,40.597973,38.610634,36.623295,41.753677,46.880157,52.006638,57.133118,62.263504,62.013622,61.76374,61.51386,61.263977,61.014095,54.743626,48.47706,42.21049,35.943928,29.673458,29.443098,29.208834,28.978474,28.74421,28.51385,30.5988,32.687656,34.776512,36.86146,38.950317,36.943455,34.940495,32.93363,30.930676,28.923813,28.486519,28.049225,27.611933,27.17464,26.737347,28.267872,29.798397,31.328924,32.85945,34.38607,32.23084,30.071707,27.916475,25.757341,23.598207,24.87885,26.159494,27.44014,28.720783,30.001427,27.881336,25.761246,23.641155,21.521065,19.400974,19.756275,20.11548,20.470781,20.829987,21.189192,21.681147,22.1731,22.665054,23.15701,23.648964,22.024733,20.400501,18.77627,17.152039,15.523903,15.418485,15.313066,15.211552,15.1061325,15.000713,15.336493,15.676175,16.011953,16.351637,16.687416,16.39068,16.093946,15.793307,15.4965725,15.199838,14.473619,13.751305,13.025085,12.298867,11.576552,11.916236,12.259823,12.603411,12.943093,13.286681,13.360865,13.431144,13.505327,13.575606,13.64979,14.090988,14.53609,14.977287,15.418485,15.863586,16.359446,16.8514,17.34726,17.843119,18.338978,19.041769,19.748466,20.45126,21.157955,21.860748,21.688955,21.51716,21.345367,21.173573,21.00178,21.00178,21.005684,21.005684,21.009588,21.013493,21.349272,21.681147,22.016924,22.352703,22.688482,22.04035,21.39222,20.74409,20.095959,19.451733,19.20966,18.97149,18.729418,18.49125,18.249176,17.316025,16.386776,15.453624,14.520472,13.58732,14.356487,15.125654,15.8987255,16.667892,17.437061,16.539047,15.641035,14.743023,13.848915,12.950902,12.2793455,11.611692,10.940135,10.268578,9.600925,8.609207,7.621393,6.629675,5.6418614,4.650143,5.493494,6.336845,7.1762915,8.019642,8.862993,9.796145,10.733202,11.666354,12.603411,13.536563,0.9019169,0.92534333,0.94876975,0.97610056,0.999527,1.0268579,1.0268579,1.0268579,1.0268579,1.0268579,1.0268579,1.038571,1.0502841,1.0619974,1.0737107,1.0893283,1.1361811,1.1869383,1.2376955,1.2884527,1.33921,1.3235924,1.3118792,1.3001659,1.2884527,1.2767396,1.3001659,1.3235924,1.3509232,1.3743496,1.4016805,1.4133936,1.4290112,1.4446288,1.4602464,1.475864,1.5110037,1.5461433,1.5812829,1.6164225,1.6515622,3.06886,4.4861584,5.903456,7.320754,8.738052,11.045554,13.353056,15.660558,17.96806,20.27556,17.128613,13.981665,10.8308115,7.6838636,4.5369153,3.7989833,3.057147,2.3192148,1.5773785,0.8394465,0.81211567,0.78868926,0.76135844,0.737932,0.7106012,0.61689556,0.5192855,0.42167544,0.3240654,0.22645533,0.21474212,0.20693332,0.19522011,0.1835069,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.75354964,1.3353056,1.9131571,2.494913,3.076669,3.619381,4.1581883,4.7009,5.2436123,5.786324,6.364176,6.9381227,7.5120697,8.086017,8.663869,9.354948,10.046027,10.741011,11.43209,12.123169,11.642927,11.158782,10.67854,10.194394,9.714153,11.166591,12.622932,14.079274,15.531713,16.988054,16.179844,15.371632,14.56342,13.759113,12.950902,11.806912,10.6590185,9.515028,8.371038,7.223144,6.774138,6.3251314,5.8761253,5.423215,4.9742084,5.466163,5.9542136,6.446168,6.9342184,7.426173,7.8205175,8.214863,8.609207,9.0035515,9.4018,8.781001,8.164105,7.5472097,6.930314,6.3134184,6.13772,5.9620223,5.786324,5.610626,5.4388323,5.8487945,6.262661,6.676528,7.08649,7.5003567,7.141152,6.7819467,6.4188375,6.0596323,5.700427,5.4856853,5.270943,5.056201,4.841459,4.6267166,4.478349,4.3338866,4.1894236,4.044961,3.900498,3.8965936,3.8887846,3.8848803,3.8809757,3.873167,4.084005,4.290938,4.4978714,4.704805,4.911738,5.364649,5.8175592,6.27047,6.7233806,7.1762915,7.5120697,7.8517528,8.187531,8.52331,8.862993,8.734148,8.601398,8.472553,8.343708,8.210958,8.335898,8.460839,8.58578,8.710721,8.835662,8.4257,8.011833,7.601871,7.1880045,6.774138,7.8556576,8.933272,10.0147915,11.096312,12.173926,10.151445,8.125061,6.098676,4.0761957,2.0498111,3.3187418,4.5837684,5.852699,7.1216297,8.386656,9.386183,10.38571,11.389141,12.388668,13.388195,14.0831785,14.778163,15.473146,16.168129,16.863113,15.726933,14.586847,13.450665,12.31058,11.174399,10.666827,10.155351,9.643873,9.136301,8.624825,8.75367,8.878611,9.007456,9.136301,9.261242,8.991838,8.722435,8.453031,8.183627,7.914223,8.402273,8.894228,9.382278,9.874233,10.362284,10.42085,10.479416,10.534078,10.592644,10.651209,12.103647,13.556085,15.008522,16.46096,17.913397,20.990067,24.066736,27.143404,30.223978,33.300648,30.778402,28.256159,25.733915,23.211672,20.685524,16.863113,13.036799,9.2104845,5.388075,1.5617609,1.2494087,0.93705654,0.62470436,0.31235218,0.0,0.3318742,0.6637484,0.9956226,1.3314011,1.6632754,3.619381,5.579391,7.535496,9.491602,11.4516115,13.2788725,15.1061325,16.933393,18.760653,20.587914,20.911978,21.236044,21.564014,21.888079,22.212145,18.928543,15.641035,12.357433,9.073831,5.786324,6.899079,8.011833,9.124588,10.237343,11.350098,10.990892,10.6355915,10.276386,9.921086,9.561881,9.921086,10.276386,10.6355915,10.990892,11.350098,10.553599,9.753197,8.956698,8.160201,7.363703,7.1489606,6.9342184,6.715572,6.5008297,6.2860875,6.6960497,7.1060123,7.5159745,7.9259367,8.335898,8.941081,9.546264,10.151445,10.756628,11.361811,11.053363,10.741011,10.432563,10.124115,9.811763,9.120684,8.4257,7.734621,7.043542,6.348558,6.7233806,7.094299,7.4691215,7.8400397,8.210958,6.8405128,5.473972,4.1035266,2.7330816,1.3626363,1.1713207,0.98390937,0.79259366,0.60127795,0.41386664,0.3318742,0.24597734,0.1639849,0.08199245,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.25378615,0.21083772,0.1639849,0.12103647,0.07418364,0.113227665,0.15617609,0.19522011,0.23426414,0.27330816,0.60518235,0.93315214,1.2650263,1.5969005,1.9248703,2.2723622,2.619854,2.9673457,3.3148375,3.6623292,4.095718,4.5291066,4.958591,5.3919797,5.825368,5.4583545,5.0913405,4.7243266,4.3534083,3.9863946,4.415879,4.8492675,5.278752,5.708236,6.13772,5.911265,5.6809053,5.45445,5.2279944,5.001539,5.8175592,6.6335793,7.453504,8.269524,9.085544,8.866898,8.648251,8.4257,8.207053,7.988407,7.4691215,6.9537406,6.434455,5.919074,5.3997884,5.903456,6.4110284,6.914696,7.4183645,7.9259367,9.163632,10.405232,11.6468315,12.884527,14.126127,15.246691,16.36335,17.483913,18.604477,5052.0,19.900738,20.076437,20.24823,20.423927,20.599627,21.193096,21.790468,22.383938,22.981312,23.574781,23.86761,24.16044,24.453272,24.746101,25.03893,25.058455,25.077976,25.097498,25.11702,25.136541,26.233679,27.326912,28.42405,29.51728,30.610514,33.46463,36.31875,39.168964,42.023083,44.873295,46.345253,47.81331,49.28527,50.753326,52.225285,52.45174,52.678196,52.908554,53.13501,53.361465,46.157845,38.958126,31.754503,24.55088,17.351164,15.785499,14.223738,12.661977,11.100216,9.538455,16.492195,23.445936,30.40358,37.357323,44.31106,43.76054,43.213924,42.663403,42.112885,41.562363,46.981674,52.40098,57.824196,63.243507,68.66282,65.05125,61.43577,57.824196,54.212624,50.60105,45.084133,39.571117,34.054195,28.54118,23.02426,25.452799,27.881336,30.305971,32.73451,35.163048,37.65015,40.137257,42.62436,45.111465,47.598568,43.936237,40.270004,36.60377,32.94144,29.275208,29.087797,28.900385,28.712975,28.525562,28.338152,29.115128,29.892103,30.669079,31.446056,32.22303,30.641748,29.056562,27.471375,25.886187,24.300999,26.190731,28.080462,29.970192,31.859922,33.749653,31.141512,28.529467,25.921326,23.309282,20.701141,21.146242,21.59525,22.044254,22.489357,22.938364,23.516214,24.094067,24.671917,25.245865,25.823717,23.63725,21.450787,19.26432,17.073952,14.8874855,15.070992,15.258404,15.441911,15.629322,15.812829,16.36335,16.91387,17.464392,18.011007,18.56153,18.206228,17.850927,17.495626,17.14423,16.788929,15.687888,14.586847,13.4858055,12.388668,11.287627,11.588266,11.892809,12.193448,12.497992,12.798631,12.654168,12.509705,12.365242,12.220779,12.076316,12.216875,12.353529,12.494087,12.634645,12.775204,13.786445,14.79378,15.80502,16.816261,17.823597,18.74113,19.65476,20.568392,21.485926,22.399555,22.134056,21.864653,21.599154,21.32975,21.06425,20.931501,20.802654,20.67381,20.54106,20.412214,20.915882,21.423454,21.927124,22.430792,22.938364,22.383938,21.82561,21.271183,20.716759,20.162333,19.818747,19.471254,19.127666,18.784079,18.436588,17.690847,16.941202,16.195461,15.445815,14.700074,15.18422,15.668366,16.156416,16.640562,17.124708,16.281357,15.438006,14.59856,13.755209,12.911859,12.603411,12.291059,11.982611,11.674163,11.361811,10.155351,8.94889,7.7385254,6.532065,5.3256044,6.114294,6.9068875,7.6955767,8.484266,9.276859,10.042123,10.81129,11.576552,12.34572,13.110983,0.93705654,0.96438736,0.9878138,1.0112402,1.038571,1.0619974,1.0619974,1.0619974,1.0619974,1.0619974,1.0619974,1.0737107,1.0893283,1.1010414,1.1127546,1.1244678,1.1869383,1.2494087,1.3118792,1.3743496,1.43682,1.4133936,1.3860629,1.3626363,1.33921,1.3118792,1.33921,1.3626363,1.3860629,1.4133936,1.43682,1.43682,1.43682,1.43682,1.43682,1.43682,1.4016805,1.3626363,1.3235924,1.2884527,1.2494087,2.9361105,4.6267166,6.3134184,8.00012,9.686822,11.588266,13.4858055,15.387249,17.288692,19.186234,16.086138,12.986042,9.885946,6.785851,3.6857557,3.1235218,2.5612879,1.999054,1.43682,0.8745861,0.8238289,0.77307165,0.7262188,0.6754616,0.62470436,0.5388075,0.44900626,0.3631094,0.27330816,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.7106012,1.3626363,2.0107672,2.6628022,3.310933,3.8263142,4.337791,4.8492675,5.3607445,5.8761253,6.461786,7.0513506,7.6370106,8.226576,8.812236,9.612638,10.413041,11.213444,12.013845,12.814248,12.076316,11.338385,10.600452,9.86252,9.124588,10.413041,11.701493,12.986042,14.274494,15.562947,14.813302,14.063657,13.314012,12.564366,11.810817,10.588739,9.362757,8.136774,6.910792,5.688714,5.473972,5.263134,5.0483923,4.8375545,4.6267166,5.3607445,6.098676,6.8366084,7.57454,8.312472,8.648251,8.987934,9.323712,9.663396,9.999174,9.112875,8.226576,7.336372,6.4500723,5.563773,5.423215,5.2865605,5.1499066,5.0132523,4.8765984,5.473972,6.0752497,6.676528,7.2739015,7.8751793,7.4105554,6.949836,6.4891167,6.0244927,5.563773,5.036679,4.513489,3.9863946,3.4632049,2.9361105,3.049338,3.1625657,3.2757936,3.3890212,3.4983444,3.4983444,3.4983444,3.4983444,3.4983444,3.4983444,3.78727,4.0761957,4.3612175,4.650143,4.939069,5.3997884,5.8644123,6.3251314,6.785851,7.250475,7.6370106,8.023546,8.413987,8.800523,9.187058,9.023073,8.862993,8.699008,8.538928,8.374943,8.324185,8.273428,8.226576,8.175818,8.125061,7.8634663,7.601871,7.336372,7.0747766,6.813182,7.648724,8.488171,9.323712,10.163159,10.998701,9.311999,7.6252975,5.938596,4.251894,2.5612879,3.8106966,5.0640097,6.3134184,7.562827,8.812236,9.811763,10.81129,11.810817,12.814248,13.813775,14.836729,15.863586,16.88654,17.913397,18.936352,17.562002,16.187653,14.813302,13.438952,12.0606985,11.475039,10.889378,10.299813,9.714153,9.124588,9.311999,9.499411,9.686822,9.874233,10.061645,9.714153,9.362757,9.01136,8.663869,8.312472,8.800523,9.288573,9.776623,10.260769,10.748819,10.838621,10.924518,11.014318,11.100216,11.186112,12.712734,14.239355,15.762072,17.288692,18.81141,22.087204,25.362997,28.63879,31.910679,35.186474,31.723269,28.263968,24.800762,21.337559,17.874353,14.625891,11.373524,8.125061,4.8765984,1.6242313,1.3001659,0.97610056,0.6481308,0.3240654,0.0,0.39824903,0.80040246,1.1986516,1.6008049,1.999054,4.037152,6.0752497,8.113348,10.151445,12.185639,13.688834,15.188125,16.687416,18.186707,19.685997,19.326792,18.963682,18.600573,18.237463,17.874353,15.000713,12.123169,9.249529,6.375889,3.4983444,5.349031,7.1997175,9.050405,10.901091,12.751778,12.013845,11.275913,10.537982,9.80005,9.062118,9.686822,10.311526,10.936231,11.560935,12.185639,11.361811,10.537982,9.714153,8.886419,8.062591,7.7619514,7.461313,7.1606736,6.8639393,6.5633,6.899079,7.238762,7.57454,7.914223,8.250002,8.874706,9.499411,10.124115,10.748819,11.373524,10.826907,10.276386,9.725866,9.175345,8.624825,8.413987,8.1992445,7.988407,7.773665,7.562827,8.086017,8.6131115,9.136301,9.663396,10.186585,8.238289,6.2860875,4.337791,2.3855898,0.43729305,0.42557985,0.41386664,0.39824903,0.38653582,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.5622339,0.93705654,1.3118792,1.6867018,2.0615244,2.1864653,2.3114061,2.436347,2.5612879,2.6862288,2.9243972,3.1625657,3.4007344,3.638903,3.873167,3.5256753,3.174279,2.8267872,2.475391,2.1239948,2.2996929,2.475391,2.6510892,2.8267872,2.998581,2.8385005,2.6745155,2.514435,2.35045,2.1864653,3.4514916,4.7126136,5.9737353,7.238762,8.499884,8.086017,7.676055,7.262188,6.8483214,6.4383593,5.950309,5.462259,4.9742084,4.4861584,3.998108,4.6735697,5.349031,6.0244927,6.699954,7.375416,8.511597,9.651682,10.787864,11.924045,13.06413,14.098797,15.137367,16.175938,17.210606,18.249176,17.913397,17.573715,17.237936,16.898252,16.562475,17.413633,18.26089,19.11205,19.96321,20.81437,21.2868,21.763138,22.23557,22.711908,23.188246,22.37613,21.564014,20.751898,19.935879,19.123762,20.67381,22.223858,23.773905,25.323954,26.874,31.02438,35.17476,39.325138,43.475517,47.6259,48.88702,50.148144,51.41317,52.67429,53.939316,52.18624,50.43707,48.687897,46.938725,45.185646,39.250957,33.31236,27.373764,21.439074,15.500477,14.637604,13.774731,12.911859,12.0489855,11.186112,17.362877,23.535736,29.712502,35.889267,42.062126,42.948425,43.838627,44.724926,45.61123,46.50143,52.21357,57.925713,63.63785,69.34999,75.06213,68.08887,61.111706,54.138443,47.161274,40.18801,35.42464,30.66127,25.901804,21.138433,16.375063,21.4625,26.549934,31.637371,36.724808,41.812244,44.7015,47.586853,50.476112,53.361465,56.250725,50.925117,45.599514,40.27391,34.948303,29.626604,29.689075,29.751545,29.814016,29.876486,29.938957,29.962383,29.98581,30.01314,30.036566,30.063898,29.048752,28.037512,27.026272,26.011127,24.999887,27.498705,30.001427,32.500244,34.99906,37.501785,34.401688,31.301594,28.201498,25.101402,22.001307,22.53621,23.075018,23.613825,24.148727,24.687536,25.351284,26.011127,26.674877,27.338625,27.998468,25.24977,22.50107,19.748466,16.999767,14.251068,14.723501,15.199838,15.676175,16.148607,16.624945,17.386303,18.151566,18.912924,19.674282,20.435642,20.025679,19.611813,19.20185,18.787983,18.374117,16.898252,15.426293,13.950429,12.4745655,10.998701,11.2642,11.525795,11.787391,12.0489855,12.31058,11.951375,11.588266,11.225157,10.862047,10.498938,10.338858,10.174872,10.010887,9.850807,9.686822,11.213444,12.73616,14.262781,15.785499,17.31212,18.436588,19.561056,20.689428,21.813896,22.938364,22.575254,22.212145,21.849035,21.485926,21.12672,20.861221,20.599627,20.338032,20.076437,19.810938,20.486399,21.16186,21.837322,22.512783,23.188246,22.723621,22.262901,21.798277,21.337559,20.876839,20.423927,19.974922,19.525915,19.07691,18.623999,18.061766,17.49953,16.937298,16.375063,15.812829,16.011953,16.211079,16.414106,16.613232,16.812357,16.023666,15.238882,14.450192,13.661504,12.8767185,12.923572,12.974329,13.025085,13.075843,13.1266,11.701493,10.276386,8.85128,7.426173,6.001066,6.7389984,7.47693,8.210958,8.94889,9.686822,10.2881,10.889378,11.486752,12.08803,12.689307,0.999527,1.0190489,1.038571,1.0580931,1.0815194,1.1010414,1.1049459,1.1088502,1.116659,1.1205635,1.1244678,1.1478943,1.1713207,1.1908426,1.2142692,1.2376955,1.2728351,1.3079748,1.3431144,1.3782539,1.4133936,1.4016805,1.3938715,1.3821584,1.3743496,1.3626363,1.3743496,1.3860629,1.4016805,1.4133936,1.4251068,1.4133936,1.4016805,1.3860629,1.3743496,1.3626363,1.3118792,1.261122,1.2142692,1.1635119,1.1127546,3.6857557,6.262661,8.835662,11.412568,13.985569,14.438479,14.89139,15.344301,15.797212,16.250122,13.68493,11.119738,8.554545,5.989353,3.4241607,2.893162,2.358259,1.8272603,1.2962615,0.76135844,0.7262188,0.6871748,0.6481308,0.61299115,0.57394713,0.5036679,0.43338865,0.3631094,0.29673457,0.22645533,0.20302892,0.1796025,0.15617609,0.13665408,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.57394713,1.1010414,1.6242313,2.1513257,2.6745155,3.2055142,3.736513,4.263607,4.794606,5.3256044,5.883934,6.446168,7.0044975,7.5667315,8.125061,8.913751,9.698535,10.487225,11.275913,12.0606985,11.400854,10.737106,10.073358,9.413514,8.749765,9.663396,10.58093,11.49456,12.408191,13.325725,12.658072,11.994324,11.330575,10.666827,9.999174,9.21439,8.429605,7.6448197,6.860035,6.0752497,6.0713453,6.0635366,6.0596323,6.055728,6.0518236,6.7663293,7.4847393,8.203149,8.921559,9.636065,9.86252,10.088976,10.311526,10.537982,10.764437,9.811763,8.862993,7.914223,6.9615493,6.012779,5.883934,5.7511845,5.6223392,5.493494,5.3607445,5.840986,6.3173227,6.79366,7.2739015,7.7502384,7.3832245,7.0201154,6.6531014,6.289992,5.9268827,5.3138914,4.704805,4.095718,3.4866312,2.87364,3.049338,3.2250361,3.4007344,3.5764325,3.7482262,3.7521305,3.7560349,3.7560349,3.7599394,3.7638438,3.998108,4.2323723,4.466636,4.7009,4.939069,5.388075,5.840986,6.2938967,6.746807,7.1997175,7.558923,7.914223,8.273428,8.628729,8.987934,8.784905,8.581876,8.378847,8.175818,7.9766936,7.8868923,7.793187,7.703386,7.6135845,7.523783,7.426173,7.3246584,7.223144,7.125534,7.0240197,7.5979667,8.171914,8.741957,9.315904,9.885946,8.468649,7.0513506,5.6340523,4.2167544,2.7994564,4.1035266,5.4036927,6.707763,8.011833,9.311999,10.100689,10.889378,11.674163,12.4628525,13.251541,14.008995,14.770353,15.531713,16.289165,17.050524,15.851873,14.649317,13.450665,12.24811,11.0494585,10.631687,10.2100115,9.788337,9.370565,8.94889,9.218294,9.491602,9.761005,10.03041,10.299813,10.0382185,9.776623,9.511124,9.249529,8.987934,9.296382,9.600925,9.909373,10.217821,10.526268,10.721489,10.920613,11.115833,11.314958,11.514082,13.903577,16.29307,18.682566,21.07206,23.461554,25.476225,27.490896,29.509472,31.524143,33.538815,29.829634,26.124355,22.415173,18.705992,15.000713,12.302772,9.60483,6.9068875,4.2089458,1.5110037,1.2494087,0.9878138,0.7262188,0.46071947,0.19912452,0.57394713,0.94876975,1.3235924,1.698415,2.0732377,3.7443218,5.4154058,7.08649,8.75367,10.424754,12.236397,14.048039,15.863586,17.675228,19.486872,19.29165,19.096432,18.90121,18.705992,18.51077,16.03538,13.556085,11.080693,8.601398,6.126007,7.3168497,8.503788,9.694631,10.885473,12.076316,11.256392,10.4403715,9.6243515,8.804427,7.988407,8.624825,9.261242,9.901564,10.537982,11.174399,10.475512,9.780528,9.081639,8.386656,7.687768,7.480835,7.2739015,7.0630636,6.8561306,6.649197,6.984976,7.320754,7.656533,7.988407,8.324185,8.777096,9.230007,9.682918,10.135828,10.588739,10.198298,9.807858,9.4174185,9.026978,8.636538,8.39056,8.148487,7.90251,7.656533,7.4105554,8.109444,8.804427,9.499411,10.194394,10.889378,8.894228,6.899079,4.903929,2.9087796,0.9136301,0.79649806,0.679366,0.5583295,0.44119745,0.3240654,0.26159495,0.19522011,0.12884527,0.06637484,0.0,0.0,0.0,0.0,0.0,0.0,0.042948425,0.08589685,0.12884527,0.1717937,0.21083772,0.26940376,0.3240654,0.37872702,0.43338865,0.48805028,0.8706817,1.2572175,1.6437533,2.0263848,2.4129205,2.475391,2.5378613,2.6003318,2.6628022,2.7252727,2.8853533,3.0454338,3.2055142,3.3655949,3.5256753,3.2094188,2.893162,2.5808098,2.2645533,1.9482968,2.077142,2.2059872,2.330928,2.4597735,2.5886188,2.5027218,2.416825,2.330928,2.2489357,2.1630387,3.3070288,4.4510183,5.5989127,6.7429028,7.8868923,7.5550184,7.223144,6.89127,6.559396,6.223617,5.677001,5.1303844,4.5837684,4.0332475,3.4866312,4.1464753,4.802415,5.4583545,6.1181984,6.774138,8.054782,9.335425,10.61607,11.896713,13.173453,13.813775,14.450192,15.086611,15.726933,16.36335,16.183748,16.004145,15.820638,15.641035,15.461433,16.617136,17.772839,18.928543,20.084246,21.236044,21.118912,20.997875,20.876839,20.755802,20.63867,20.166237,19.69771,19.229181,18.756748,18.28822,20.201378,22.118439,24.031595,25.948658,27.861814,31.816975,35.76823,39.719482,43.67074,47.6259,48.55905,49.49611,50.42926,51.366318,52.29947,50.52687,48.754272,46.981674,45.209072,43.436474,37.646248,31.852114,26.057981,20.267752,14.473619,13.895767,13.314012,12.73616,12.154405,11.576552,16.375063,21.173573,25.975988,30.774498,35.576912,36.377316,37.18162,37.982025,38.78633,39.586735,44.412575,49.23842,54.06426,58.886196,63.712036,57.874954,52.037872,46.20079,40.363712,34.52663,31.243027,27.96333,24.683632,21.403933,18.124235,22.559637,26.991133,31.42263,35.854126,40.28562,42.72197,45.158318,47.59076,50.027107,52.46345,47.61809,42.77663,37.935173,33.09371,28.24835,28.287394,28.326439,28.361578,28.400621,28.435762,28.369387,28.299107,28.228828,28.158548,28.08827,27.447948,26.807627,26.167303,25.526981,24.88666,26.94428,28.997995,31.051712,33.10933,35.163048,32.48072,29.798397,27.116074,24.43375,21.751425,22.27071,22.789995,23.309282,23.828568,24.351757,24.48841,24.62897,24.769527,24.910086,25.050644,22.67677,20.306797,17.93292,15.559043,13.189071,13.821584,14.458001,15.0944195,15.726933,16.36335,17.042715,17.722082,18.401447,19.080814,19.764084,19.283842,18.8036,18.32336,17.843119,17.362877,16.316498,15.274021,14.227642,13.181262,12.138786,12.2793455,12.415999,12.556558,12.697116,12.837675,12.349625,11.861574,11.373524,10.889378,10.401327,10.459893,10.518459,10.58093,10.639496,10.698062,12.006037,13.310107,14.614178,15.918248,17.226223,18.54591,19.865599,21.185287,22.504974,23.824663,23.461554,23.09454,22.73143,22.364416,22.001307,21.548395,21.095486,20.642574,20.189665,19.736753,20.423927,21.111103,21.798277,22.489357,23.176533,22.821232,22.46593,22.11063,21.75533,21.400028,20.986162,20.568392,20.154524,19.740658,19.326792,18.791887,18.25308,17.718178,17.183275,16.64837,16.952915,17.253553,17.558098,17.858736,18.163279,17.101282,16.039284,14.973383,13.911386,12.849388,12.728352,12.611219,12.490183,12.369146,12.24811,11.084598,9.921086,8.75367,7.590158,6.426646,7.0630636,7.699481,8.335898,8.976221,9.612638,10.2334385,10.858143,11.478943,12.103647,12.724447,1.0619974,1.077615,1.0932326,1.1088502,1.1205635,1.1361811,1.1478943,1.1557031,1.1674163,1.1791295,1.1869383,1.2181735,1.2533131,1.2845483,1.3157835,1.3509232,1.358732,1.3665408,1.3743496,1.3782539,1.3860629,1.3938715,1.397776,1.4016805,1.4055848,1.4133936,1.4133936,1.4133936,1.4133936,1.4133936,1.4133936,1.3860629,1.3626363,1.33921,1.3118792,1.2884527,1.2259823,1.1635119,1.1010414,1.038571,0.97610056,4.4393053,7.898606,11.361811,14.825015,18.28822,17.292597,16.296974,15.3013525,14.30573,13.314012,11.283723,9.253433,7.223144,5.192855,3.1625657,2.6588979,2.1591344,1.6554666,1.1517987,0.6481308,0.62470436,0.60127795,0.57394713,0.5505207,0.5231899,0.47243267,0.42167544,0.3670138,0.31625658,0.26159495,0.23035973,0.19912452,0.1639849,0.13274968,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.43729305,0.8355421,1.2376955,1.6359446,2.0380979,2.5847144,3.1313305,3.6818514,4.2284675,4.775084,5.3060827,5.840986,6.3719845,6.9068875,7.437886,8.210958,8.987934,9.761005,10.537982,11.311053,10.725393,10.135828,9.550168,8.960603,8.374943,8.917655,9.460366,10.003078,10.545791,11.088503,10.506746,9.928895,9.347139,8.769287,8.187531,7.843944,7.4964523,7.152865,6.8092775,6.461786,6.6648145,6.8678436,7.0708723,7.2739015,7.47693,8.171914,8.870802,9.565785,10.264673,10.963562,11.076789,11.186112,11.29934,11.412568,11.525795,10.510651,9.499411,8.488171,7.47693,6.461786,6.3407493,6.2158084,6.094772,5.9737353,5.8487945,6.2040954,6.559396,6.914696,7.269997,7.6252975,7.355894,7.0903945,6.8209906,6.5554914,6.2860875,5.591104,4.8961205,4.2011366,3.506153,2.8111696,3.049338,3.2875066,3.5256753,3.7638438,3.998108,4.0059166,4.009821,4.0137253,4.0215344,4.025439,4.2089458,4.388548,4.572055,4.755562,4.939069,5.380266,5.8214636,6.266566,6.707763,7.1489606,7.47693,7.8049,8.13287,8.460839,8.78881,8.546737,8.300759,8.058686,7.816613,7.57454,7.445695,7.3168497,7.1841,7.055255,6.9264097,6.98888,7.0513506,7.113821,7.1762915,7.238762,7.5433054,7.8517528,8.160201,8.468649,8.773191,7.629202,6.481308,5.3334136,4.185519,3.0376248,4.3924527,5.74728,7.1021075,8.456935,9.811763,10.38571,10.963562,11.537509,12.111456,12.689307,13.181262,13.677121,14.17298,14.668839,15.160794,14.13784,13.110983,12.08803,11.061172,10.0382185,9.784432,9.530646,9.280765,9.026978,8.773191,9.128492,9.479889,9.8312845,10.186585,10.537982,10.362284,10.186585,10.010887,9.839094,9.663396,9.788337,9.917182,10.046027,10.170968,10.299813,10.608261,10.916709,11.221252,11.5297,11.838148,15.090515,18.346786,21.603058,24.85933,28.111696,28.86915,29.6227,30.37625,31.133703,31.887253,27.935999,23.980839,20.029583,16.07833,12.123169,9.979652,7.8361354,5.688714,3.5451972,1.4016805,1.1986516,0.999527,0.80040246,0.60127795,0.39824903,0.74964523,1.1010414,1.4485333,1.7999294,2.1513257,3.4514916,4.755562,6.055728,7.3597984,8.663869,10.787864,12.911859,15.035853,17.163752,19.287746,19.260416,19.233086,19.205755,19.178425,19.151093,17.070047,14.989,12.911859,10.8308115,8.749765,9.280765,9.811763,10.338858,10.869856,11.400854,10.502842,9.60483,8.706817,7.8088045,6.910792,7.562827,8.210958,8.862993,9.511124,10.163159,9.593117,9.023073,8.453031,7.882988,7.3129454,7.195813,7.082586,6.969358,6.852226,6.7389984,7.0708723,7.4027467,7.734621,8.066495,8.398369,8.679486,8.960603,9.24172,9.518932,9.80005,9.56969,9.339331,9.108971,8.878611,8.648251,8.371038,8.093826,7.816613,7.5394006,7.262188,8.128965,8.991838,9.858616,10.721489,11.588266,9.546264,7.5081654,5.466163,3.4280653,1.3860629,1.1635119,0.94096094,0.71841,0.4958591,0.27330816,0.21864653,0.1639849,0.10932326,0.05466163,0.0,0.0,0.0,0.0,0.0,0.0,0.08589685,0.1717937,0.25378615,0.339683,0.42557985,0.4958591,0.5700427,0.6442264,0.7145056,0.78868926,1.183034,1.5773785,1.9717231,2.366068,2.7643168,2.7643168,2.7643168,2.7643168,2.7643168,2.7643168,2.8463092,2.9283018,3.0102942,3.0922866,3.174279,2.893162,2.6159496,2.3348327,2.0537157,1.7765031,1.8545911,1.9365835,2.0146716,2.096664,2.174752,2.1669433,2.1591344,2.1513257,2.1435168,2.135708,3.1664703,4.193328,5.2201858,6.2470436,7.2739015,7.0240197,6.7702336,6.5164475,6.266566,6.012779,5.4036927,4.7985106,4.1894236,3.5842414,2.9751544,3.6154766,4.2557983,4.8961205,5.5364423,6.1767645,7.5979667,9.019169,10.444276,11.8654785,13.286681,13.524849,13.763018,14.001186,14.239355,14.473619,14.454097,14.430671,14.407245,14.383818,14.364296,15.820638,17.280884,18.74113,20.201378,21.661623,20.947119,20.232613,19.518106,18.8036,18.089096,17.96025,17.831406,17.706465,17.57762,17.448774,19.728945,22.009115,24.289286,26.569458,28.849628,32.605663,36.3617,40.11383,43.869865,47.6259,48.231083,48.840168,49.449253,50.054436,50.663525,48.8675,47.071472,45.279354,43.48333,41.6873,36.04154,30.391867,24.746101,19.096432,13.450665,13.153932,12.853292,12.556558,12.259823,11.963089,15.387249,18.81141,22.239475,25.663635,29.087797,29.806208,30.520712,31.239122,31.957533,32.67594,36.61158,40.55112,44.48676,48.4263,52.36194,47.661037,42.964043,38.26314,33.56224,28.861341,27.065317,25.26929,23.469362,21.673336,19.873407,23.652868,27.428427,31.207888,34.983444,38.762905,40.74634,42.725872,44.70931,46.692745,48.67618,44.314964,39.953747,35.596436,31.235218,26.874,26.885714,26.90133,26.913044,26.924759,26.936472,26.772486,26.608501,26.440613,26.276627,26.112642,25.843239,25.57774,25.308336,25.042835,24.773432,26.38595,27.994564,29.603178,31.215696,32.82431,30.559757,28.295202,26.03065,23.766096,21.501543,22.001307,22.504974,23.008642,23.508406,24.012074,23.629442,23.24681,22.86418,22.481548,22.098917,20.103767,18.108618,16.113468,14.118319,12.123169,12.919667,13.716166,14.508759,15.305257,16.101755,16.69913,17.296501,17.893875,18.49125,19.088623,18.538101,17.991486,17.44487,16.898252,16.351637,15.734741,15.12175,14.504854,13.891863,13.274967,13.2905855,13.310107,13.325725,13.345247,13.360865,12.751778,12.138786,11.525795,10.912805,10.299813,10.58093,10.865952,11.147068,11.428185,11.713207,12.798631,13.884054,14.969479,16.050997,17.136421,18.651329,20.166237,21.681147,23.196054,24.710962,24.343948,23.976934,23.60992,23.242907,22.875893,22.231667,21.591345,20.947119,20.306797,19.662569,20.361458,21.06425,21.763138,22.462027,23.160913,22.914936,22.668959,22.419077,22.1731,21.923218,21.54449,21.165764,20.783133,20.404406,20.025679,19.518106,19.010534,18.502962,17.99539,17.487818,17.893875,18.296028,18.702087,19.108145,19.514202,18.174992,16.835783,15.500477,14.161267,12.825961,12.533132,12.244205,11.955279,11.666354,11.373524,10.471607,9.565785,8.659965,7.7541428,6.8483214,7.387129,7.9259367,8.460839,8.999647,9.538455,10.182681,10.826907,11.471134,12.119265,12.763491,1.1244678,1.1361811,1.1439898,1.1557031,1.1635119,1.175225,1.1908426,1.2064602,1.2181735,1.2337911,1.2494087,1.2923572,1.3353056,1.3782539,1.4212024,1.4641509,1.4407244,1.4212024,1.4016805,1.3821584,1.3626363,1.3821584,1.4016805,1.4212024,1.4407244,1.4641509,1.4485333,1.43682,1.4251068,1.4133936,1.4016805,1.3626363,1.3235924,1.2884527,1.2494087,1.2142692,1.1361811,1.0619974,0.9878138,0.9136301,0.8394465,5.1889505,9.538455,13.887959,18.237463,22.586967,20.146715,17.70256,15.258404,12.818152,10.373997,8.878611,7.3832245,5.891743,4.396357,2.900971,2.4285383,1.9561055,1.4836729,1.0112402,0.5388075,0.5231899,0.5114767,0.4997635,0.48805028,0.47633708,0.44119745,0.40605783,0.3709182,0.3357786,0.30063897,0.25769055,0.21474212,0.1717937,0.12884527,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.30063897,0.57394713,0.8511597,1.1244678,1.4016805,1.9639144,2.5300527,3.096191,3.6584249,4.224563,4.728231,5.2358036,5.7394714,6.2431393,6.7507114,7.5120697,8.273428,9.0386915,9.80005,10.561408,10.049932,9.538455,9.023073,8.511597,8.00012,8.171914,8.339804,8.511597,8.679486,8.85128,8.355421,7.859562,7.363703,6.871748,6.375889,6.4695945,6.5633,6.66091,6.754616,6.8483214,7.2582836,7.6682463,8.078208,8.488171,8.898132,9.577498,10.256865,10.932326,11.611692,12.287154,12.287154,12.287154,12.287154,12.287154,12.287154,11.213444,10.135828,9.062118,7.988407,6.910792,6.7975645,6.6843367,6.5672045,6.453977,6.336845,6.571109,6.801469,7.0357327,7.266093,7.5003567,7.328563,7.1606736,6.98888,6.8209906,6.649197,5.8683167,5.0913405,4.31046,3.5295796,2.7486992,3.049338,3.349977,3.6506162,3.951255,4.251894,4.2557983,4.263607,4.271416,4.279225,4.2870336,4.415879,4.548629,4.677474,4.806319,4.939069,5.368553,5.801942,6.2353306,6.6687193,7.098203,7.3988423,7.6955767,7.9923115,8.289046,8.58578,8.304664,8.023546,7.7385254,7.4574084,7.1762915,7.0044975,6.8366084,6.6648145,6.4969254,6.3251314,6.551587,6.774138,7.000593,7.223144,7.4495993,7.492548,7.535496,7.578445,7.621393,7.6643414,6.785851,5.9073606,5.02887,4.154284,3.2757936,4.6813784,6.0908675,7.4964523,8.905942,10.311526,10.674636,11.037745,11.400854,11.763964,12.123169,12.353529,12.583888,12.814248,13.044608,13.274967,12.423808,11.576552,10.725393,9.874233,9.023073,8.941081,8.855185,8.769287,8.683391,8.601398,9.034787,9.468176,9.905469,10.338858,10.77615,10.686349,10.600452,10.510651,10.424754,10.338858,10.284196,10.2334385,10.178777,10.128019,10.073358,10.491129,10.9089,11.326671,11.744442,12.162213,16.281357,20.400501,24.52355,28.642694,32.76184,32.25817,31.750599,31.246931,30.743263,30.235691,26.038458,21.841227,17.643993,13.446761,9.249529,7.656533,6.0635366,4.4705405,2.8814487,1.2884527,1.1517987,1.0112402,0.8745861,0.737932,0.60127795,0.92534333,1.2494087,1.5734742,1.901444,2.2255092,3.1586614,4.095718,5.02887,5.9659266,6.899079,9.339331,11.775677,14.212025,16.64837,19.088623,19.229181,19.365835,19.506393,19.646952,19.78751,18.104713,16.421915,14.739119,13.056321,11.373524,11.2446785,11.115833,10.983084,10.8542385,10.725393,9.749292,8.769287,7.793187,6.813182,5.8370814,6.5008297,7.1606736,7.824422,8.488171,9.151918,8.706817,8.265619,7.824422,7.37932,6.9381227,6.914696,6.89127,6.871748,6.8483214,6.824895,7.1567693,7.4847393,7.816613,8.144583,8.476458,8.581876,8.691199,8.796618,8.905942,9.01136,8.941081,8.870802,8.804427,8.734148,8.663869,8.351517,8.043069,7.7307167,7.422269,7.113821,8.148487,9.183154,10.217821,11.252487,12.287154,10.202203,8.117252,6.0323014,3.9473507,1.8623998,1.53443,1.2064602,0.8784905,0.5544251,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.12884527,0.25378615,0.38263142,0.5114767,0.63641757,0.7262188,0.8160201,0.9058213,0.9956226,1.0893283,1.4914817,1.8975395,2.3035975,2.7057507,3.1118085,3.049338,2.9868677,2.9243972,2.8619268,2.7994564,2.803361,2.8111696,2.815074,2.8189783,2.8267872,2.5808098,2.3348327,2.0888553,1.8467822,1.6008049,1.6320401,1.6632754,1.698415,1.7296503,1.7608855,1.8311646,1.901444,1.9717231,2.0420024,2.1122816,3.0220075,3.9317331,4.841459,5.7511845,6.66091,6.4891167,6.3173227,6.1455293,5.9737353,5.801942,5.134289,4.466636,3.7989833,3.1313305,2.463678,3.084478,3.7091823,4.3299823,4.950782,5.575486,7.141152,8.706817,10.268578,11.834243,13.399908,13.235924,13.075843,12.911859,12.751778,12.587793,12.724447,12.857197,12.993851,13.1266,13.263254,15.028045,16.792833,18.557625,20.322414,22.087204,20.779228,19.46735,18.159374,16.847496,15.535617,15.754263,15.969006,16.183748,16.398489,16.613232,19.256512,21.903696,24.546976,27.194162,29.837442,33.394352,36.951263,40.508175,44.06899,47.6259,47.90311,48.184227,48.465343,48.746464,49.023674,47.208126,45.388676,43.573128,41.753677,39.93813,34.432922,28.931622,23.430319,17.929016,12.423808,12.408191,12.396477,12.380859,12.365242,12.349625,14.399435,16.449247,18.499058,20.548868,22.59868,23.231194,23.863707,24.49622,25.128733,25.761246,28.81449,31.863827,34.913166,37.9625,41.01184,37.451027,33.886307,30.325493,26.760773,23.199959,22.883701,22.57135,22.255093,21.938837,21.626484,24.746101,27.869623,30.993145,34.11667,37.236286,38.76681,40.297337,41.82786,43.358387,44.888912,41.00794,37.130867,33.253796,29.376722,25.499651,25.487938,25.476225,25.460608,25.448895,25.437181,25.175587,24.917894,24.6563,24.39861,24.137014,24.242434,24.347853,24.453272,24.558691,24.664108,25.827621,26.991133,28.158548,29.322062,30.485573,28.63879,26.792007,24.945227,23.098444,21.251661,21.735807,22.219954,22.7041,23.188246,23.676296,22.770473,21.864653,20.958832,20.056915,19.151093,17.530766,15.914344,14.297921,12.681499,11.061172,12.01775,12.974329,13.927003,14.883581,15.836256,16.351637,16.867018,17.382399,17.89778,18.41316,17.796265,17.183275,16.56638,15.953387,15.336493,15.152986,14.965574,14.782067,14.59856,14.411149,14.30573,14.204215,14.098797,13.993378,13.887959,13.150026,12.412095,11.674163,10.936231,10.198298,10.705871,11.209538,11.713207,12.220779,12.724447,13.591225,14.454097,15.320874,16.183748,17.050524,18.760653,20.470781,22.18091,23.891037,25.601166,25.230247,24.85933,24.48841,24.121397,23.750479,22.91884,22.0833,21.251661,20.420023,19.588387,20.298986,21.013493,21.724094,22.4386,23.1492,23.008642,22.868084,22.73143,22.590872,22.450314,22.106726,21.759233,21.415646,21.068155,20.724567,20.244326,19.764084,19.283842,18.8036,18.32336,18.830933,19.338505,19.846077,20.35365,20.861221,19.248703,17.636185,16.023666,14.411149,12.798631,12.341816,11.881096,11.420377,10.959657,10.498938,9.854712,9.2104845,8.566258,7.918128,7.2739015,7.7111945,8.148487,8.58578,9.023073,9.464272,10.131924,10.795672,11.4633255,12.130978,12.798631,1.1869383,1.1908426,1.1986516,1.2025559,1.2064602,1.2142692,1.2337911,1.2533131,1.2728351,1.2923572,1.3118792,1.3665408,1.4172981,1.4680552,1.5227169,1.5734742,1.5266213,1.4797685,1.4329157,1.3860629,1.33921,1.3743496,1.4055848,1.4407244,1.475864,1.5110037,1.4875772,1.4641509,1.43682,1.4133936,1.3860629,1.33921,1.2884527,1.2376955,1.1869383,1.1361811,1.0502841,0.96438736,0.8745861,0.78868926,0.698888,5.938596,11.174399,16.414106,21.64991,26.885714,22.99693,19.108145,15.215456,11.326671,7.437886,6.477403,5.5169206,4.5564375,3.5959544,2.639376,2.194274,1.7530766,1.3118792,0.8667773,0.42557985,0.42557985,0.42557985,0.42557985,0.42557985,0.42557985,0.40605783,0.39044023,0.3709182,0.3553006,0.3357786,0.28502136,0.23426414,0.1796025,0.12884527,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.1639849,0.31235218,0.46071947,0.61299115,0.76135844,1.3431144,1.9287747,2.5105307,3.0922866,3.6740425,4.154284,4.630621,5.1069584,5.5832953,6.0635366,6.813182,7.562827,8.312472,9.062118,9.811763,9.37447,8.937177,8.499884,8.062591,7.6252975,7.422269,7.2192397,7.016211,6.813182,6.6140575,6.2040954,5.794133,5.3841705,4.9742084,4.564246,5.099149,5.6340523,6.168956,6.703859,7.238762,7.8556576,8.472553,9.089449,9.706344,10.323239,10.983084,11.639023,12.298867,12.954806,13.610746,13.501423,13.388195,13.274967,13.16174,13.048512,11.912332,10.77615,9.636065,8.499884,7.363703,7.2543793,7.1489606,7.039637,6.9342184,6.824895,6.9342184,7.043542,7.1567693,7.266093,7.375416,7.3012323,7.230953,7.1567693,7.08649,7.012306,6.1494336,5.282656,4.415879,3.5530062,2.6862288,3.049338,3.4124475,3.775557,4.138666,4.5017757,4.5095844,4.521298,4.5291066,4.5408196,4.548629,4.6267166,4.704805,4.7828927,4.860981,4.939069,5.3607445,5.7824197,6.2040954,6.6257706,7.0513506,7.3168497,7.5862536,7.8517528,8.121157,8.386656,8.066495,7.7424297,7.4183645,7.098203,6.774138,6.5633,6.356367,6.1455293,5.9346914,5.7238536,6.114294,6.5008297,6.8873653,7.2739015,7.6643414,7.4417906,7.2192397,6.996689,6.774138,6.551587,5.9425,5.3334136,4.728231,4.1191444,3.513962,4.9742084,6.4305506,7.890797,9.351044,10.81129,10.963562,11.111929,11.2642,11.412568,11.560935,11.525795,11.490656,11.45942,11.424281,11.389141,10.71368,10.0382185,9.362757,8.687295,8.011833,8.093826,8.175818,8.261715,8.343708,8.4257,8.941081,9.460366,9.975748,10.495033,11.014318,11.014318,11.014318,11.014318,11.014318,11.014318,10.780055,10.545791,10.315431,10.081166,9.850807,10.377901,10.904996,11.43209,11.959184,12.486279,17.4722,22.458122,27.444044,32.42606,37.411983,35.647194,33.882404,32.117615,30.352823,28.588034,24.144823,19.701614,15.258404,10.819098,6.375889,5.3334136,4.2948427,3.2562714,2.2137961,1.175225,1.1010414,1.0268579,0.94876975,0.8745861,0.80040246,1.1010414,1.4016805,1.698415,1.999054,2.2996929,2.8658314,3.435874,4.0020123,4.5681505,5.138193,7.8868923,10.6355915,13.388195,16.136894,18.885593,19.194042,19.50249,19.810938,20.119385,20.423927,19.13938,17.854832,16.570284,15.285735,14.001186,13.208592,12.419904,11.631214,10.838621,10.049932,8.991838,7.9337454,6.8756523,5.8214636,4.7633705,5.4388323,6.114294,6.785851,7.461313,8.136774,7.8205175,7.5081654,7.191909,6.8756523,6.5633,6.6335793,6.703859,6.774138,6.844417,6.910792,7.238762,7.5667315,7.8947015,8.2226715,8.550641,8.484266,8.421796,8.355421,8.289046,8.226576,8.316377,8.406178,8.495979,8.58578,8.675582,8.331994,7.988407,7.648724,7.3051367,6.9615493,8.16801,9.370565,10.577025,11.783486,12.986042,10.858143,8.726339,6.5984397,4.466636,2.338737,1.9053483,1.4719596,1.038571,0.60908675,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.0,0.0,0.0,0.0,0.0,0.1717937,0.339683,0.5114767,0.679366,0.8511597,0.95657855,1.0659018,1.1713207,1.2806439,1.3860629,1.8038338,2.2177005,2.631567,3.049338,3.4632049,3.338264,3.213323,3.0883822,2.9634414,2.8385005,2.7643168,2.6940374,2.619854,2.5456703,2.475391,2.2645533,2.0537157,1.8467822,1.6359446,1.4251068,1.4094892,1.3938715,1.3782539,1.3665408,1.3509232,1.4992905,1.6437533,1.7921207,1.9404879,2.0888553,2.8814487,3.6740425,4.466636,5.2592297,6.0518236,5.958118,5.8644123,5.7707067,5.6809053,5.5871997,4.860981,4.1308575,3.4046388,2.67842,1.9482968,2.5534792,3.1586614,3.7638438,4.369026,4.9742084,6.6843367,8.39056,10.096785,11.806912,13.513136,12.950902,12.388668,11.826434,11.2642,10.698062,10.990892,11.283723,11.576552,11.869383,12.162213,14.231546,16.300879,18.374117,20.44345,22.512783,20.607435,18.702087,16.796738,14.89139,12.986042,13.544372,14.102701,14.661031,15.21936,15.773785,18.784079,21.794373,24.804668,27.814962,30.825256,34.186947,37.54473,40.90642,44.26421,47.6259,47.579044,47.52829,47.481438,47.43458,47.38773,45.548756,43.70588,41.866905,40.02793,38.188957,32.828213,27.471375,22.114534,16.757694,11.400854,11.666354,11.935758,12.201257,12.470661,12.73616,13.411622,14.087084,14.762545,15.438006,16.113468,16.660084,17.206701,17.753317,18.303837,18.850454,21.013493,23.176533,25.335667,27.498705,29.661743,27.23711,24.812477,22.387842,19.96321,17.538574,18.705992,19.873407,21.040823,22.20824,23.375656,25.843239,28.310822,30.778402,33.245987,35.713566,36.791183,37.868797,38.94641,40.02403,41.101643,37.70481,34.311886,30.915056,27.518227,24.125301,24.086258,24.051117,24.012074,23.97303,23.937891,23.58259,23.22729,22.871988,22.516687,22.161386,22.641628,23.117966,23.594303,24.07064,24.55088,25.26929,25.991606,26.710016,27.428427,28.15074,26.72173,25.288813,23.859802,22.430792,21.00178,21.466404,21.934933,22.40346,22.868084,23.336613,21.911505,20.482494,19.053482,17.628376,16.199366,14.96167,13.72007,12.47847,11.240774,9.999174,11.115833,12.228588,13.345247,14.458001,15.57466,16.008049,16.441439,16.870922,17.30431,17.7377,17.054428,16.371159,15.6917925,15.008522,14.325252,14.571229,14.813302,15.059279,15.305257,15.551234,15.320874,15.0944195,14.867964,14.641508,14.411149,13.548276,12.689307,11.826434,10.963562,10.100689,10.826907,11.553126,12.28325,13.009468,13.735687,14.383818,15.028045,15.672271,16.316498,16.960724,18.866072,20.77142,22.67677,24.582117,26.487465,26.116547,25.741724,25.370806,24.995983,24.625065,23.602112,22.579159,21.556206,20.53325,19.514202,20.236517,20.962736,21.688955,22.411268,23.137487,23.106253,23.071114,23.039877,23.008642,22.973503,22.665054,22.356607,22.044254,21.735807,21.423454,20.970545,20.521538,20.068628,19.615717,19.162806,19.771893,20.38098,20.99397,21.603058,22.212145,20.326319,18.436588,16.55076,14.661031,12.775204,12.146595,11.514082,10.885473,10.256865,9.6243515,9.24172,8.855185,8.468649,8.086017,7.699481,8.039165,8.374943,8.710721,9.050405,9.386183,10.077262,10.768341,11.45942,12.146595,12.837675,1.2494087,1.2494087,1.2494087,1.2494087,1.2494087,1.2494087,1.2767396,1.3001659,1.3235924,1.3509232,1.3743496,1.43682,1.4992905,1.5617609,1.6242313,1.6867018,1.6125181,1.5383345,1.4641509,1.3860629,1.3118792,1.3626363,1.4133936,1.4641509,1.5110037,1.5617609,1.5266213,1.4875772,1.4485333,1.4133936,1.3743496,1.3118792,1.2494087,1.1869383,1.1244678,1.0619974,0.96438736,0.8628729,0.76135844,0.6637484,0.5622339,6.688241,12.814248,18.936352,25.062359,31.188366,25.851048,20.51373,15.176412,9.839094,4.5017757,4.0761957,3.6506162,3.2250361,2.7994564,2.3738766,1.9639144,1.5500476,1.1361811,0.7262188,0.31235218,0.3240654,0.3357786,0.3513962,0.3631094,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.7262188,1.3235924,1.9248703,2.5261483,3.1235218,3.5764325,4.025439,4.474445,4.9234514,5.376362,6.114294,6.8483214,7.5862536,8.324185,9.062118,8.699008,8.335898,7.9766936,7.6135845,7.250475,6.676528,6.098676,5.5247293,4.950782,4.376835,4.0488653,3.7247996,3.4007344,3.076669,2.7486992,3.7247996,4.7009,5.6730967,6.649197,7.6252975,8.449126,9.276859,10.100689,10.924518,11.748346,12.388668,13.025085,13.661504,14.301826,14.938243,14.711788,14.489237,14.262781,14.036326,13.813775,12.611219,11.412568,10.213917,9.01136,7.812709,7.7111945,7.6135845,7.5120697,7.4105554,7.3129454,7.3012323,7.2856145,7.2739015,7.262188,7.250475,7.2739015,7.3012323,7.3246584,7.348085,7.375416,6.426646,5.473972,4.5252023,3.5764325,2.6237583,3.049338,3.474918,3.900498,4.3260775,4.7516575,4.7633705,4.775084,4.786797,4.7985106,4.814128,4.8375545,4.860981,4.8883114,4.911738,4.939069,5.349031,5.7628975,6.1767645,6.5867267,7.000593,7.238762,7.47693,7.7111945,7.9493628,8.187531,7.824422,7.461313,7.098203,6.7389984,6.375889,6.126007,5.8761253,5.6262436,5.376362,5.12648,5.6730967,6.223617,6.774138,7.3246584,7.8751793,7.387129,6.899079,6.4110284,5.9268827,5.4388323,5.099149,4.7633705,4.423688,4.087909,3.7482262,5.263134,6.774138,8.289046,9.80005,11.311053,11.248583,11.186112,11.123642,11.061172,10.998701,10.698062,10.401327,10.100689,9.80005,9.499411,8.999647,8.499884,8.00012,7.5003567,7.000593,7.250475,7.5003567,7.7502384,8.00012,8.250002,8.85128,9.448653,10.049932,10.651209,11.248583,11.338385,11.424281,11.514082,11.599979,11.685876,11.275913,10.862047,10.44818,10.0382185,9.6243515,10.260769,10.901091,11.537509,12.173926,12.814248,18.663042,24.511837,30.364536,36.21333,42.062126,39.036213,36.014206,32.988297,29.962383,26.936472,22.251188,17.562002,12.8767185,8.187531,3.4983444,3.0141985,2.5261483,2.0380979,1.5500476,1.0619974,1.0502841,1.038571,1.0268579,1.0112402,0.999527,1.2767396,1.5500476,1.8233559,2.1005683,2.3738766,2.5769055,2.77603,2.9751544,3.174279,3.3734035,6.4383593,9.499411,12.564366,15.625418,18.68647,19.162806,19.639143,20.111576,20.587914,21.06425,20.174046,19.287746,18.401447,17.511244,16.624945,15.176412,13.723974,12.27544,10.826907,9.37447,8.238289,7.098203,5.9620223,4.825841,3.6857557,4.376835,5.0640097,5.7511845,6.4383593,7.125534,6.9381227,6.7507114,6.5633,6.375889,6.1884775,6.348558,6.5125427,6.676528,6.8366084,7.000593,7.3246584,7.648724,7.9766936,8.300759,8.624825,8.386656,8.148487,7.914223,7.676055,7.437886,7.687768,7.9376497,8.187531,8.437413,8.687295,8.312472,7.9376497,7.562827,7.1880045,6.813182,8.187531,9.561881,10.936231,12.31058,13.688834,11.514082,9.339331,7.1606736,4.985922,2.8111696,2.2762666,1.737459,1.1986516,0.6637484,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.21083772,0.42557985,0.63641757,0.8511597,1.0619974,1.1869383,1.3118792,1.43682,1.5617609,1.6867018,2.1122816,2.5378613,2.9634414,3.3890212,3.8106966,3.6232853,3.435874,3.2484627,3.0610514,2.87364,2.7252727,2.5769055,2.4246337,2.2762666,2.1239948,1.9482968,1.7765031,1.6008049,1.4251068,1.2494087,1.1869383,1.1244678,1.0619974,0.999527,0.93705654,1.1635119,1.3860629,1.6125181,1.8389735,2.0615244,2.736986,3.4124475,4.087909,4.7633705,5.4388323,5.423215,5.4115014,5.3997884,5.388075,5.376362,4.5876727,3.7989833,3.0141985,2.2255092,1.43682,2.0263848,2.612045,3.2016098,3.78727,4.376835,6.223617,8.074304,9.924991,11.775677,13.626364,12.661977,11.701493,10.737106,9.776623,8.812236,9.261242,9.714153,10.163159,10.612165,11.061172,13.438952,15.812829,18.186707,20.564487,22.938364,20.435642,17.936825,15.438006,12.939189,10.436467,11.338385,12.236397,13.138313,14.036326,14.938243,18.311647,21.688955,25.062359,28.435762,31.81307,34.975636,38.138203,41.300766,44.463333,47.6259,47.251076,46.876255,46.50143,46.12661,45.751785,43.885483,42.026985,40.160683,38.298283,36.435883,31.223505,26.011127,20.79875,15.586374,10.373997,10.924518,11.475039,12.025558,12.576079,13.1266,12.423808,11.72492,11.0260315,10.323239,9.6243515,10.088976,10.549695,11.014318,11.475039,11.935758,13.212498,14.489237,15.762072,17.03881,18.311647,17.023193,15.738646,14.450192,13.16174,11.873287,14.524376,17.175465,19.826555,22.47374,25.124828,26.936472,28.748114,30.563662,32.375305,34.186947,34.81165,35.436356,36.061058,36.685764,37.314373,34.401688,31.489004,28.57632,25.663635,22.750952,22.688482,22.62601,22.563541,22.50107,22.4386,21.98569,21.536682,21.087677,20.63867,20.18576,21.036919,21.888079,22.739239,23.586494,24.437654,24.710962,24.988174,25.261482,25.538694,25.812004,24.800762,23.785618,22.774378,21.763138,20.751898,21.200905,21.64991,22.098917,22.551826,23.000834,21.048632,19.100336,17.148134,15.199838,13.251541,12.388668,11.525795,10.662923,9.80005,8.937177,10.213917,11.486752,12.763491,14.036326,15.313066,15.664462,16.011953,16.36335,16.710842,17.062239,16.312593,15.562947,14.813302,14.063657,13.314012,13.989473,14.661031,15.336493,16.011953,16.687416,16.33602,15.988527,15.637131,15.285735,14.938243,13.950429,12.962616,11.974802,10.986988,9.999174,10.951848,11.900618,12.849388,13.798158,14.750832,15.176412,15.598087,16.023666,16.449247,16.874826,18.975395,21.075964,23.176533,25.273195,27.373764,26.998941,26.624119,26.249296,25.874474,25.499651,24.289286,23.075018,21.860748,20.650383,19.436115,20.174046,20.911978,21.64991,22.387842,23.125774,23.199959,23.274141,23.348326,23.426414,23.500597,23.223385,22.950077,22.67677,22.399555,22.126247,21.700668,21.275087,20.849508,20.423927,19.998348,20.712854,21.423454,22.13796,22.848562,23.563068,21.400028,19.23699,17.073952,14.9109125,12.751778,11.951375,11.150972,10.350571,9.550168,8.749765,8.624825,8.499884,8.374943,8.250002,8.125061,8.36323,8.601398,8.835662,9.073831,9.311999,10.0265045,10.737106,11.4516115,12.162213,12.8767185,1.261122,1.2728351,1.2806439,1.2923572,1.3040704,1.3118792,1.3274968,1.3431144,1.358732,1.3743496,1.3860629,1.4407244,1.4914817,1.5461433,1.5969005,1.6515622,1.5812829,1.5149081,1.4485333,1.3782539,1.3118792,1.3509232,1.3938715,1.4329157,1.4719596,1.5110037,1.4680552,1.4212024,1.3782539,1.3314011,1.2884527,1.2415999,1.1908426,1.1439898,1.097137,1.0502841,0.98390937,0.92143893,0.8550641,0.78868926,0.7262188,6.1221027,11.517986,16.917774,22.31366,27.713448,23.028164,18.346786,13.665408,8.98403,4.298747,3.9317331,3.5608149,3.1898966,2.8189783,2.4480603,2.05762,1.6632754,1.2728351,0.8784905,0.48805028,0.46071947,0.43338865,0.40605783,0.37872702,0.3513962,0.3435874,0.339683,0.3357786,0.3318742,0.3240654,0.26940376,0.21474212,0.16008049,0.10541886,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.62470436,1.1517987,1.6749885,2.1981785,2.7252727,3.1430438,3.5647192,3.9863946,4.4041657,4.825841,5.575486,6.3251314,7.0747766,7.824422,8.574067,8.242193,7.910319,7.578445,7.2465706,6.910792,6.426646,5.938596,5.4505453,4.9624953,4.474445,4.169902,3.8653584,3.5608149,3.2562714,2.951728,3.8614538,4.7711797,5.6809053,6.590631,7.5003567,8.460839,9.421323,10.381805,11.338385,12.298867,12.70102,13.09927,13.501423,13.899672,14.301826,13.989473,13.6810255,13.368673,13.0602255,12.751778,11.721016,10.694158,9.6673,8.640442,7.6135845,7.453504,7.297328,7.141152,6.9810715,6.824895,6.89127,6.9615493,7.027924,7.094299,7.1606736,7.1567693,7.152865,7.1489606,7.141152,7.137247,6.356367,5.579391,4.7985106,4.01763,3.2367494,3.533484,3.8263142,4.123049,4.415879,4.7126136,4.716518,4.7243266,4.728231,4.732136,4.73604,4.7907014,4.841459,4.8961205,4.9468775,5.001539,5.349031,5.700427,6.0518236,6.3993154,6.7507114,6.918601,7.0903945,7.2582836,7.4300776,7.601871,7.328563,7.055255,6.7819467,6.5086384,6.239235,5.9073606,5.579391,5.2475166,4.9156423,4.5876727,5.087436,5.5871997,6.086963,6.5867267,7.08649,6.860035,6.6335793,6.4032197,6.1767645,5.950309,5.493494,5.036679,4.575959,4.1191444,3.6623292,5.4036927,7.141152,8.882515,10.6238785,12.361338,11.943566,11.521891,11.10412,10.682445,10.260769,10.053836,9.8429985,9.63216,9.421323,9.21439,8.847376,8.484266,8.117252,7.7541428,7.387129,7.5940623,7.7970915,8.0040245,8.207053,8.413987,9.112875,9.811763,10.510651,11.213444,11.912332,12.072412,12.232492,12.392572,12.552653,12.712734,12.517513,12.322293,12.127073,11.931853,11.736633,12.373051,13.013372,13.64979,14.286208,14.92653,20.67381,26.42109,32.16837,37.91565,43.66293,40.09821,36.537395,32.97658,29.411861,25.851048,21.341463,16.835783,12.326198,7.8205175,3.310933,3.0141985,2.717464,2.4207294,2.1239948,1.8233559,1.9053483,1.9834363,2.0654287,2.1435168,2.2255092,2.3348327,2.4441557,2.5534792,2.6667068,2.77603,3.252367,3.7287042,4.2089458,4.6852827,5.1616197,7.7775693,10.393518,13.009468,15.621513,18.237463,18.45611,18.678661,18.897306,19.115953,19.338505,19.197947,19.057388,18.916828,18.77627,18.635712,17.17937,15.719124,14.258877,12.798631,11.338385,10.159255,8.98403,7.8049,6.6257706,5.4505453,6.153338,6.860035,7.5667315,8.269524,8.976221,8.640442,8.304664,7.968885,7.633106,7.3012323,7.2934237,7.2856145,7.277806,7.269997,7.262188,7.5433054,7.8283267,8.109444,8.39056,8.675582,8.831758,8.991838,9.148014,9.304191,9.464272,9.600925,9.741484,9.882042,10.0226,10.163159,9.503315,8.847376,8.191436,7.531592,6.8756523,7.699481,8.52331,9.351044,10.174872,10.998701,9.4018,7.8049,6.2079997,4.6110992,3.0141985,2.4831998,1.9522011,1.4212024,0.8941081,0.3631094,0.28892577,0.21864653,0.14446288,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.19131571,0.38653582,0.57785153,0.76916724,0.96438736,1.1908426,1.4172981,1.6437533,1.8741131,2.1005683,2.4441557,2.7838387,3.1274261,3.4710135,3.8106966,3.5998588,3.3890212,3.174279,2.9634414,2.7486992,2.6549935,2.5612879,2.463678,2.3699722,2.2762666,2.0380979,1.7999294,1.5617609,1.3235924,1.0893283,1.0893283,1.0932326,1.0932326,1.097137,1.1010414,1.2923572,1.4836729,1.678893,1.8702087,2.0615244,2.6471848,3.232845,3.8185053,4.4041657,4.985922,4.860981,4.73604,4.6110992,4.4861584,4.3612175,3.7208953,3.0805733,2.4441557,1.8038338,1.1635119,1.6710842,2.1786566,2.6862288,3.193801,3.7013733,5.298274,6.899079,8.499884,10.100689,11.701493,11.2642,10.8308115,10.393518,9.96013,9.526741,10.081166,10.6355915,11.190017,11.744442,12.298867,14.016804,15.734741,17.452679,19.170614,20.888552,18.549814,16.211079,13.8762455,11.537509,9.198771,10.163159,11.131451,12.095839,13.0602255,14.024612,17.714273,21.403933,25.093594,28.783253,32.476818,35.291893,38.11087,40.925945,43.744923,46.5639,46.665417,46.76693,46.868446,46.97386,47.07538,44.322773,41.57017,38.817566,36.064964,33.31236,28.630981,23.9457,19.26432,14.582942,9.901564,10.541886,11.178304,11.818625,12.458947,13.09927,12.076316,11.0494585,10.0265045,8.999647,7.9766936,8.343708,8.710721,9.077735,9.444749,9.811763,11.701493,13.591225,15.480955,17.370686,19.26432,18.74113,18.217941,17.694752,17.17156,16.64837,17.686943,18.72161,19.756275,20.790941,21.82561,23.301472,24.773432,26.249296,27.72516,29.201025,30.141985,31.086851,32.027813,32.968773,33.91364,31.926298,29.938957,27.951616,25.964275,23.976934,23.348326,22.719717,22.091108,21.466404,20.837795,20.38098,19.92807,19.471254,19.018343,18.56153,19.604004,20.646479,21.688955,22.73143,23.773905,24.527454,25.281004,26.03065,26.784199,27.537748,26.143877,24.75391,23.360039,21.966167,20.5762,21.009588,21.446882,21.88027,22.31366,22.750952,21.122816,19.49468,17.866545,16.238409,14.614178,13.466284,12.322293,11.178304,10.034314,8.886419,10.09288,11.29934,12.501896,13.708356,14.9109125,15.391153,15.867491,16.343828,16.82407,17.300406,16.476578,15.656653,14.832824,14.008995,13.189071,13.759113,14.33306,14.903104,15.477051,16.050997,15.836256,15.625418,15.410676,15.199838,14.989,14.133936,13.282777,12.431617,11.576552,10.725393,11.471134,12.216875,12.958711,13.704452,14.450192,14.879677,15.309161,15.738646,16.168129,16.601519,18.436588,20.271656,22.106726,23.941795,25.776863,25.644114,25.515268,25.386423,25.253674,25.124828,23.891037,22.653341,21.41955,20.18576,18.948065,19.701614,20.455164,21.208714,21.958359,22.711908,22.82904,22.946173,23.063305,23.184341,23.301472,22.977407,22.653341,22.333181,22.009115,21.688955,21.091581,20.498112,19.900738,19.30727,18.7138,19.506393,20.30289,21.09939,21.891983,22.688482,20.693333,18.698183,16.703033,14.707883,12.712734,12.025558,11.338385,10.651209,9.964035,9.276859,9.089449,8.905942,8.718531,8.535024,8.351517,8.52331,8.695104,8.866898,9.0386915,9.21439,9.874233,10.534078,11.193921,11.8537655,12.513609,1.2767396,1.2962615,1.3157835,1.3353056,1.3548276,1.3743496,1.3782539,1.3860629,1.3899672,1.3938715,1.4016805,1.4407244,1.4836729,1.5266213,1.5695697,1.6125181,1.5539521,1.4914817,1.4329157,1.3743496,1.3118792,1.3431144,1.3743496,1.4016805,1.4329157,1.4641509,1.4094892,1.358732,1.3040704,1.2533131,1.1986516,1.1674163,1.1361811,1.1010414,1.0698062,1.038571,1.0073358,0.97610056,0.94876975,0.91753453,0.8862993,5.5559645,10.22563,14.899199,19.568865,24.23853,20.209187,16.183748,12.154405,8.128965,4.0996222,3.7833657,3.4710135,3.154757,2.8385005,2.5261483,2.1513257,1.7804074,1.4055848,1.0346665,0.6637484,0.59346914,0.5270943,0.46071947,0.39434463,0.3240654,0.31625658,0.30454338,0.29673457,0.28502136,0.27330816,0.22645533,0.1796025,0.13274968,0.08589685,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.5231899,0.97610056,1.4251068,1.8741131,2.3231194,2.7135596,3.1039999,3.49444,3.8848803,4.2753205,5.036679,5.7980375,6.5633,7.3246584,8.086017,7.785378,7.480835,7.180196,6.8756523,6.575013,6.1767645,5.774611,5.376362,4.9742084,4.575959,4.290938,4.0059166,3.7208953,3.435874,3.1508527,3.9942036,4.841459,5.6848097,6.5281606,7.375416,8.468649,9.565785,10.6590185,11.756155,12.849388,13.013372,13.173453,13.337439,13.501423,13.661504,13.2671585,12.872814,12.47847,12.084125,11.685876,10.8308115,9.975748,9.120684,8.265619,7.4105554,7.195813,6.9810715,6.7663293,6.551587,6.336845,6.4852123,6.6335793,6.7819467,6.9264097,7.0747766,7.039637,7.0044975,6.969358,6.9342184,6.899079,6.289992,5.6809053,5.0718184,4.4588275,3.8497405,4.0137253,4.181615,4.3455997,4.5095844,4.6735697,4.6735697,4.6696653,4.6657605,4.6657605,4.661856,4.743849,4.8219366,4.903929,4.9820175,5.0640097,5.349031,5.6379566,5.9268827,6.211904,6.5008297,6.602344,6.703859,6.8092775,6.910792,7.012306,6.8287997,6.649197,6.46569,6.282183,6.098676,5.688714,5.278752,4.8687897,4.4588275,4.0488653,4.5017757,4.950782,5.3997884,5.8487945,6.3017054,6.3329406,6.364176,6.3993154,6.4305506,6.461786,5.883934,5.3060827,4.728231,4.154284,3.5764325,5.5442514,7.5081654,9.475985,11.443803,13.411622,12.634645,11.85767,11.080693,10.303718,9.526741,9.405705,9.284669,9.163632,9.0465,8.925464,8.695104,8.464745,8.234385,8.0040245,7.773665,7.9337454,8.093826,8.253906,8.413987,8.574067,9.37447,10.174872,10.975275,11.775677,12.576079,12.806439,13.040704,13.271063,13.505327,13.735687,13.759113,13.78254,13.805966,13.829392,13.848915,14.489237,15.125654,15.762072,16.398489,17.03881,22.680674,28.326439,33.972202,39.61797,45.263737,41.164112,37.06449,32.960964,28.861341,24.761719,20.435642,16.109564,11.779582,7.453504,3.1235218,3.018103,2.9087796,2.803361,2.6940374,2.5886188,2.7604125,2.9322062,3.1039999,3.2757936,3.4514916,3.39683,3.338264,3.2836022,3.2289407,3.174279,3.9317331,4.6852827,5.4388323,6.196286,6.949836,9.116779,11.283723,13.450665,15.621513,17.788456,17.753317,17.718178,17.683039,17.647898,17.612759,18.221846,18.827028,19.436115,20.041296,20.650383,19.178425,17.71037,16.238409,14.770353,13.298394,12.084125,10.865952,9.647778,8.429605,7.211431,7.9337454,8.65606,9.378374,10.100689,10.826907,10.342762,9.858616,9.378374,8.894228,8.413987,8.234385,8.058686,7.8790836,7.703386,7.523783,7.7658563,8.0040245,8.246098,8.484266,8.726339,9.276859,9.8312845,10.381805,10.936231,11.486752,11.517986,11.549222,11.576552,11.607788,11.639023,10.698062,9.757101,8.81614,7.8790836,6.9381227,7.211431,7.4886436,7.7619514,8.039165,8.312472,7.2934237,6.2743745,5.251421,4.2323723,3.213323,2.690133,2.1669433,1.6437533,1.1205635,0.60127795,0.48024148,0.359205,0.23816854,0.12103647,0.0,0.0,0.0,0.0,0.0,0.0,0.1717937,0.3435874,0.5192855,0.6910792,0.8628729,1.1908426,1.5227169,1.8506867,2.182561,2.514435,2.7721257,3.0337205,3.2914112,3.5530062,3.8106966,3.5764325,3.338264,3.1000953,2.8619268,2.6237583,2.5847144,2.5456703,2.5066261,2.463678,2.4246337,2.1239948,1.8233559,1.5266213,1.2259823,0.92534333,0.9917182,1.0580931,1.1283722,1.1947471,1.261122,1.4212024,1.5812829,1.7413634,1.901444,2.0615244,2.5573835,3.0532427,3.5491016,4.041056,4.5369153,4.298747,4.0605783,3.8263142,3.5881457,3.349977,2.8580225,2.366068,1.8741131,1.3782539,0.8862993,1.3157835,1.7413634,2.1708477,2.5964274,3.0259118,4.376835,5.7238536,7.0747766,8.4257,9.776623,9.866425,9.96013,10.053836,10.143637,10.237343,10.897186,11.557031,12.216875,12.8767185,13.536563,14.59856,15.656653,16.71865,17.776743,18.838741,16.663988,14.489237,12.31058,10.135828,7.9610763,8.991838,10.0226,11.053363,12.084125,13.110983,17.1169,21.122816,25.128733,29.130745,33.13666,35.612053,38.083538,40.555027,43.026512,45.501904,46.079754,46.66151,47.239365,47.821117,48.39897,44.756165,41.113358,37.470547,33.831646,30.188839,26.034554,21.884174,17.72989,13.575606,9.425227,10.155351,10.885473,11.615597,12.34572,13.075843,11.72492,10.373997,9.023073,7.676055,6.3251314,6.5984397,6.871748,7.141152,7.4144597,7.687768,10.194394,12.697116,15.203742,17.706465,20.21309,20.455164,20.697237,20.93931,21.181383,21.423454,20.845604,20.263847,19.685997,19.10424,18.526388,19.662569,20.79875,21.938837,23.075018,24.211199,25.47232,26.733442,27.99066,29.251781,30.512903,29.450907,28.388908,27.326912,26.26101,25.199013,24.00817,22.813423,21.62258,20.431738,19.23699,18.77627,18.315552,17.858736,17.398016,16.937298,18.171087,19.408783,20.642574,21.876366,23.114061,24.343948,25.573835,26.803722,28.033607,29.263494,27.490896,25.718298,23.9457,22.1731,20.400501,20.818274,21.239948,21.661623,22.079395,22.50107,21.193096,19.889025,18.584955,17.280884,15.976814,14.547803,13.118792,11.693685,10.264673,8.835662,9.971844,11.108025,12.244205,13.376482,14.512663,15.117846,15.723028,16.32821,16.933393,17.538574,16.640562,15.746454,14.852346,13.958238,13.06413,13.532659,14.001186,14.473619,14.942147,15.410676,15.336493,15.262308,15.188125,15.113941,15.035853,14.321347,13.602938,12.884527,12.166118,11.4516115,11.990419,12.529227,13.0719385,13.610746,14.149553,14.586847,15.020235,15.453624,15.890917,16.324306,17.893875,19.463446,21.036919,22.60649,24.17606,24.289286,24.406418,24.519646,24.636778,24.750006,23.492788,22.23557,20.978354,19.721136,18.463919,19.229181,19.998348,20.76361,21.532778,22.301945,22.458122,22.618202,22.778282,22.938364,23.098444,22.73143,22.360512,21.989594,21.618675,21.251661,20.486399,19.721136,18.955873,18.19061,17.425346,18.303837,19.178425,20.056915,20.935406,21.813896,19.986635,18.15547,16.32821,14.50095,12.67369,12.099743,11.525795,10.951848,10.373997,9.80005,9.554072,9.308095,9.066022,8.8200445,8.574067,8.683391,8.78881,8.898132,9.0035515,9.112875,9.721962,10.327144,10.936231,11.541413,12.150499,1.2884527,1.3157835,1.3470187,1.3782539,1.4055848,1.43682,1.4329157,1.4290112,1.4212024,1.4172981,1.4133936,1.4446288,1.475864,1.5110037,1.542239,1.5734742,1.5227169,1.4680552,1.4172981,1.3665408,1.3118792,1.3314011,1.3509232,1.3743496,1.3938715,1.4133936,1.3509232,1.2923572,1.2337911,1.1713207,1.1127546,1.0932326,1.077615,1.0580931,1.0424755,1.0268579,1.0307622,1.0346665,1.038571,1.0463798,1.0502841,4.9937305,8.933272,12.8767185,16.820166,20.76361,17.390207,14.016804,10.6434,7.2739015,3.900498,3.638903,3.3812122,3.1196175,2.8619268,2.6003318,2.2489357,1.893635,1.542239,1.1908426,0.8394465,0.7301232,0.62079996,0.5153811,0.40605783,0.30063897,0.28502136,0.26940376,0.25378615,0.23816854,0.22645533,0.1835069,0.14446288,0.10541886,0.06637484,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.42557985,0.80040246,1.175225,1.5500476,1.9248703,2.2840753,2.6432803,3.0063896,3.3655949,3.7247996,4.5017757,5.2748475,6.0518236,6.824895,7.601871,7.328563,7.055255,6.7819467,6.5086384,6.239235,5.9268827,5.610626,5.298274,4.985922,4.6735697,4.40807,4.1464753,3.8809757,3.6154766,3.349977,4.1308575,4.911738,5.688714,6.4695945,7.250475,8.480362,9.710248,10.940135,12.170022,13.399908,13.325725,13.251541,13.173453,13.09927,13.025085,12.544845,12.064603,11.584361,11.10412,10.6238785,9.940608,9.261242,8.577971,7.8947015,7.211431,6.9381227,6.6687193,6.395411,6.1221027,5.8487945,6.0791545,6.3056097,6.532065,6.75852,6.98888,6.9225054,6.8561306,6.79366,6.727285,6.66091,6.223617,5.7824197,5.3412223,4.903929,4.462732,4.4978714,4.533011,4.5681505,4.60329,4.6384296,4.6267166,4.618908,4.607195,4.5993857,4.5876727,4.6930914,4.802415,4.911738,5.017157,5.12648,5.349031,5.575486,5.801942,6.0244927,6.250948,6.2860875,6.321227,6.356367,6.3915067,6.426646,6.3329406,6.239235,6.1494336,6.055728,5.9620223,5.473972,4.9820175,4.493967,4.0020123,3.513962,3.912211,4.3143644,4.7126136,5.1108627,5.5130157,5.805846,6.098676,6.3915067,6.6843367,6.9732623,6.278279,5.579391,4.884407,4.185519,3.4866312,5.6809053,7.8790836,10.073358,12.267632,14.461906,13.325725,12.193448,11.057267,9.921086,8.78881,8.757574,8.726339,8.699008,8.667773,8.636538,8.542832,8.449126,8.351517,8.257811,8.164105,8.277332,8.39056,8.507692,8.62092,8.738052,9.636065,10.537982,11.435994,12.337912,13.235924,13.544372,13.848915,14.153459,14.458001,14.762545,15.000713,15.242786,15.480955,15.723028,15.961197,16.601519,17.237936,17.874353,18.51077,19.151093,24.69144,30.235691,35.77604,41.32029,46.860638,42.22611,37.58768,32.94925,28.310822,23.676296,19.525915,15.37944,11.232965,7.08649,2.9361105,3.018103,3.1039999,3.1859922,3.2679846,3.349977,3.6154766,3.8809757,4.1464753,4.40807,4.6735697,4.454923,4.2362766,4.0137253,3.795079,3.5764325,4.607195,5.6418614,6.6726236,7.703386,8.738052,10.455989,12.177831,13.895767,15.617609,17.33945,17.04662,16.757694,16.46877,16.175938,15.8870125,17.24184,18.596668,19.951496,21.306324,22.66115,21.181383,19.701614,18.221846,16.742077,15.262308,14.005091,12.747873,11.490656,10.2334385,8.976221,9.714153,10.455989,11.193921,11.935758,12.67369,12.045081,11.416472,10.783959,10.155351,9.526741,9.17925,8.831758,8.484266,8.136774,7.7892823,7.984503,8.183627,8.378847,8.577971,8.773191,9.721962,10.670732,11.615597,12.564366,13.513136,13.431144,13.353056,13.271063,13.192975,13.110983,11.888905,10.666827,9.444749,8.2226715,7.000593,6.7233806,6.4500723,6.1767645,5.899552,5.6262436,5.181142,4.7399445,4.298747,3.853645,3.4124475,2.8970666,2.3816853,1.8663043,1.3509232,0.8394465,0.6715572,0.5036679,0.3357786,0.1678893,0.0,0.0,0.0,0.0,0.0,0.0,0.15227169,0.30454338,0.45681506,0.60908675,0.76135844,1.1947471,1.6281357,2.0615244,2.4910088,2.9243972,3.1039999,3.279698,3.4593005,3.6349986,3.8106966,3.5491016,3.2875066,3.0259118,2.7643168,2.4988174,2.514435,2.5300527,2.5456703,2.5612879,2.5769055,2.2137961,1.8506867,1.4875772,1.1244678,0.76135844,0.8941081,1.0268579,1.1596074,1.2923572,1.4251068,1.5539521,1.678893,1.8077383,1.9365835,2.0615244,2.4675822,2.87364,3.2757936,3.6818514,4.087909,3.736513,3.3890212,3.0376248,2.6862288,2.338737,1.9912452,1.6476578,1.3040704,0.95657855,0.61299115,0.96048295,1.3079748,1.6554666,2.0029583,2.35045,3.4514916,4.548629,5.64967,6.7507114,7.8517528,8.468649,9.089449,9.710248,10.331048,10.951848,11.713207,12.47847,13.243732,14.008995,14.774258,15.176412,15.578565,15.980719,16.386776,16.788929,14.774258,12.763491,10.748819,8.738052,6.7233806,7.8205175,8.913751,10.010887,11.10412,12.201257,16.519526,20.8417,25.159967,29.478237,33.80041,35.92831,38.05621,40.18411,42.3081,44.436,45.494095,46.55219,47.610283,48.668373,49.726467,45.193455,40.660446,36.127434,31.594423,27.061413,23.438128,19.818747,16.195461,12.572175,8.94889,9.768814,10.588739,11.408664,12.228588,13.048512,11.373524,9.698535,8.023546,6.348558,4.6735697,4.853172,5.02887,5.2084727,5.3841705,5.563773,8.683391,11.803008,14.922626,18.042242,21.16186,22.169195,23.176533,24.183868,25.191204,26.19854,24.004265,21.809992,19.615717,17.421442,15.223265,16.023666,16.82407,17.624472,18.424873,19.225277,20.802654,22.380033,23.957413,25.53479,27.11217,26.975515,26.838861,26.698303,26.56165,26.424995,24.668013,22.911032,21.15405,19.393166,17.636185,17.17156,16.706938,16.242313,15.77769,15.313066,16.738173,18.167183,19.596195,21.021301,22.450314,24.156536,25.866665,27.57289,29.279112,30.98924,28.834011,26.682686,24.531359,22.37613,20.224804,20.630861,21.036919,21.439074,21.84513,22.251188,21.267279,20.28337,19.303364,18.319456,17.335546,15.629322,13.919194,12.209065,10.498938,8.78881,9.850807,10.916709,11.982611,13.048512,14.114414,14.844538,15.578565,16.30869,17.042715,17.776743,16.808453,15.84016,14.871868,13.903577,12.939189,13.306203,13.673217,14.040231,14.407245,14.774258,14.836729,14.899199,14.96167,15.024139,15.086611,14.504854,13.923099,13.341343,12.755682,12.173926,12.509705,12.845484,13.181262,13.513136,13.848915,14.2901125,14.73131,15.168603,15.6098,16.050997,17.355068,18.659138,19.96321,21.271183,22.575254,22.93446,23.293663,23.656773,24.015978,24.375183,23.09454,21.813896,20.53325,19.256512,17.975868,18.756748,19.541533,20.322414,21.103294,21.888079,22.091108,22.294136,22.493261,22.696291,22.899319,22.481548,22.063778,21.646006,21.228235,20.81437,19.877312,18.94416,18.007103,17.073952,16.136894,17.097378,18.057861,19.018343,19.978827,20.93931,19.276033,17.616663,15.957292,14.297921,12.63855,12.173926,11.713207,11.248583,10.787864,10.323239,10.018696,9.714153,9.40961,9.105066,8.800523,8.843472,8.886419,8.929368,8.968412,9.01136,9.565785,10.124115,10.67854,11.232965,11.787391,1.3001659,1.33921,1.3782539,1.4212024,1.4602464,1.4992905,1.4836729,1.4680552,1.456342,1.4407244,1.4251068,1.4485333,1.4680552,1.4914817,1.5149081,1.5383345,1.4914817,1.4485333,1.4016805,1.358732,1.3118792,1.3235924,1.3314011,1.3431144,1.3509232,1.3626363,1.2962615,1.2259823,1.1596074,1.0932326,1.0268579,1.0229534,1.0190489,1.0190489,1.0151446,1.0112402,1.0541886,1.0932326,1.1322767,1.1713207,1.2142692,4.4275923,7.6409154,10.858143,14.0714655,17.288692,14.571229,11.8537655,9.136301,6.4188375,3.7013733,3.49444,3.2914112,3.084478,2.8814487,2.6745155,2.3426414,2.0107672,1.678893,1.3431144,1.0112402,0.8667773,0.71841,0.5700427,0.42167544,0.27330816,0.25378615,0.23426414,0.21474212,0.19522011,0.1756981,0.14055848,0.10932326,0.078088045,0.046852827,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.3240654,0.62470436,0.92534333,1.2259823,1.5266213,1.8545911,2.1864653,2.514435,2.8463092,3.174279,3.9629683,4.7516575,5.5364423,6.3251314,7.113821,6.871748,6.6257706,6.3836975,6.141625,5.899552,5.6730967,5.4505453,5.22409,5.001539,4.775084,4.5291066,4.283129,4.041056,3.795079,3.5491016,4.263607,4.9781127,5.6965227,6.4110284,7.125534,8.488171,9.854712,11.221252,12.583888,13.950429,13.638077,13.325725,13.013372,12.70102,12.388668,11.82253,11.256392,10.694158,10.128019,9.561881,9.054309,8.542832,8.031356,7.523783,7.012306,6.6843367,6.3524623,6.0205884,5.6926184,5.3607445,5.6691923,5.9776397,6.2860875,6.590631,6.899079,6.805373,6.7116675,6.6140575,6.520352,6.426646,6.153338,5.883934,5.6145306,5.3451266,5.0757227,4.9781127,4.884407,4.7907014,4.6930914,4.5993857,4.5837684,4.564246,4.548629,4.5291066,4.513489,4.646239,4.7828927,4.9156423,5.0522966,5.1889505,5.349031,5.5130157,5.6730967,5.8370814,6.001066,5.9659266,5.9346914,5.903456,5.8683167,5.8370814,5.833177,5.833177,5.8292727,5.8292727,5.825368,5.2553253,4.6852827,4.11524,3.5451972,2.9751544,3.3265507,3.6740425,4.025439,4.376835,4.7243266,5.278752,5.8292727,6.3836975,6.9342184,7.4886436,6.6687193,5.852699,5.036679,4.2167544,3.4007344,5.8214636,8.246098,10.666827,13.091461,15.51219,14.020708,12.529227,11.033841,9.542359,8.050878,8.109444,8.171914,8.23048,8.289046,8.351517,8.39056,8.429605,8.468649,8.511597,8.550641,8.62092,8.691199,8.761478,8.831758,8.898132,9.901564,10.901091,11.900618,12.900145,13.899672,14.278399,14.653222,15.031949,15.410676,15.789403,16.246218,16.703033,17.159847,17.616663,18.073479,18.7138,19.350218,19.986635,20.626957,21.263374,26.702208,32.14104,37.583775,43.02261,48.46144,43.28811,38.11087,32.93754,27.764204,22.586967,18.620094,14.653222,10.686349,6.715572,2.7486992,3.0220075,3.2953155,3.5686235,3.8419318,4.1113358,4.4705405,4.825841,5.185046,5.5442514,5.899552,5.5169206,5.1303844,4.743849,4.3612175,3.9746814,5.2865605,6.5945354,7.9064145,9.21439,10.526268,11.799104,13.068034,14.34087,15.613705,16.88654,16.343828,15.797212,15.250595,14.707883,14.161267,16.26574,18.366308,20.470781,22.57135,24.675823,23.184341,21.696764,20.205282,18.7138,17.226223,15.926057,14.629795,13.333533,12.033368,10.737106,11.49456,12.252014,13.009468,13.766922,14.524376,13.7474,12.970425,12.193448,11.416472,10.6355915,10.120211,9.600925,9.085544,8.566258,8.050878,8.203149,8.359325,8.515501,8.671678,8.823949,10.167064,11.510178,12.853292,14.196406,15.535617,15.348206,15.15689,14.965574,14.778163,14.586847,13.083652,11.576552,10.073358,8.566258,7.0630636,6.239235,5.4115014,4.5876727,3.7638438,2.9361105,3.0727646,3.2094188,3.3421683,3.4788225,3.611572,3.1039999,2.5964274,2.0888553,1.5812829,1.0737107,0.8589685,0.6442264,0.42948425,0.21474212,0.0,0.0,0.0,0.0,0.0,0.0,0.13274968,0.26549935,0.39824903,0.5309987,0.6637484,1.1986516,1.7335546,2.2684577,2.803361,3.338264,3.4319696,3.5256753,3.6232853,3.716991,3.8106966,3.5256753,3.2367494,2.951728,2.6628022,2.3738766,2.4441557,2.514435,2.5847144,2.6549935,2.7252727,2.2996929,1.8741131,1.4485333,1.0268579,0.60127795,0.79649806,0.9956226,1.1908426,1.3899672,1.5890918,1.6827974,1.7765031,1.8741131,1.9678187,2.0615244,2.377781,2.6940374,3.0063896,3.3226464,3.638903,3.174279,2.7135596,2.2489357,1.7882162,1.3235924,1.1283722,0.92924774,0.7340276,0.5349031,0.3357786,0.60518235,0.8706817,1.1400855,1.4055848,1.6749885,2.5261483,3.3734035,4.224563,5.0757227,5.9268827,7.0708723,8.218767,9.366661,10.514555,11.66245,12.533132,13.403813,14.274494,15.141272,16.011953,15.758167,15.504381,15.246691,14.992905,14.739119,12.888432,11.037745,9.187058,7.336372,5.4856853,6.649197,7.8088045,8.968412,10.128019,11.287627,15.9221525,20.556679,25.191204,29.82573,34.464157,36.244568,38.028877,39.809284,41.593597,43.374004,44.908436,46.44677,47.9812,49.51563,51.05006,45.626846,40.20363,34.780415,29.361105,23.937891,20.845604,17.753317,14.661031,11.568744,8.476458,9.386183,10.295909,11.205634,12.11536,13.025085,11.0260315,9.026978,7.0240197,5.024966,3.0259118,3.1079042,3.1898966,3.2718892,3.3538816,3.435874,7.172387,10.9089,14.641508,18.378021,22.11063,23.883228,25.655827,27.428427,29.201025,30.973623,27.162926,23.356134,19.545437,15.734741,11.924045,12.388668,12.849388,13.314012,13.774731,14.239355,16.13299,18.026625,19.924164,21.8178,23.711435,24.500124,25.288813,26.073599,26.862288,27.650976,25.327858,23.004738,20.68162,18.3585,16.039284,15.566852,15.098324,14.625891,14.157363,13.688834,15.309161,16.925583,18.54591,20.166237,21.786564,23.97303,26.15559,28.342056,30.52852,32.711082,30.18103,27.647072,25.113115,22.583063,20.049105,20.439547,20.829987,21.220427,21.610867,22.001307,21.341463,20.68162,20.021774,19.36193,18.698183,16.706938,14.7156925,12.720543,10.729298,8.738052,9.733675,10.729298,11.721016,12.716639,13.712261,14.571229,15.434102,16.29307,17.152039,18.011007,16.972437,15.933866,14.89139,13.852819,12.814248,13.075843,13.341343,13.606842,13.872341,14.13784,14.336966,14.53609,14.739119,14.938243,15.137367,14.688361,14.243259,13.794253,13.349152,12.900145,13.028991,13.16174,13.2905855,13.419431,13.548276,13.993378,14.438479,14.883581,15.328683,15.773785,16.816261,17.854832,18.893402,19.935879,20.97445,21.579632,22.184814,22.789995,23.395178,24.00036,22.696291,21.396124,20.092054,18.791887,17.487818,18.284315,19.080814,19.881216,20.677715,21.474213,21.72019,21.966167,22.20824,22.454218,22.700195,22.23557,21.770947,21.306324,20.8417,20.37317,19.268225,18.163279,17.058334,15.953387,14.848442,15.890917,16.933393,17.975868,19.018343,20.06082,18.569338,17.077856,15.586374,14.090988,12.599506,12.24811,11.900618,11.549222,11.20173,10.850334,10.48332,10.120211,9.753197,9.390087,9.023073,9.0035515,8.980125,8.956698,8.933272,8.913751,9.413514,9.917182,10.42085,10.920613,11.424281,1.3118792,1.3626363,1.4133936,1.4641509,1.5110037,1.5617609,1.5383345,1.5110037,1.4875772,1.4641509,1.43682,1.4485333,1.4641509,1.475864,1.4875772,1.4992905,1.4641509,1.4251068,1.3860629,1.3509232,1.3118792,1.3118792,1.3118792,1.3118792,1.3118792,1.3118792,1.2376955,1.1635119,1.0893283,1.0112402,0.93705654,0.94876975,0.96438736,0.97610056,0.9878138,0.999527,1.0737107,1.1517987,1.2259823,1.3001659,1.3743496,3.8614538,6.348558,8.835662,11.326671,13.813775,11.748346,9.686822,7.6252975,5.563773,3.4983444,3.349977,3.2016098,3.049338,2.900971,2.7486992,2.436347,2.1239948,1.8116426,1.4992905,1.1869383,0.999527,0.81211567,0.62470436,0.43729305,0.24988174,0.22645533,0.19912452,0.1756981,0.14836729,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22645533,0.44900626,0.6754616,0.9019169,1.1244678,1.4251068,1.7257458,2.0263848,2.3231194,2.6237583,3.4241607,4.224563,5.024966,5.825368,6.6257706,6.4110284,6.2001905,5.989353,5.774611,5.563773,5.423215,5.2865605,5.1499066,5.0132523,4.8765984,4.650143,4.423688,4.2011366,3.9746814,3.7482262,4.4002614,5.0483923,5.700427,6.348558,7.000593,8.499884,9.999174,11.498465,13.001659,14.50095,13.950429,13.399908,12.849388,12.298867,11.748346,11.100216,10.44818,9.80005,9.151918,8.499884,8.164105,7.824422,7.4886436,7.1489606,6.813182,6.426646,6.036206,5.64967,5.263134,4.8765984,5.263134,5.64967,6.036206,6.426646,6.813182,6.688241,6.5633,6.4383593,6.3134184,6.1884775,6.086963,5.989353,5.8878384,5.786324,5.688714,5.462259,5.2358036,5.0132523,4.786797,4.564246,4.5369153,4.513489,4.4861584,4.462732,4.4393053,4.5993857,4.7633705,4.9234514,5.087436,5.251421,5.349031,5.4505453,5.548156,5.64967,5.7511845,5.64967,5.548156,5.4505453,5.349031,5.251421,5.337318,5.423215,5.5130157,5.5989127,5.688714,5.036679,4.388548,3.736513,3.0883822,2.436347,2.736986,3.0376248,3.338264,3.638903,3.9356375,4.7516575,5.563773,6.375889,7.1880045,8.00012,7.0630636,6.126007,5.1889505,4.251894,3.310933,5.9620223,8.6131115,11.2642,13.911386,16.562475,14.711788,12.861101,11.014318,9.163632,7.3129454,7.461313,7.6135845,7.7619514,7.914223,8.062591,8.238289,8.413987,8.58578,8.761478,8.937177,8.960603,8.987934,9.01136,9.0386915,9.062118,10.163159,11.2642,12.361338,13.462379,14.56342,15.012426,15.461433,15.914344,16.36335,16.812357,17.487818,18.163279,18.838741,19.514202,20.18576,20.826082,21.4625,22.098917,22.739239,23.375656,28.712975,34.050293,39.38761,44.724926,50.062244,44.350105,38.637966,32.925823,27.213684,21.501543,17.714273,13.927003,10.135828,6.348558,2.5612879,3.0259118,3.4866312,3.951255,4.4119744,4.8765984,5.3256044,5.774611,6.223617,6.676528,7.125534,6.575013,6.0244927,5.473972,4.9234514,4.376835,5.9620223,7.551114,9.136301,10.725393,12.31058,13.138313,13.962143,14.785972,15.613705,16.437534,15.637131,14.836729,14.036326,13.235924,12.439425,15.285735,18.135948,20.986162,23.836376,26.68659,25.1873,23.68801,22.188719,20.689428,19.186234,17.850927,16.511717,15.176412,13.837202,12.501896,13.274967,14.048039,14.825015,15.598087,16.375063,15.449719,14.524376,13.599033,12.67369,11.748346,11.061172,10.373997,9.686822,8.999647,8.312472,8.4257,8.538928,8.648251,8.761478,8.874706,10.612165,12.349625,14.087084,15.824542,17.562002,17.261362,16.960724,16.663988,16.36335,16.062712,14.274494,12.486279,10.698062,8.913751,7.125534,5.7511845,4.376835,2.998581,1.6242313,0.24988174,0.96438736,1.6749885,2.3855898,3.1000953,3.8106966,3.310933,2.8111696,2.3114061,1.8116426,1.3118792,1.0502841,0.78868926,0.5231899,0.26159495,0.0,0.0,0.0,0.0,0.0,0.0,0.113227665,0.22645533,0.3357786,0.44900626,0.5622339,1.1986516,1.8389735,2.475391,3.1118085,3.7482262,3.7638438,3.775557,3.78727,3.7989833,3.8106966,3.4983444,3.1859922,2.87364,2.5612879,2.2489357,2.3738766,2.4988174,2.6237583,2.7486992,2.87364,2.3855898,1.901444,1.4133936,0.92534333,0.43729305,0.698888,0.96438736,1.2259823,1.4875772,1.7491722,1.8116426,1.8741131,1.9365835,1.999054,2.0615244,2.2879796,2.514435,2.736986,2.9634414,3.1859922,2.612045,2.0380979,1.4641509,0.8862993,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.24988174,0.43729305,0.62470436,0.81211567,0.999527,1.6008049,2.1981785,2.7994564,3.4007344,3.998108,5.677001,7.348085,9.026978,10.701966,12.373051,13.349152,14.325252,15.3013525,16.273548,17.24965,16.33602,15.426293,14.512663,13.599033,12.689307,10.998701,9.311999,7.6252975,5.938596,4.251894,5.473972,6.699954,7.9259367,9.151918,10.373997,15.324779,20.27556,25.226343,30.173222,35.124004,36.56082,38.00155,39.438366,40.875187,42.312008,44.32668,46.337444,48.348213,50.362885,52.373653,46.060234,39.75072,33.4373,27.123882,20.81437,18.249176,15.687888,13.1266,10.561408,8.00012,8.999647,9.999174,10.998701,11.998228,13.001659,10.674636,8.351517,6.0244927,3.7013733,1.3743496,1.3626363,1.3509232,1.33921,1.3235924,1.3118792,5.661383,10.010887,14.364296,18.7138,23.063305,25.601166,28.139027,30.67689,33.210846,35.748707,30.325493,24.898373,19.475159,14.048039,8.624825,8.749765,8.874706,8.999647,9.124588,9.249529,11.4633255,13.673217,15.8870125,18.10081,20.310701,22.024733,23.738766,25.448895,27.162926,28.873055,25.987701,23.098444,20.21309,17.323833,14.438479,13.962143,13.4858055,13.013372,12.537036,12.0606985,13.8762455,15.687888,17.49953,19.311174,21.12672,23.789522,26.448421,29.111223,31.774025,34.43683,31.524143,28.61146,25.698776,22.78609,19.873407,20.24823,20.623053,21.00178,21.376602,21.751425,21.411741,21.075964,20.73628,20.400501,20.06082,17.788456,15.51219,13.235924,10.963562,8.687295,9.612638,10.537982,11.4633255,12.388668,13.314012,14.301826,15.285735,16.273548,17.261362,18.249176,17.136421,16.023666,14.9109125,13.798158,12.689307,12.849388,13.013372,13.173453,13.337439,13.501423,13.837202,14.176885,14.512663,14.848442,15.188125,14.875772,14.56342,14.251068,13.938716,13.626364,13.548276,13.4740925,13.399908,13.325725,13.251541,13.700547,14.149553,14.59856,15.051471,15.500477,16.273548,17.050524,17.823597,18.600573,19.373644,20.224804,21.075964,21.923218,22.774378,23.625538,22.29804,20.97445,19.650856,18.32336,16.999767,17.811884,18.623999,19.436115,20.24823,21.06425,21.349272,21.638197,21.923218,22.212145,22.50107,21.98569,21.474213,20.962736,20.45126,19.935879,18.663042,17.386303,16.113468,14.836729,13.563893,14.688361,15.812829,16.937298,18.061766,19.186234,17.86264,16.539047,15.211552,13.887959,12.564366,12.326198,12.08803,11.849861,11.611692,11.373524,10.951848,10.526268,10.100689,9.675109,9.249529,9.163632,9.073831,8.987934,8.898132,8.812236,9.261242,9.714153,10.163159,10.612165,11.061172,1.3118792,1.3665408,1.4172981,1.4680552,1.5227169,1.5734742,1.5500476,1.5266213,1.4992905,1.475864,1.4485333,1.4641509,1.4797685,1.4953861,1.5110037,1.5266213,1.4836729,1.4446288,1.4055848,1.3665408,1.3235924,1.3314011,1.3353056,1.33921,1.3431144,1.3509232,1.2806439,1.2103647,1.1400855,1.0698062,0.999527,0.9956226,0.9956226,0.9917182,0.9917182,0.9878138,1.4719596,1.9561055,2.4441557,2.9283018,3.4124475,5.2045684,6.996689,8.78881,10.58093,12.373051,10.549695,8.726339,6.899079,5.0757227,3.2484627,3.1039999,2.959537,2.815074,2.6706111,2.5261483,2.2840753,2.0380979,1.796025,1.5539521,1.3118792,1.1127546,0.9136301,0.7106012,0.5114767,0.31235218,0.28111696,0.24597734,0.21474212,0.1835069,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19912452,0.39434463,0.59346914,0.78868926,0.9878138,1.2884527,1.5890918,1.8858263,2.1864653,2.4871042,3.3070288,4.126953,4.9468775,5.7668023,6.5867267,6.477403,6.36808,6.2587566,6.1494336,6.036206,5.8292727,5.6223392,5.4154058,5.2084727,5.001539,4.7711797,4.5447245,4.318269,4.0918136,3.8614538,4.493967,5.12648,5.758993,6.3915067,7.0240197,8.179723,9.335425,10.491129,11.6468315,12.798631,12.369146,11.939662,11.510178,11.080693,10.651209,10.163159,9.675109,9.187058,8.699008,8.210958,7.941554,7.6682463,7.394938,7.1216297,6.8483214,6.606249,6.3602715,6.114294,5.8683167,5.6262436,5.930787,6.239235,6.547683,6.8561306,7.1606736,7.094299,7.0240197,6.9537406,6.883461,6.813182,6.699954,6.5867267,6.473499,6.364176,6.250948,5.9737353,5.6965227,5.4193106,5.138193,4.860981,4.775084,4.689187,4.5993857,4.513489,4.423688,4.630621,4.83365,5.040583,5.2436123,5.4505453,5.7238536,6.001066,6.2743745,6.551587,6.824895,6.699954,6.575013,6.4500723,6.3251314,6.2001905,6.1181984,6.04011,5.958118,5.8800297,5.801942,5.196759,4.5954814,3.9942036,3.3890212,2.787743,2.9868677,3.1859922,3.3890212,3.5881457,3.78727,4.5408196,5.298274,6.0518236,6.8092775,7.562827,6.89127,6.223617,5.55206,4.884407,4.21285,6.2314262,8.246098,10.264673,12.28325,14.301826,13.571702,12.841579,12.111456,11.381332,10.651209,10.331048,10.010887,9.690726,9.370565,9.050405,9.565785,10.081166,10.596548,11.111929,11.623405,11.572648,11.521891,11.46723,11.416472,11.361811,12.28325,13.200784,14.122223,15.043662,15.961197,16.41801,16.870922,17.327738,17.780647,18.237463,19.065197,19.89293,20.720663,21.548395,22.37613,23.160913,23.9457,24.730484,25.515268,26.300053,30.879917,35.45978,40.039646,44.61951,49.19937,43.76835,38.34123,32.910206,27.479183,22.048159,18.526388,15.004618,11.482847,7.9610763,4.4393053,4.7907014,5.1460023,5.5013027,5.8566036,6.211904,6.46569,6.715572,6.969358,7.223144,7.47693,6.9342184,6.3915067,5.8487945,5.3060827,4.7633705,6.1181984,7.473026,8.827853,10.182681,11.537509,12.845484,14.153459,15.461433,16.769407,18.073479,17.085665,16.093946,15.1061325,14.114414,13.1266,15.371632,17.616663,19.861694,22.106726,24.351757,23.242907,22.134056,21.02911,19.92026,18.81141,17.991486,17.167656,16.343828,15.523903,14.700074,15.090515,15.480955,15.871395,16.261835,16.64837,15.9104395,15.168603,14.430671,13.688834,12.950902,12.185639,11.424281,10.662923,9.901564,9.136301,9.600925,10.061645,10.526268,10.986988,11.4516115,13.25935,15.070992,16.87873,18.690374,20.498112,19.365835,18.233559,17.101282,15.969006,14.836729,13.833297,12.825961,11.82253,10.819098,9.811763,8.32809,6.8483214,5.364649,3.8809757,2.4012074,2.7213683,3.0415294,3.3616903,3.6818514,3.998108,3.5959544,3.1898966,2.7838387,2.3816853,1.9756275,1.5812829,1.1869383,0.78868926,0.39434463,0.0,0.0,0.0,0.0,0.0,0.0,0.12103647,0.24597734,0.3670138,0.48805028,0.61299115,1.1517987,1.6906061,2.233318,2.7721257,3.310933,3.2875066,3.2640803,3.2367494,3.213323,3.1859922,2.9283018,2.6706111,2.416825,2.1591344,1.901444,2.077142,2.2567444,2.4324427,2.6081407,2.787743,2.3855898,1.9834363,1.5812829,1.1791295,0.77307165,0.9917182,1.2103647,1.4290112,1.6437533,1.8623998,1.9443923,2.0224805,2.1005683,2.182561,2.260649,2.3894942,2.5183394,2.6432803,2.7721257,2.900971,2.455869,2.0146716,1.5734742,1.1283722,0.6871748,0.60127795,0.5114767,0.42557985,0.3357786,0.24988174,0.5192855,0.78868926,1.0580931,1.3314011,1.6008049,2.2059872,2.8111696,3.416352,4.0215344,4.6267166,6.4969254,8.36323,10.2334385,12.103647,13.973856,14.50095,15.024139,15.551234,16.074425,16.601519,15.457528,14.313539,13.173453,12.029464,10.889378,9.694631,8.503788,7.309041,6.1181984,4.9234514,6.3993154,7.8751793,9.351044,10.826907,12.298867,17.128613,21.954454,26.784199,31.61004,36.435883,37.732143,39.028404,40.320763,41.617023,42.913284,44.0807,45.24812,46.415535,47.58295,48.750366,42.88205,37.013733,31.145416,25.281004,19.412687,17.608854,15.801116,13.997282,12.193448,10.38571,10.436467,10.487225,10.537982,10.588739,10.6355915,8.94889,7.2582836,5.5676775,3.8770714,2.1864653,2.9087796,3.6271896,4.3455997,5.067914,5.786324,9.6243515,13.462379,17.300406,21.138433,24.976461,27.16683,29.361105,31.551476,33.74575,35.93612,31.68032,27.428427,23.172626,18.916828,14.661031,14.992905,15.320874,15.652749,15.980719,16.312593,18.647425,20.982258,23.317091,25.651922,27.986755,28.923813,29.856964,30.79402,31.727173,32.66423,30.067802,27.471375,24.87885,22.282423,19.685997,19.151093,18.61619,18.081287,17.546383,17.01148,18.163279,19.318983,20.470781,21.62258,22.774378,25.0116,27.248823,29.486046,31.723269,33.964394,31.293783,28.627077,25.960371,23.293663,20.623053,20.728472,20.829987,20.931501,21.036919,21.138433,21.16186,21.181383,21.20481,21.228235,21.251661,19.018343,16.785025,14.551707,12.318389,10.088976,10.6355915,11.186112,11.736633,12.287154,12.837675,13.548276,14.262781,14.973383,15.687888,16.398489,16.023666,15.648844,15.274021,14.899199,14.524376,14.512663,14.50095,14.489237,14.473619,14.461906,14.231546,13.997282,13.766922,13.532659,13.298394,13.325725,13.349152,13.376482,13.399908,13.423335,13.493614,13.563893,13.634172,13.704452,13.774731,14.204215,14.629795,15.059279,15.484859,15.914344,16.394585,16.87873,17.358973,17.843119,18.32336,19.07691,19.83046,20.58401,21.333654,22.087204,21.275087,20.462973,19.650856,18.838741,18.026625,18.577147,19.13157,19.682093,20.236517,20.787037,21.165764,21.54449,21.919313,22.29804,22.67677,22.161386,21.646006,21.130625,20.615244,20.099863,18.948065,17.800169,16.64837,15.500477,14.348679,15.473146,16.601519,17.725986,18.850454,19.974922,18.74113,17.503435,16.269644,15.035853,13.798158,13.2905855,12.779109,12.271536,11.760059,11.248583,10.944039,10.6355915,10.327144,10.018696,9.714153,9.585307,9.456462,9.331521,9.202676,9.073831,9.362757,9.651682,9.936704,10.22563,10.510651,1.3118792,1.3665408,1.4212024,1.475864,1.53443,1.5890918,1.5617609,1.5383345,1.5110037,1.4875772,1.4641509,1.4797685,1.4992905,1.5149081,1.53443,1.5500476,1.5070993,1.4641509,1.4212024,1.3782539,1.33921,1.3470187,1.358732,1.3665408,1.3782539,1.3860629,1.3235924,1.2572175,1.1908426,1.1283722,1.0619974,1.0463798,1.0268579,1.0112402,0.9917182,0.97610056,1.8702087,2.7643168,3.6584249,4.5564375,5.4505453,6.547683,7.6448197,8.741957,9.839094,10.936231,9.351044,7.7619514,6.1767645,4.5876727,2.998581,2.8619268,2.7213683,2.5808098,2.4402514,2.2996929,2.1278992,1.9561055,1.7843118,1.6086137,1.43682,1.2259823,1.0112402,0.80040246,0.58566034,0.37482262,0.3357786,0.29673457,0.25378615,0.21474212,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1717937,0.339683,0.5114767,0.679366,0.8511597,1.1517987,1.4485333,1.7491722,2.0498111,2.35045,3.1898966,4.029343,4.8687897,5.708236,6.551587,6.5437784,6.5359693,6.5281606,6.520352,6.5125427,6.2353306,5.958118,5.6809053,5.4036927,5.12648,4.8961205,4.6657605,4.435401,4.2050414,3.9746814,4.591577,5.2045684,5.8214636,6.434455,7.0513506,7.859562,8.671678,9.479889,10.2881,11.100216,10.791768,10.479416,10.170968,9.858616,9.550168,9.226103,8.898132,8.574067,8.250002,7.9259367,7.719003,7.5081654,7.3012323,7.094299,6.8873653,6.785851,6.6843367,6.578918,6.477403,6.375889,6.602344,6.8287997,7.0591593,7.2856145,7.5120697,7.4964523,7.480835,7.4691215,7.453504,7.437886,7.3129454,7.1880045,7.0630636,6.9381227,6.813182,6.481308,6.153338,5.8214636,5.493494,5.1616197,5.0132523,4.860981,4.7126136,4.564246,4.4119744,4.661856,4.9078336,5.153811,5.4036927,5.64967,6.098676,6.551587,7.000593,7.4495993,7.898606,7.7502384,7.601871,7.4495993,7.3012323,7.1489606,6.902983,6.6531014,6.407124,6.1611466,5.911265,5.35684,4.802415,4.2479897,3.6935644,3.1391394,3.2367494,3.338264,3.435874,3.5373883,3.638903,4.3338866,5.0327744,5.7316628,6.426646,7.125534,6.7233806,6.321227,5.919074,5.5169206,5.1108627,6.4969254,7.882988,9.269051,10.651209,12.037272,12.427712,12.818152,13.208592,13.599033,13.989473,13.196879,12.408191,11.615597,10.826907,10.0382185,10.893282,11.748346,12.603411,13.458474,14.313539,14.180789,14.051944,13.923099,13.794253,13.661504,14.40334,15.141272,15.883108,16.62104,17.362877,17.823597,18.284315,18.74113,19.20185,19.662569,20.642574,21.62258,22.602585,23.58259,24.562595,25.495747,26.4289,27.358147,28.291298,29.224451,33.04686,36.86927,40.69168,44.51409,48.3365,43.1905,38.044495,32.89459,27.748587,22.59868,19.34241,16.086138,12.825961,9.56969,6.3134184,6.559396,6.8092775,7.055255,7.3012323,7.551114,7.605776,7.660437,7.715099,7.7697606,7.824422,7.289519,6.754616,6.2197127,5.6848097,5.1499066,6.2743745,7.394938,8.519405,9.639969,10.764437,12.552653,14.34087,16.13299,17.921206,19.713327,18.534197,17.351164,16.172033,14.992905,13.813775,15.453624,17.093473,18.733322,20.37317,22.01302,21.298513,20.58401,19.865599,19.151093,18.436588,18.12814,17.823597,17.515148,17.206701,16.898252,16.906061,16.909966,16.91387,16.921679,16.925583,16.371159,15.816733,15.258404,14.703979,14.149553,13.314012,12.4745655,11.639023,10.799577,9.964035,10.77615,11.588266,12.400381,13.212498,14.024612,15.906535,17.788456,19.674282,21.556206,23.438128,21.474213,19.506393,17.542479,15.578565,13.610746,13.388195,13.165645,12.943093,12.724447,12.501896,10.9089,9.319808,7.7307167,6.141625,4.548629,4.478349,4.4041657,4.3338866,4.2597027,4.1894236,3.8770714,3.5686235,3.2562714,2.9478238,2.639376,2.1083772,1.5812829,1.0541886,0.5270943,0.0,0.0,0.0,0.0,0.0,0.0,0.13274968,0.26549935,0.39824903,0.5309987,0.6637484,1.1049459,1.5461433,1.9912452,2.4324427,2.87364,2.8111696,2.7486992,2.6862288,2.6237583,2.5612879,2.358259,2.1591344,1.9561055,1.7530766,1.5500476,1.7804074,2.0107672,2.241127,2.4714866,2.7018464,2.3816853,2.0654287,1.7491722,1.4290112,1.1127546,1.2845483,1.456342,1.6281357,1.8038338,1.9756275,2.0732377,2.1708477,2.2684577,2.366068,2.463678,2.4910088,2.522244,2.5534792,2.5808098,2.612045,2.3035975,1.9912452,1.6827974,1.3743496,1.0619974,0.93705654,0.81211567,0.6871748,0.5622339,0.43729305,0.78868926,1.1439898,1.4953861,1.8467822,2.1981785,2.8111696,3.4202564,4.029343,4.6384296,5.251421,7.3168497,9.378374,11.443803,13.509232,15.57466,15.648844,15.726933,15.801116,15.875299,15.949483,14.579038,13.204688,11.834243,10.459893,9.085544,8.39056,7.6916723,6.996689,6.297801,5.5989127,7.3246584,9.050405,10.77615,12.501896,14.223738,18.928543,23.633347,28.342056,33.04686,37.751667,38.903465,40.055264,41.20706,42.35886,43.51066,43.834724,44.15879,44.47895,44.803017,45.123177,39.703865,34.28065,28.857437,23.434223,18.011007,16.964628,15.918248,14.871868,13.821584,12.775204,11.873287,10.975275,10.073358,9.175345,8.273428,7.2192397,6.165051,5.1108627,4.056674,2.998581,4.4510183,5.903456,7.355894,8.8083315,10.260769,13.58732,16.91387,20.236517,23.563068,26.885714,28.7364,30.583183,32.429966,34.27675,36.12353,33.03905,29.954575,26.870096,23.785618,20.701141,21.236044,21.770947,22.305851,22.840754,23.375656,25.831526,28.291298,30.747168,33.20694,35.66281,35.818985,35.979065,36.135242,36.29142,36.4515,34.147903,31.844305,29.540707,27.241014,24.937418,24.343948,23.746574,23.153105,22.555733,21.962263,22.454218,22.946173,23.438128,23.933987,24.425941,26.237583,28.049225,29.860868,31.676416,33.48806,31.063425,28.642694,26.218061,23.79733,21.376602,21.20481,21.036919,20.865126,20.693333,20.525442,20.908073,21.290705,21.673336,22.05597,22.4386,20.24823,18.057861,15.867491,13.677121,11.486752,11.66245,11.838148,12.013845,12.185639,12.361338,12.798631,13.235924,13.673217,14.11051,14.551707,14.9109125,15.274021,15.637131,16.00024,16.36335,16.175938,15.988527,15.801116,15.613705,15.426293,14.621986,13.821584,13.017277,12.216875,11.412568,11.775677,12.138786,12.501896,12.861101,13.224211,13.438952,13.653695,13.868437,14.0831785,14.301826,14.703979,15.110037,15.516094,15.918248,16.324306,16.515621,16.706938,16.894348,17.085665,17.273075,17.929016,18.584955,19.240894,19.896833,20.548868,20.24823,19.951496,19.650856,19.350218,19.049578,19.34241,19.635239,19.92807,20.2209,20.51373,20.978354,21.446882,21.91541,22.383938,22.848562,22.333181,21.813896,21.298513,20.779228,20.263847,19.23699,18.214037,17.18718,16.164225,15.137367,16.261835,17.386303,18.51077,19.639143,20.76361,19.615717,18.471727,17.327738,16.183748,15.035853,14.254972,13.4740925,12.689307,11.908427,11.123642,10.936231,10.744915,10.553599,10.366188,10.174872,10.006983,9.839094,9.671205,9.503315,9.339331,9.464272,9.589212,9.714153,9.839094,9.964035,1.3118792,1.3704453,1.4290112,1.4836729,1.542239,1.6008049,1.5734742,1.5500476,1.5266213,1.4992905,1.475864,1.4953861,1.5149081,1.53443,1.5539521,1.5734742,1.5305257,1.4836729,1.4407244,1.3938715,1.3509232,1.3665408,1.3782539,1.3938715,1.4094892,1.4251068,1.3665408,1.3040704,1.2455044,1.1869383,1.1244678,1.0932326,1.0580931,1.0268579,0.9956226,0.96438736,2.2684577,3.5725281,4.8765984,6.180669,7.4886436,7.890797,8.292951,8.695104,9.097258,9.499411,8.148487,6.801469,5.4505453,4.0996222,2.7486992,2.6159496,2.4792955,2.3465457,2.2098918,2.0732377,1.9717231,1.8702087,1.7686942,1.6632754,1.5617609,1.33921,1.1127546,0.8862993,0.6637484,0.43729305,0.39044023,0.3435874,0.29673457,0.24597734,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14055848,0.28502136,0.42557985,0.5700427,0.7106012,1.0112402,1.3118792,1.6125181,1.9131571,2.2137961,3.0727646,3.9317331,4.7907014,5.6535745,6.5125427,6.606249,6.703859,6.7975645,6.89127,6.98888,6.6413884,6.2938967,5.9464045,5.5989127,5.251421,5.017157,4.786797,4.552533,4.318269,4.087909,4.6852827,5.282656,5.8800297,6.477403,7.0747766,7.5394006,8.0040245,8.468649,8.933272,9.4018,9.2104845,9.019169,8.831758,8.640442,8.449126,8.289046,8.125061,7.9610763,7.800996,7.6370106,7.4964523,7.3519893,7.211431,7.066968,6.9264097,6.9654536,7.0044975,7.043542,7.08649,7.125534,7.2739015,7.4183645,7.5667315,7.715099,7.8634663,7.90251,7.941554,7.9805984,8.023546,8.062591,7.9259367,7.7892823,7.648724,7.5120697,7.375416,6.9927845,6.610153,6.2275214,5.84489,5.462259,5.251421,5.036679,4.825841,4.6110992,4.4002614,4.689187,4.9781127,5.270943,5.559869,5.8487945,6.473499,7.098203,7.726812,8.351517,8.976221,8.800523,8.624825,8.449126,8.273428,8.101635,7.6838636,7.269997,6.8561306,6.4383593,6.0244927,5.5169206,5.009348,4.5017757,3.9942036,3.4866312,3.4866312,3.4866312,3.4866312,3.4866312,3.4866312,4.126953,4.7672753,5.407597,6.0479193,6.688241,6.551587,6.4188375,6.282183,6.1494336,6.012779,6.7663293,7.5159745,8.269524,9.023073,9.776623,11.283723,12.794726,14.30573,15.816733,17.323833,16.066616,14.805493,13.544372,12.28325,11.0260315,12.220779,13.415526,14.610273,15.80502,16.999767,16.792833,16.585901,16.378967,16.168129,15.961197,16.52343,17.08176,17.643993,18.202324,18.760653,19.229181,19.693806,20.158428,20.623053,21.087677,22.219954,23.35223,24.484507,25.616783,26.74906,27.83058,28.908194,29.989714,31.071234,32.14885,35.213802,38.27876,41.343716,44.408672,47.473625,42.60874,37.74386,32.87897,28.014086,23.1492,20.158428,17.163752,14.17298,11.178304,8.187531,8.32809,8.468649,8.609207,8.745861,8.886419,8.745861,8.601398,8.460839,8.316377,8.175818,7.648724,7.1216297,6.590631,6.0635366,5.5364423,6.426646,7.3168497,8.207053,9.097258,9.987461,12.259823,14.532186,16.804546,19.07691,21.349272,19.978827,18.608381,17.24184,15.871395,14.50095,15.535617,16.570284,17.60495,18.639616,19.674282,19.354122,19.030056,18.705992,18.38583,18.061766,18.268698,18.475632,18.68647,18.893402,19.100336,18.72161,18.338978,17.96025,17.581524,17.198893,16.831879,16.46096,16.090042,15.719124,15.348206,14.438479,13.524849,12.611219,11.701493,10.787864,11.951375,13.110983,14.274494,15.438006,16.601519,18.553719,20.509825,22.46593,24.41813,26.374237,23.578686,20.779228,17.983677,15.18422,12.388668,12.946998,13.509232,14.067561,14.625891,15.188125,13.48971,11.791295,10.096785,8.398369,6.699954,6.2353306,5.7707067,5.3060827,4.841459,4.376835,4.1581883,3.9434462,3.7287042,3.513962,3.2992198,2.639376,1.979532,1.319688,0.659844,0.0,0.0,0.0,0.0,0.0,0.0,0.14055848,0.28502136,0.42557985,0.5700427,0.7106012,1.0580931,1.4016805,1.7491722,2.0927596,2.436347,2.338737,2.2372224,2.135708,2.0380979,1.9365835,1.7882162,1.6437533,1.4953861,1.3470187,1.1986516,1.4836729,1.7647898,2.0459068,2.330928,2.612045,2.3816853,2.1474214,1.9131571,1.6827974,1.4485333,1.5773785,1.7062237,1.8311646,1.9600099,2.0888553,2.2020829,2.3192148,2.4324427,2.5456703,2.6628022,2.5964274,2.5261483,2.4597735,2.3933985,2.3231194,2.1474214,1.9717231,1.7921207,1.6164225,1.43682,1.2767396,1.1127546,0.94876975,0.78868926,0.62470436,1.0580931,1.4953861,1.9287747,2.366068,2.7994564,3.416352,4.029343,4.646239,5.2592297,5.8761253,8.136774,10.393518,12.654168,14.914817,17.175465,16.800642,16.42582,16.050997,15.676175,15.3013525,13.696643,12.095839,10.491129,8.890324,7.2856145,7.08649,6.883461,6.6804323,6.477403,6.2743745,8.250002,10.22563,12.201257,14.176885,16.148607,20.732376,25.316145,29.896008,34.479774,39.063545,40.07088,41.08212,42.09336,43.100697,44.11194,43.588745,43.06946,42.546272,42.023083,41.499893,36.52178,31.543665,26.565554,21.591345,16.613232,16.324306,16.031475,15.74255,15.453624,15.160794,13.314012,11.4633255,9.612638,7.7619514,5.911265,5.493494,5.0718184,4.6540475,4.2323723,3.8106966,5.997162,8.183627,10.366188,12.552653,14.739119,17.550287,20.361458,23.176533,25.987701,28.79887,30.302067,31.805262,33.308456,34.81165,36.31094,34.397785,32.48072,30.567566,28.650503,26.737347,27.479183,28.217115,28.958952,29.696884,30.43872,33.01953,35.596436,38.177246,40.758057,43.338863,42.718063,42.097263,41.476463,40.855667,40.23877,38.228,36.217236,34.206467,32.1957,30.188839,29.532898,28.876959,28.22102,27.568985,26.913044,26.745155,26.577267,26.409376,26.241488,26.073599,27.463566,28.849628,30.235691,31.625658,33.011723,30.833065,28.658312,26.479656,24.300999,22.126247,21.681147,21.239948,20.79875,20.35365,19.91245,20.654287,21.396124,22.141865,22.883701,23.625538,21.478117,19.330696,17.183275,15.035853,12.888432,12.689307,12.486279,12.287154,12.08803,11.888905,12.0489855,12.212971,12.376955,12.537036,12.70102,13.798158,14.899199,16.00024,17.101282,18.19842,17.839214,17.476105,17.112995,16.749886,16.386776,15.016331,13.641981,12.271536,10.897186,9.526741,10.22563,10.924518,11.623405,12.326198,13.025085,13.384291,13.743496,14.106606,14.465811,14.825015,15.207646,15.590279,15.97291,16.355541,16.738173,16.636658,16.531239,16.429726,16.32821,16.226696,16.78112,17.33945,17.89778,18.45611,19.014439,19.225277,19.436115,19.650856,19.861694,20.076437,20.107672,20.138906,20.174046,20.205282,20.236517,20.794846,21.353176,21.911505,22.46593,23.02426,22.504974,21.98569,21.466404,20.943214,20.423927,19.525915,18.623999,17.725986,16.82407,15.926057,17.050524,18.174992,19.29946,20.423927,21.548395,20.494207,19.44002,18.38583,17.331642,16.273548,15.21936,14.165172,13.110983,12.056794,10.998701,10.928422,10.8542385,10.783959,10.709775,10.6355915,10.4286585,10.221725,10.0147915,9.807858,9.600925,9.561881,9.526741,9.487698,9.448653,9.413514,1.3118792,1.3743496,1.4329157,1.4914817,1.5539521,1.6125181,1.5890918,1.5617609,1.5383345,1.5110037,1.4875772,1.5110037,1.53443,1.5539521,1.5773785,1.6008049,1.5539521,1.5031948,1.456342,1.4094892,1.3626363,1.3821584,1.4016805,1.4212024,1.4407244,1.4641509,1.4055848,1.3509232,1.2962615,1.2415999,1.1869383,1.1400855,1.0932326,1.0463798,0.9956226,0.94876975,2.6667068,4.380739,6.094772,7.8088045,9.526741,9.2339115,8.941081,8.648251,8.355421,8.062591,6.949836,5.8370814,4.7243266,3.611572,2.4988174,2.3699722,2.241127,2.1083772,1.979532,1.8506867,1.815547,1.7843118,1.7530766,1.7218413,1.6867018,1.4485333,1.2142692,0.97610056,0.737932,0.4997635,0.44510186,0.39044023,0.3357786,0.28111696,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.113227665,0.23035973,0.3435874,0.46071947,0.57394713,0.8745861,1.175225,1.475864,1.7765031,2.0732377,2.9556324,3.8341231,4.716518,5.5950084,6.473499,6.6726236,6.871748,7.066968,7.266093,7.461313,7.043542,6.6257706,6.211904,5.794133,5.376362,5.138193,4.903929,4.6696653,4.435401,4.2011366,4.7789884,5.3607445,5.938596,6.520352,7.098203,7.2192397,7.3402762,7.461313,7.578445,7.699481,7.629202,7.558923,7.4886436,7.4183645,7.348085,7.348085,7.348085,7.348085,7.348085,7.348085,7.2739015,7.195813,7.1177254,7.039637,6.9615493,7.1450562,7.328563,7.5081654,7.6916723,7.8751793,7.941554,8.011833,8.078208,8.144583,8.210958,8.308568,8.402273,8.495979,8.59359,8.687295,8.538928,8.386656,8.238289,8.086017,7.9376497,7.504261,7.066968,6.6335793,6.196286,5.7628975,5.4856853,5.212377,4.939069,4.661856,4.388548,4.7204223,5.0522966,5.3841705,5.716045,6.0518236,6.8483214,7.648724,8.449126,9.249529,10.049932,9.850807,9.651682,9.448653,9.249529,9.050405,8.468649,7.8868923,7.3012323,6.719476,6.13772,5.677001,5.2162814,4.755562,4.298747,3.8380275,3.736513,3.638903,3.5373883,3.435874,3.338264,3.9200199,4.5017757,5.083532,5.6691923,6.250948,6.3836975,6.5164475,6.649197,6.7819467,6.910792,7.0318284,7.152865,7.2739015,7.3910336,7.5120697,10.143637,12.771299,15.402867,18.034433,20.662096,18.932447,17.202797,15.473146,13.743496,12.013845,13.548276,15.0827055,16.617136,18.151566,19.685997,19.400974,19.115953,18.830933,18.54591,18.26089,18.64352,19.022247,19.400974,19.783606,20.162333,20.630861,21.103294,21.571823,22.044254,22.512783,23.79733,25.08188,26.366428,27.650976,28.93943,30.165411,31.391394,32.62128,33.847263,35.073246,37.38075,39.688248,41.99575,44.303253,46.610756,42.03089,37.44712,32.863354,28.28349,23.699722,20.97445,18.245272,15.516094,12.790822,10.061645,10.096785,10.128019,10.159255,10.194394,10.22563,9.885946,9.546264,9.20658,8.866898,8.52331,8.0040245,7.4847393,6.9654536,6.446168,5.9268827,6.5828223,7.238762,7.898606,8.554545,9.21439,11.966993,14.723501,17.476105,20.232613,22.98912,21.42736,19.869503,18.307743,16.745981,15.188125,15.617609,16.047092,16.476578,16.906061,17.335546,17.405825,17.476105,17.546383,17.616663,17.686943,18.409256,19.13157,19.853886,20.5762,21.298513,20.53325,19.771893,19.00663,18.241367,17.476105,17.288692,17.105186,16.921679,16.734268,16.55076,15.562947,14.575133,13.58732,12.599506,11.611692,13.1266,14.637604,16.148607,17.663515,19.174519,21.200905,23.231194,25.257578,27.283962,29.314253,25.683159,22.052063,18.420969,14.79378,11.162686,12.5058,13.848915,15.188125,16.531239,17.874353,16.07052,14.2666855,12.458947,10.655114,8.85128,7.9923115,7.1333427,6.278279,5.4193106,4.564246,4.4432096,4.322173,4.2011366,4.084005,3.9629683,3.1703746,2.377781,1.5851873,0.79259366,0.0,0.0,0.0,0.0,0.0,0.0,0.15227169,0.30454338,0.45681506,0.60908675,0.76135844,1.0112402,1.2572175,1.5031948,1.7530766,1.999054,1.8623998,1.7257458,1.5890918,1.4485333,1.3118792,1.2181735,1.1283722,1.0346665,0.94096094,0.8511597,1.1869383,1.5188124,1.8545911,2.1903696,2.5261483,2.377781,2.2294137,2.0810463,1.9365835,1.7882162,1.8702087,1.9522011,2.0341935,2.1161861,2.1981785,2.330928,2.463678,2.5964274,2.7291772,2.8619268,2.697942,2.533957,2.366068,2.2020829,2.0380979,1.9912452,1.9482968,1.901444,1.8584955,1.8116426,1.6125181,1.4133936,1.2142692,1.0112402,0.81211567,1.3314011,1.8467822,2.366068,2.8814487,3.4007344,4.0215344,4.6384296,5.2592297,5.8800297,6.5008297,8.956698,11.408664,13.864532,16.320402,18.77627,17.948538,17.124708,16.300879,15.473146,14.649317,12.818152,10.986988,9.151918,7.320754,5.4856853,5.7785153,6.0713453,6.364176,6.657006,6.949836,9.175345,11.400854,13.626364,15.851873,18.073479,22.53621,26.995037,31.453865,35.916595,40.375423,41.242203,42.10898,42.975754,43.846436,44.713215,43.346672,41.976227,40.609688,39.24315,37.876606,33.343594,28.810585,24.277573,19.744562,15.211552,15.680079,16.148607,16.613232,17.08176,17.550287,14.750832,11.951375,9.148014,6.348558,3.5491016,3.7638438,3.978586,4.193328,4.40807,4.6267166,7.5433054,10.459893,13.376482,16.296974,19.213564,21.513256,23.81295,26.112642,28.412334,30.712029,31.871635,33.02734,34.186947,35.342648,36.498352,35.756516,35.010777,34.265034,33.519295,32.773552,33.71842,34.663284,35.612053,36.55692,37.501785,40.20363,42.905476,45.607323,48.30917,51.011017,49.61324,48.219368,46.82159,45.423817,44.02604,42.3081,40.590164,38.87223,37.154293,35.436356,34.721848,34.007343,33.29284,32.57833,31.863827,31.036093,30.20836,29.380627,28.552895,27.72516,28.685644,29.65003,30.614418,31.574902,32.539288,30.60661,28.673931,26.741251,24.808573,22.875893,22.161386,21.446882,20.728472,20.013966,19.29946,20.404406,21.505447,22.60649,23.711435,24.812477,22.708004,20.60353,18.499058,16.394585,14.286208,13.712261,13.138313,12.564366,11.986515,11.412568,11.29934,11.186112,11.076789,10.963562,10.850334,12.689307,14.524376,16.36335,18.19842,20.037392,19.498585,18.963682,18.424873,17.886066,17.351164,15.406772,13.466284,11.521891,9.581403,7.6370106,8.675582,9.714153,10.748819,11.787391,12.825961,13.329629,13.833297,14.34087,14.844538,15.348206,15.711315,16.07052,16.429726,16.788929,17.148134,16.75379,16.359446,15.965101,15.570756,15.176412,15.633226,16.093946,16.554665,17.015385,17.476105,18.19842,18.924637,19.650856,20.37317,21.09939,20.872934,20.646479,20.416119,20.189665,19.96321,20.61134,21.25947,21.903696,22.551826,23.199959,22.67677,22.153578,21.634293,21.111103,20.587914,19.810938,19.037865,18.26089,17.487818,16.710842,17.839214,18.963682,20.08815,21.212618,22.337086,21.372698,20.40831,19.443924,18.475632,17.511244,16.183748,14.856251,13.528754,12.201257,10.87376,10.920613,10.963562,11.010414,11.053363,11.100216,10.8542385,10.604357,10.358379,10.108498,9.86252,9.663396,9.464272,9.261242,9.062118,8.862993,1.3118792,1.3743496,1.43682,1.4992905,1.5617609,1.6242313,1.6008049,1.5734742,1.5500476,1.5266213,1.4992905,1.5266213,1.5500476,1.5734742,1.6008049,1.6242313,1.5734742,1.5266213,1.475864,1.4251068,1.3743496,1.4016805,1.4251068,1.4485333,1.475864,1.4992905,1.4485333,1.4016805,1.3509232,1.3001659,1.2494087,1.1869383,1.1244678,1.0619974,0.999527,0.93705654,3.0610514,5.1889505,7.3129454,9.43694,11.560935,10.573121,9.589212,8.601398,7.6135845,6.6257706,5.7511845,4.8765984,3.998108,3.1235218,2.2489357,2.1239948,1.999054,1.8741131,1.7491722,1.6242313,1.6632754,1.698415,1.737459,1.7765031,1.8116426,1.5617609,1.3118792,1.0619974,0.81211567,0.5622339,0.4997635,0.43729305,0.37482262,0.31235218,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.737932,1.038571,1.33921,1.6359446,1.9365835,2.8385005,3.736513,4.6384296,5.5364423,6.4383593,6.7389984,7.0357327,7.336372,7.6370106,7.9376497,7.4495993,6.9615493,6.473499,5.989353,5.5013027,5.263134,5.024966,4.786797,4.548629,4.3143644,4.8765984,5.4388323,6.001066,6.5633,7.125534,6.899079,6.676528,6.4500723,6.223617,6.001066,6.0518236,6.098676,6.1494336,6.2001905,6.250948,6.4110284,6.575013,6.7389984,6.899079,7.0630636,7.0513506,7.0357327,7.0240197,7.012306,7.000593,7.3246584,7.648724,7.9766936,8.300759,8.624825,8.6131115,8.601398,8.58578,8.574067,8.562354,8.710721,8.862993,9.01136,9.163632,9.311999,9.151918,8.987934,8.823949,8.663869,8.499884,8.011833,7.523783,7.0357327,6.551587,6.0635366,5.7238536,5.388075,5.0483923,4.7126136,4.376835,4.7516575,5.12648,5.5013027,5.8761253,6.250948,7.223144,8.1992445,9.175345,10.151445,11.123642,10.901091,10.674636,10.44818,10.22563,9.999174,9.249529,8.499884,7.7502384,7.000593,6.250948,5.8370814,5.423215,5.0132523,4.5993857,4.1894236,3.9863946,3.78727,3.5881457,3.3890212,3.1859922,3.7130866,4.2362766,4.7633705,5.2865605,5.813655,6.211904,6.6140575,7.012306,7.4105554,7.812709,7.3012323,6.785851,6.2743745,5.7628975,5.251421,8.999647,12.751778,16.500004,20.24823,24.00036,21.798277,19.6001,17.398016,15.199838,13.001659,14.875772,16.749886,18.623999,20.498112,22.37613,22.01302,21.64991,21.2868,20.92369,20.560583,20.76361,20.962736,21.16186,21.360985,21.564014,22.036446,22.512783,22.98912,23.461554,23.937891,25.37471,26.811531,28.24835,29.689075,31.125895,32.500244,33.874596,35.248943,36.623295,38.00155,39.551594,41.101643,42.65169,44.201736,45.751785,41.449135,37.150387,32.85164,28.548988,24.250242,21.786564,19.326792,16.863113,14.399435,11.935758,11.861574,11.787391,11.713207,11.639023,11.560935,11.0260315,10.487225,9.948417,9.413514,8.874706,8.36323,7.8517528,7.336372,6.824895,6.3134184,6.7389984,7.1606736,7.5862536,8.011833,8.437413,11.674163,14.9109125,18.151566,21.388315,24.625065,22.875893,21.12672,19.373644,17.624472,15.875299,15.699601,15.523903,15.348206,15.176412,15.000713,15.461433,15.926057,16.386776,16.8514,17.31212,18.549814,19.78751,21.025206,22.262901,23.500597,22.348799,21.200905,20.049105,18.90121,17.749413,17.749413,17.749413,17.749413,17.749413,17.749413,16.687416,15.625418,14.56342,13.501423,12.439425,14.301826,16.164225,18.026625,19.889025,21.751425,23.851994,25.948658,28.049225,30.149794,32.250362,27.78763,23.3249,18.862167,14.399435,9.936704,12.0606985,14.188598,16.312593,18.436588,20.560583,18.651329,16.738173,14.825015,12.911859,10.998701,9.749292,8.499884,7.250475,6.001066,4.7516575,4.7243266,4.7009,4.6735697,4.650143,4.6267166,3.7013733,2.77603,1.8506867,0.92534333,0.0,0.0,0.0,0.0,0.0,0.0,0.1639849,0.3240654,0.48805028,0.6481308,0.81211567,0.96438736,1.1127546,1.261122,1.4133936,1.5617609,1.3860629,1.2142692,1.038571,0.8628729,0.6871748,0.6481308,0.61299115,0.57394713,0.5388075,0.4997635,0.8862993,1.2767396,1.6632754,2.0498111,2.436347,2.3738766,2.3114061,2.2489357,2.1864653,2.1239948,2.1630387,2.1981785,2.2372224,2.2762666,2.3114061,2.463678,2.612045,2.7643168,2.912684,3.0610514,2.7994564,2.5378613,2.2762666,2.0107672,1.7491722,1.8389735,1.9248703,2.0107672,2.1005683,2.1864653,1.9482968,1.7140326,1.475864,1.2376955,0.999527,1.6008049,2.1981785,2.7994564,3.4007344,3.998108,4.6267166,5.251421,5.8761253,6.5008297,7.125534,9.776623,12.423808,15.074897,17.725986,20.37317,19.100336,17.823597,16.55076,15.274021,14.001186,11.935758,9.874233,7.812709,5.7511845,3.6857557,4.474445,5.263134,6.0518236,6.8366084,7.6252975,10.100689,12.576079,15.051471,17.526861,19.998348,24.33614,28.673931,33.011723,37.34951,41.6873,42.41352,43.135838,43.862057,44.588272,45.31059,43.100697,40.8869,38.673103,36.46321,34.249416,30.161507,26.073599,21.98569,17.901684,13.813775,15.035853,16.261835,17.487818,18.7138,19.935879,16.187653,12.439425,8.687295,4.939069,1.1869383,2.0380979,2.8892577,3.736513,4.5876727,5.4388323,9.089449,12.73616,16.386776,20.037392,23.68801,25.476225,27.260536,29.048752,30.83697,32.625187,33.4373,34.249416,35.06153,35.87365,36.685764,37.111343,37.536922,37.9625,38.388084,38.813663,39.961555,41.113358,42.26125,43.413048,44.560944,47.38773,50.210613,53.0374,55.86419,58.68707,56.512318,54.337566,52.162815,49.988064,47.81331,46.388203,44.963097,43.53799,42.112885,40.687775,39.9108,39.13773,38.360752,37.58768,36.810703,35.323128,33.839455,32.351875,30.8643,29.376722,29.911625,30.450434,30.98924,31.524143,32.06295,30.37625,28.685644,26.998941,25.31224,23.625538,22.637724,21.64991,20.662096,19.674282,18.68647,20.15062,21.610867,23.075018,24.539167,25.999414,23.937891,21.876366,19.810938,17.749413,15.687888,14.739119,13.786445,12.837675,11.888905,10.936231,10.549695,10.163159,9.776623,9.386183,8.999647,11.576552,14.149553,16.72646,19.29946,21.876366,21.16186,20.45126,19.736753,19.026152,18.311647,15.801116,13.286681,10.77615,8.261715,5.7511845,7.125534,8.499884,9.874233,11.248583,12.626837,13.274967,13.923099,14.575133,15.223265,15.875299,16.211079,16.55076,16.88654,17.226223,17.562002,16.874826,16.187653,15.500477,14.813302,14.126127,14.489237,14.848442,15.211552,15.57466,15.93777,17.175465,18.41316,19.650856,20.888552,22.126247,21.638197,21.150146,20.662096,20.174046,19.685997,20.423927,21.16186,21.899792,22.637724,23.375656,22.848562,22.325373,21.798277,21.275087,20.751898,20.099863,19.451733,18.799696,18.151566,17.49953,18.623999,19.748466,20.876839,22.001307,23.125774,22.251188,21.376602,20.498112,19.623526,18.74894,17.148134,15.551234,13.950429,12.349625,10.748819,10.912805,11.076789,11.23687,11.400854,11.560935,11.275913,10.986988,10.698062,10.413041,10.124115,9.761005,9.4018,9.0386915,8.675582,8.312472,1.3509232,1.4016805,1.456342,1.5070993,1.5617609,1.6125181,1.5890918,1.5656652,1.5461433,1.5227169,1.4992905,1.5188124,1.5383345,1.5617609,1.5812829,1.6008049,1.5461433,1.4953861,1.4407244,1.3899672,1.33921,1.3704453,1.4016805,1.43682,1.4680552,1.4992905,1.4719596,1.4446288,1.4172981,1.3899672,1.3626363,1.2806439,1.1986516,1.116659,1.0307622,0.94876975,3.3655949,5.786324,8.203149,10.619974,13.036799,11.6351185,10.2334385,8.831758,7.426173,6.0244927,5.3138914,4.5993857,3.8887846,3.174279,2.463678,2.2723622,2.0810463,1.893635,1.7023194,1.5110037,1.5305257,1.5461433,1.5656652,1.5812829,1.6008049,1.4094892,1.2181735,1.0307622,0.8394465,0.6481308,0.5622339,0.47633708,0.38653582,0.30063897,0.21083772,0.1717937,0.12884527,0.08589685,0.042948425,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07027924,0.14055848,0.21083772,0.28111696,0.3513962,0.59346914,0.8355421,1.077615,1.319688,1.5617609,2.541766,3.5178664,4.493967,5.473972,6.4500723,6.621866,6.7897553,6.9615493,7.1294384,7.3012323,6.871748,6.4383593,6.008875,5.579391,5.1499066,4.9624953,4.775084,4.5876727,4.4002614,4.21285,4.7516575,5.2865605,5.825368,6.364176,6.899079,6.703859,6.504734,6.3056097,6.1103897,5.911265,5.9229784,5.930787,5.9425,5.9542136,5.9620223,6.1064854,6.2470436,6.3915067,6.532065,6.676528,6.602344,6.5281606,6.4578815,6.3836975,6.3134184,6.66091,7.012306,7.363703,7.7111945,8.062591,8.082112,8.101635,8.121157,8.140678,8.164105,8.398369,8.632633,8.866898,9.101162,9.339331,9.14411,8.952794,8.761478,8.566258,8.374943,8.007929,7.6409154,7.2739015,6.9068875,6.5359693,6.211904,5.8878384,5.563773,5.2358036,4.911738,5.298274,5.688714,6.0752497,6.461786,6.8483214,7.890797,8.933272,9.975748,11.018223,12.0606985,12.056794,12.05289,12.0489855,12.041177,12.037272,11.39695,10.752724,10.108498,9.468176,8.823949,8.175818,7.523783,6.8756523,6.223617,5.575486,5.2865605,5.001539,4.7126136,4.423688,4.138666,4.630621,5.12648,5.6223392,6.1181984,6.6140575,6.969358,7.328563,7.6838636,8.043069,8.398369,8.078208,7.7541428,7.433982,7.1099167,6.785851,9.679013,12.572175,15.465338,18.3585,21.251661,20.092054,18.936352,17.776743,16.62104,15.461433,17.136421,18.807507,20.47859,22.153578,23.824663,23.660677,23.496693,23.328804,23.164818,23.000834,23.188246,23.37956,23.570877,23.758287,23.949604,24.17606,24.39861,24.625065,24.85152,25.074072,26.182922,27.29177,28.396717,29.505568,30.614418,32.48072,34.35093,36.221138,38.091347,39.961555,40.85176,41.741966,42.632168,43.522373,44.412575,40.234867,36.057156,31.879444,27.701735,23.524023,21.591345,19.658665,17.725986,15.793307,13.860628,14.176885,14.493141,14.809398,15.12175,15.438006,14.438479,13.442857,12.44333,11.447707,10.44818,9.741484,9.034787,8.32809,7.621393,6.910792,7.1216297,7.328563,7.535496,7.7424297,7.9493628,10.526268,13.103174,15.683984,18.26089,20.837795,19.639143,18.444397,17.245745,16.047092,14.848442,14.711788,14.575133,14.438479,14.301826,14.161267,14.754736,15.348206,15.941674,16.531239,17.124708,18.3585,19.596195,20.829987,22.063778,23.301472,22.223858,21.150146,20.076437,18.998821,17.92511,17.620567,17.316025,17.01148,16.706938,16.398489,15.594183,14.789876,13.985569,13.181262,12.373051,14.379913,16.386776,18.389734,20.396597,22.399555,23.453745,24.504028,25.558218,26.608501,27.66269,25.03893,22.411268,19.78751,17.163752,14.53609,15.250595,15.961197,16.675701,17.386303,18.10081,17.112995,16.125181,15.137367,14.149553,13.16174,12.412095,11.66245,10.912805,10.163159,9.413514,8.273428,7.1333427,5.9932575,4.853172,3.7130866,2.97125,2.233318,1.4914817,0.75354964,0.011713207,0.015617609,0.015617609,0.019522011,0.023426414,0.023426414,0.1756981,0.3318742,0.48414588,0.63641757,0.78868926,1.0737107,1.3626363,1.6515622,1.9365835,2.2255092,2.05762,1.8897307,1.7218413,1.5539521,1.3860629,1.3274968,1.2689307,1.2064602,1.1478943,1.0893283,1.475864,1.8663043,2.2567444,2.6471848,3.0376248,2.8970666,2.7565079,2.6159496,2.4792955,2.338737,2.4090161,2.4831998,2.5534792,2.6276627,2.7018464,2.7213683,2.7447948,2.7682211,2.7916477,2.8111696,2.5886188,2.366068,2.1435168,1.9209659,1.698415,2.0888553,2.4792955,2.8697357,3.260176,3.6506162,3.521771,3.3890212,3.260176,3.1313305,2.998581,3.7599394,4.521298,5.278752,6.04011,6.801469,7.1333427,7.465217,7.7970915,8.128965,8.460839,10.522364,12.583888,14.641508,16.703033,18.760653,17.50734,16.254026,14.996809,13.743496,12.486279,10.819098,9.151918,7.4847393,5.8175592,4.1503797,5.1108627,6.0713453,7.0318284,7.988407,8.94889,11.951375,14.949956,17.948538,20.951023,23.949604,27.233206,30.516808,33.796505,37.08011,40.363712,41.88643,43.413048,44.935764,46.462387,47.98901,44.084606,40.18411,36.279705,32.379208,28.474806,25.503555,22.53621,19.56496,16.59371,13.626364,14.555612,15.488764,16.421915,17.355068,18.28822,15.453624,12.622932,9.788337,6.957645,4.126953,5.8566036,7.5862536,9.315904,11.045554,12.775204,15.8870125,18.998821,22.114534,25.226343,28.338152,29.493855,30.645653,31.801357,32.957058,34.112762,35.073246,36.03373,36.994213,37.95079,38.911274,39.293903,39.676537,40.059166,40.4418,40.82443,41.67559,42.52675,43.374004,44.225163,45.076324,47.251076,49.425827,51.60058,53.775333,55.950085,54.279,52.61182,50.940735,49.269653,47.598568,46.618565,45.634655,44.650745,43.67074,42.68683,41.456944,40.227055,38.99717,37.767284,36.537395,35.21771,33.89802,32.57833,31.258644,29.938957,30.454338,30.965815,31.481195,31.996576,32.51196,30.610514,28.712975,26.811531,24.91399,23.012547,21.82561,20.642574,19.455637,18.272602,17.085665,18.514675,19.943687,21.368793,22.797804,24.226816,22.723621,21.220427,19.717232,18.214037,16.710842,15.867491,15.024139,14.176885,13.333533,12.486279,11.927949,11.365715,10.807385,10.249056,9.686822,11.66245,13.638077,15.613705,17.585428,19.561056,19.315079,19.069101,18.81922,18.573242,18.32336,16.378967,14.430671,12.482374,10.534078,8.58578,9.390087,10.194394,10.994797,11.799104,12.599506,13.032895,13.466284,13.895767,14.329156,14.762545,15.133463,15.5082855,15.879204,16.254026,16.624945,15.801116,14.981192,14.157363,13.333533,12.513609,12.8650055,13.216402,13.571702,13.923099,14.274494,15.320874,16.36335,17.409729,18.45611,19.498585,19.400974,19.303364,19.205755,19.108145,19.014439,19.635239,20.256039,20.880743,21.501543,22.126247,21.630388,21.13453,20.63867,20.146715,19.650856,19.256512,18.858263,18.463919,18.069574,17.675228,18.772366,19.869503,20.96664,22.063778,23.160913,22.325373,21.485926,20.650383,19.810938,18.975395,17.573715,16.175938,14.774258,13.376482,11.974802,11.955279,11.935758,11.916236,11.896713,11.873287,11.443803,11.014318,10.584834,10.155351,9.725866,9.499411,9.269051,9.042596,8.81614,8.58578,1.3860629,1.4290112,1.4719596,1.5149081,1.5578566,1.6008049,1.5812829,1.5617609,1.5383345,1.5188124,1.4992905,1.5149081,1.5305257,1.5461433,1.5617609,1.5734742,1.5188124,1.4641509,1.4094892,1.3548276,1.3001659,1.33921,1.3782539,1.4212024,1.4602464,1.4992905,1.4953861,1.4914817,1.4836729,1.4797685,1.475864,1.3743496,1.2689307,1.1674163,1.0659018,0.96438736,3.6740425,6.3836975,9.093353,11.803008,14.512663,12.693212,10.877665,9.058213,7.2426662,5.423215,4.8765984,4.3260775,3.775557,3.2250361,2.6745155,2.4207294,2.1669433,1.9092526,1.6554666,1.4016805,1.397776,1.3938715,1.3938715,1.3899672,1.3860629,1.2572175,1.1283722,0.9956226,0.8667773,0.737932,0.62470436,0.5114767,0.39824903,0.28892577,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10541886,0.15617609,0.21083772,0.26159495,0.44900626,0.63251317,0.8160201,1.0034313,1.1869383,2.241127,3.2992198,4.3534083,5.407597,6.461786,6.5008297,6.5437784,6.5828223,6.621866,6.66091,6.289992,5.919074,5.5442514,5.173333,4.7985106,4.661856,4.5252023,4.388548,4.251894,4.1113358,4.6267166,5.138193,5.64967,6.1611466,6.676528,6.504734,6.336845,6.165051,5.9932575,5.825368,5.794133,5.7668023,5.735567,5.704332,5.6730967,5.7980375,5.919074,6.044015,6.165051,6.2860875,6.153338,6.0205884,5.891743,5.758993,5.6262436,6.001066,6.375889,6.7507114,7.125534,7.5003567,7.551114,7.605776,7.656533,7.7111945,7.7619514,8.082112,8.402273,8.722435,9.042596,9.362757,9.140205,8.917655,8.695104,8.472553,8.250002,8.0040245,7.7541428,7.5081654,7.2582836,7.012306,6.699954,6.387602,6.0752497,5.7628975,5.4505453,5.8487945,6.250948,6.649197,7.0513506,7.4495993,8.55845,9.671205,10.780055,11.888905,13.001659,13.216402,13.431144,13.645885,13.860628,14.07537,13.540467,13.005564,12.470661,11.935758,11.400854,10.510651,9.6243515,8.738052,7.8517528,6.9615493,6.5867267,6.211904,5.8370814,5.462259,5.087436,5.55206,6.016684,6.481308,6.9459314,7.4105554,7.726812,8.043069,8.359325,8.671678,8.987934,8.855185,8.722435,8.589685,8.456935,8.324185,10.358379,12.396477,14.430671,16.464865,18.499058,18.38583,18.268698,18.15547,18.038338,17.92511,19.393166,20.865126,22.333181,23.805141,25.273195,25.308336,25.339571,25.370806,25.405945,25.437181,25.616783,25.796385,25.975988,26.15559,26.339098,26.311768,26.28834,26.26101,26.237583,26.214157,26.991133,27.768108,28.545084,29.322062,30.099037,32.465103,34.831173,37.193336,39.559402,41.925472,42.15583,42.386192,42.61655,42.84691,43.073364,39.020596,34.96392,30.911152,26.854479,22.801708,21.396124,19.994444,18.592764,17.191084,15.789403,16.492195,17.198893,17.901684,18.608381,19.311174,17.854832,16.398489,14.938243,13.481901,12.025558,11.123642,10.221725,9.315904,8.413987,7.5120697,7.504261,7.492548,7.480835,7.473026,7.461313,9.378374,11.29934,13.216402,15.133463,17.050524,16.406298,15.758167,15.113941,14.469715,13.825488,13.723974,13.626364,13.524849,13.423335,13.325725,14.048039,14.770353,15.492668,16.214983,16.937298,18.171087,19.400974,20.634766,21.868557,23.098444,22.098917,21.09939,20.099863,19.100336,18.10081,17.491722,16.87873,16.269644,15.660558,15.051471,14.50095,13.954333,13.407718,12.861101,12.31058,14.461906,16.609327,18.756748,20.90417,23.05159,23.055496,23.0594,23.063305,23.071114,23.075018,22.286327,21.501543,20.712854,19.924164,19.13938,18.436588,17.7377,17.03881,16.33602,15.637131,15.57466,15.51219,15.449719,15.387249,15.324779,15.074897,14.825015,14.575133,14.325252,14.07537,11.818625,9.565785,7.309041,5.056201,2.7994564,2.2450314,1.6906061,1.1361811,0.58175594,0.023426414,0.031235218,0.03513962,0.039044023,0.046852827,0.05075723,0.19131571,0.3357786,0.47633708,0.62079996,0.76135844,1.1869383,1.6125181,2.0380979,2.463678,2.8892577,2.7291772,2.5690966,2.4090161,2.2489357,2.0888553,2.0068626,1.9209659,1.8389735,1.756981,1.6749885,2.069333,2.4597735,2.854118,3.2445583,3.638903,3.4202564,3.2016098,2.9868677,2.7682211,2.5495746,2.6588979,2.7643168,2.87364,2.979059,3.0883822,2.9829633,2.8775444,2.7721257,2.6667068,2.5612879,2.3816853,2.1981785,2.0146716,1.8311646,1.6515622,2.3426414,3.0337205,3.7287042,4.4197836,5.1108627,5.0913405,5.067914,5.044488,5.0210614,5.001539,5.919074,6.8405128,7.7619514,8.679486,9.600925,9.639969,9.679013,9.721962,9.761005,9.80005,11.272009,12.740065,14.208119,15.680079,17.148134,15.914344,14.6805525,13.446761,12.209065,10.975275,9.702439,8.429605,7.1567693,5.883934,4.6110992,5.743376,6.8756523,8.011833,9.14411,10.276386,13.802062,17.323833,20.849508,24.375183,27.900858,30.126368,32.35578,34.58129,36.810703,39.036213,41.36324,43.686356,46.013382,48.3365,50.663525,45.068516,39.47741,33.886307,28.291298,22.700195,20.845604,18.994917,17.14423,15.289639,13.438952,14.079274,14.7156925,15.356014,15.996336,16.636658,14.723501,12.806439,10.893282,8.976221,7.0630636,9.671205,12.28325,14.89139,17.503435,20.111576,22.688482,25.261482,27.838388,30.411388,32.988297,33.511486,34.03077,34.55396,35.07715,35.600338,36.70919,37.814137,38.922985,40.031837,41.136784,41.476463,41.816147,42.15583,42.49942,42.8391,43.38572,43.936237,44.48676,45.03728,45.5878,47.11442,48.63714,50.16376,51.686478,53.213097,52.04568,50.88217,49.71866,48.551243,47.38773,46.848923,46.30621,45.767403,45.228596,44.685883,43.003086,41.316383,39.633587,37.946884,36.264088,35.108383,33.956585,32.804787,31.652988,30.50119,30.993145,31.4851,31.977055,32.46901,32.960964,30.848682,28.7364,26.624119,24.511837,22.399555,21.017397,19.635239,18.25308,16.870922,15.488764,16.87873,18.272602,19.666473,21.056442,22.450314,21.509352,20.564487,19.623526,18.678661,17.7377,16.995863,16.25793,15.516094,14.778163,14.036326,13.306203,12.572175,11.838148,11.108025,10.373997,11.748346,13.1266,14.50095,15.875299,17.24965,17.468296,17.683039,17.901684,18.12033,18.338978,16.95682,15.570756,14.188598,12.806439,11.424281,11.654641,11.885,12.11536,12.34572,12.576079,12.790822,13.005564,13.220306,13.435048,13.64979,14.055848,14.465811,14.871868,15.281831,15.687888,14.73131,13.770826,12.814248,11.85767,10.901091,11.240774,11.584361,11.927949,12.271536,12.611219,13.466284,14.317443,15.168603,16.023666,16.874826,17.167656,17.460487,17.753317,18.046146,18.338978,18.84655,19.354122,19.861694,20.369267,20.876839,20.40831,19.943687,19.479063,19.014439,18.549814,18.409256,18.268698,18.12814,17.991486,17.850927,18.920732,19.99054,21.060347,22.130152,23.199959,22.399555,21.599154,20.79875,19.998348,19.20185,17.999294,16.800642,15.598087,14.399435,13.200784,12.997755,12.794726,12.591698,12.388668,12.185639,11.615597,11.04165,10.471607,9.897659,9.323712,9.2339115,9.140205,9.0465,8.956698,8.862993,1.4251068,1.456342,1.4914817,1.5227169,1.5539521,1.5890918,1.5695697,1.5539521,1.53443,1.5188124,1.4992905,1.5110037,1.5188124,1.5305257,1.5383345,1.5500476,1.4914817,1.43682,1.3782539,1.319688,1.261122,1.3118792,1.358732,1.4055848,1.4524376,1.4992905,1.5188124,1.53443,1.5539521,1.5695697,1.5890918,1.4641509,1.3431144,1.2181735,1.097137,0.97610056,3.978586,6.9810715,9.983557,12.986042,15.988527,13.755209,11.521891,9.288573,7.0591593,4.825841,4.4393053,4.0488653,3.6623292,3.2757936,2.8892577,2.5690966,2.2489357,1.9287747,1.6086137,1.2884527,1.2650263,1.2415999,1.2181735,1.1986516,1.175225,1.1049459,1.0346665,0.96438736,0.8941081,0.8238289,0.6871748,0.5505207,0.41386664,0.27330816,0.13665408,0.10932326,0.08199245,0.05466163,0.027330816,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.30063897,0.42948425,0.5583295,0.6832704,0.81211567,1.9443923,3.076669,4.2089458,5.3412223,6.473499,6.3836975,6.2938967,6.2040954,6.114294,6.0244927,5.708236,5.395884,5.0796275,4.7633705,4.4510183,4.3612175,4.2753205,4.1894236,4.0996222,4.0137253,4.5017757,4.985922,5.473972,5.9620223,6.4500723,6.3056097,6.165051,6.0205884,5.8800297,5.735567,5.6691923,5.5989127,5.5286336,5.4583545,5.388075,5.4895897,5.591104,5.6965227,5.7980375,5.899552,5.708236,5.5169206,5.3217,5.1303844,4.939069,5.337318,5.735567,6.13772,6.5359693,6.9381227,7.0240197,7.1060123,7.191909,7.277806,7.363703,7.7658563,8.171914,8.577971,8.98403,9.386183,9.136301,8.882515,8.628729,8.378847,8.125061,7.996216,7.871275,7.7424297,7.6135845,7.4886436,7.1880045,6.8873653,6.5867267,6.2860875,5.989353,6.3993154,6.813182,7.223144,7.6370106,8.050878,9.226103,10.405232,11.584361,12.759586,13.938716,14.372105,14.809398,15.242786,15.676175,16.113468,15.683984,15.258404,14.828919,14.40334,13.973856,12.849388,11.72492,10.600452,9.475985,8.351517,7.8868923,7.426173,6.9615493,6.5008297,6.036206,6.473499,6.9068875,7.3441806,7.7775693,8.210958,8.484266,8.757574,9.030883,9.304191,9.573594,9.63216,9.690726,9.749292,9.803954,9.86252,11.04165,12.216875,13.396004,14.571229,15.750359,16.675701,17.60495,18.534197,19.459541,20.388788,21.653814,22.922745,24.191677,25.456703,26.725634,26.955994,27.186354,27.416712,27.643167,27.873528,28.04532,28.213211,28.385004,28.556799,28.724688,28.45138,28.174168,27.900858,27.623646,27.350338,27.799343,28.244446,28.693453,29.138554,29.58756,32.445583,35.30751,38.169437,41.02746,43.889385,43.455997,43.026512,42.597027,42.167545,41.73806,37.806328,33.87069,29.938957,26.007223,22.07549,21.200905,20.330223,19.455637,18.584955,17.714273,18.807507,19.900738,20.997875,22.091108,23.188246,21.271183,19.354122,17.433157,15.516094,13.599033,12.501896,11.404759,10.307622,9.2104845,8.113348,7.8868923,7.656533,7.4300776,7.2036223,6.9732623,8.234385,9.491602,10.748819,12.006037,13.263254,13.169549,13.075843,12.986042,12.892336,12.798631,12.73616,12.67369,12.611219,12.548749,12.486279,13.341343,14.192502,15.043662,15.8987255,16.749886,17.979773,19.20966,20.439547,21.669432,22.899319,21.973976,21.048632,20.12329,19.20185,18.276506,17.358973,16.445343,15.531713,14.614178,13.700547,13.411622,13.118792,12.829865,12.54094,12.24811,14.539994,16.831879,19.119858,21.411741,23.699722,22.657246,21.61477,20.572296,19.52982,18.487345,19.537628,20.587914,21.638197,22.688482,23.738766,21.626484,19.514202,17.398016,15.285735,13.173453,14.036326,14.899199,15.762072,16.624945,17.487818,17.7377,17.987581,18.237463,18.487345,18.737226,15.367727,11.998228,8.628729,5.2592297,1.8858263,1.5188124,1.1478943,0.77697605,0.40605783,0.039044023,0.046852827,0.05075723,0.058566034,0.06637484,0.07418364,0.20693332,0.339683,0.47243267,0.60518235,0.737932,1.3001659,1.8623998,2.4246337,2.9868677,3.5491016,3.39683,3.2445583,3.0922866,2.9400148,2.787743,2.6823244,2.5769055,2.4714866,2.366068,2.260649,2.6588979,3.0532427,3.4475873,3.8419318,4.2362766,3.9434462,3.6467118,3.3538816,3.057147,2.7643168,2.9048753,3.049338,3.1898966,3.3343596,3.474918,3.240654,3.0102942,2.77603,2.5456703,2.3114061,2.1708477,2.0263848,1.8858263,1.7413634,1.6008049,2.5964274,3.5881457,4.5837684,5.579391,6.575013,6.66091,6.746807,6.8287997,6.914696,7.000593,8.078208,9.159728,10.241247,11.318862,12.400381,12.146595,11.896713,11.642927,11.389141,11.139259,12.01775,12.89624,13.778636,14.657126,15.535617,14.321347,13.107079,11.892809,10.67854,9.464272,8.58578,7.70729,6.8287997,5.9542136,5.0757227,6.379793,7.6838636,8.991838,10.295909,11.599979,15.648844,19.701614,23.750479,27.799343,31.84821,33.023434,34.194756,35.366077,36.5413,37.71262,40.836143,43.96357,47.08709,50.210613,53.33804,46.056328,38.77462,31.489004,24.207294,16.925583,16.191557,15.453624,14.719597,13.985569,13.251541,13.599033,13.946525,14.294017,14.641508,14.989,13.989473,12.993851,11.994324,10.998701,9.999174,13.48971,16.980246,20.470781,23.961317,27.451853,29.486046,31.524143,33.56224,35.600338,37.63844,37.529114,37.415886,37.306564,37.19724,37.087917,38.34123,39.598446,40.85176,42.10898,43.362293,43.659027,43.95576,44.2564,44.553135,44.84987,45.09975,45.349632,45.599514,45.849396,46.099277,46.97386,47.84845,48.72694,49.601524,50.476112,49.81627,49.156425,48.496582,47.836735,47.17689,47.07928,46.981674,46.884064,46.786453,46.688843,44.54923,42.405712,40.2661,38.126488,35.986877,35.002968,34.01906,33.031242,32.047333,31.063425,31.531952,32.004387,32.47291,32.94144,33.413876,31.086851,28.763731,26.436708,24.113588,21.786564,20.209187,18.627903,17.04662,15.469242,13.887959,15.246691,16.601519,17.96025,19.318983,20.67381,20.291178,19.908546,19.525915,19.143284,18.760653,18.12814,17.491722,16.85921,16.222792,15.586374,14.6805525,13.778636,12.872814,11.966993,11.061172,11.838148,12.611219,13.388195,14.161267,14.938243,15.621513,16.300879,16.98415,17.66742,18.35069,17.530766,16.714746,15.8987255,15.078801,14.262781,13.919194,13.575606,13.235924,12.892336,12.548749,12.548749,12.544845,12.54094,12.54094,12.537036,12.978233,13.423335,13.864532,14.30573,14.750832,13.657599,12.564366,11.471134,10.381805,9.288573,9.620447,9.952321,10.284196,10.61607,10.951848,11.611692,12.271536,12.93138,13.591225,14.251068,14.934339,15.613705,16.296974,16.980246,17.663515,18.053955,18.448301,18.838741,19.233086,19.623526,19.190138,18.756748,18.319456,17.886066,17.448774,17.565907,17.679134,17.796265,17.909492,18.026625,19.069101,20.111576,21.15405,22.196527,23.239002,22.47374,21.712381,20.951023,20.18576,19.4244,18.424873,17.425346,16.42582,15.426293,14.426766,14.040231,13.653695,13.271063,12.884527,12.501896,11.783486,11.06898,10.354475,9.639969,8.925464,8.968412,9.01136,9.054309,9.093353,9.136301,1.4641509,1.4836729,1.5070993,1.5305257,1.5539521,1.5734742,1.5617609,1.5461433,1.5305257,1.5149081,1.4992905,1.5031948,1.5110037,1.5149081,1.5188124,1.5266213,1.4641509,1.4055848,1.3431144,1.2845483,1.2259823,1.2806439,1.3353056,1.3899672,1.4446288,1.4992905,1.5383345,1.5812829,1.620327,1.6593709,1.698415,1.5578566,1.4133936,1.2728351,1.1283722,0.9878138,4.283129,7.578445,10.87376,14.169076,17.464392,14.813302,12.166118,9.518932,6.871748,4.224563,3.998108,3.775557,3.5491016,3.3265507,3.1000953,2.7135596,2.330928,1.9443923,1.5617609,1.175225,1.1322767,1.0893283,1.0463798,1.0034313,0.96438736,0.95267415,0.94096094,0.93315214,0.92143893,0.9136301,0.74964523,0.58566034,0.42557985,0.26159495,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.15617609,0.22645533,0.29673457,0.3670138,0.43729305,1.6476578,2.8580225,4.068387,5.278752,6.4891167,6.266566,6.0479193,5.8292727,5.606722,5.388075,5.1303844,4.872694,4.6150036,4.357313,4.0996222,4.0605783,4.025439,3.9863946,3.951255,3.912211,4.376835,4.8375545,5.298274,5.7628975,6.223617,6.1103897,5.9932575,5.8800297,5.7668023,5.64967,5.5403466,5.4310236,5.3217,5.2084727,5.099149,5.181142,5.263134,5.349031,5.4310236,5.5130157,5.2592297,5.009348,4.755562,4.5017757,4.251894,4.6735697,5.099149,5.5247293,5.950309,6.375889,6.493021,6.610153,6.727285,6.844417,6.9615493,7.453504,7.941554,8.433509,8.921559,9.413514,9.128492,8.847376,8.566258,8.281238,8.00012,7.9923115,7.984503,7.9766936,7.968885,7.9610763,7.676055,7.387129,7.098203,6.813182,6.524256,6.949836,7.375416,7.800996,8.226576,8.648251,9.893755,11.139259,12.384764,13.630268,14.875772,15.531713,16.183748,16.839687,17.495626,18.151566,17.831406,17.511244,17.191084,16.870922,16.55076,15.188125,13.825488,12.4628525,11.100216,9.737579,9.187058,8.636538,8.086017,7.5394006,6.98888,7.3910336,7.7970915,8.203149,8.609207,9.01136,9.24172,9.47208,9.702439,9.932799,10.163159,10.409137,10.6590185,10.904996,11.150972,11.400854,11.721016,12.041177,12.361338,12.681499,13.001659,14.969479,16.941202,18.90902,20.880743,22.848562,23.914463,24.980366,26.046267,27.108265,28.174168,28.603651,29.02923,29.458715,29.884295,30.31378,30.47386,30.63394,30.79402,30.954102,31.114182,30.587088,30.063898,29.536802,29.013613,28.486519,28.603651,28.720783,28.84182,28.958952,29.076084,32.429966,35.783848,39.141632,42.495514,45.849396,44.760067,43.67074,42.58141,41.48818,40.39885,36.588154,32.78136,28.970665,25.159967,21.349272,21.005684,20.666,20.322414,19.978827,19.639143,21.122816,22.60649,24.094067,25.57774,27.061413,24.683632,22.305851,19.92807,17.554192,15.176412,13.884054,12.591698,11.29934,10.003078,8.710721,8.265619,7.824422,7.37932,6.9342184,6.4891167,7.08649,7.6838636,8.281238,8.878611,9.475985,9.936704,10.393518,10.8542385,11.314958,11.775677,11.748346,11.72492,11.701493,11.674163,11.650736,12.630741,13.614651,14.59856,15.578565,16.562475,17.788456,19.018343,20.244326,21.474213,22.700195,21.849035,21.00178,20.15062,19.29946,18.448301,17.230127,16.011953,14.789876,13.571702,12.349625,12.318389,12.28325,12.252014,12.220779,12.185639,14.621986,17.050524,19.486872,21.919313,24.351757,22.258997,20.170141,18.081287,15.988527,13.899672,16.788929,19.674282,22.563541,25.448895,28.338152,24.812477,21.2868,17.761126,14.239355,10.71368,12.501896,14.286208,16.074425,17.86264,19.650856,20.400501,21.150146,21.899792,22.649437,23.399082,18.912924,14.430671,9.944512,5.4583545,0.97610056,0.78868926,0.60518235,0.42167544,0.23426414,0.05075723,0.058566034,0.07027924,0.078088045,0.08980125,0.10151446,0.22255093,0.3435874,0.46852827,0.58956474,0.7106012,1.4133936,2.1122816,2.8111696,3.513962,4.21285,4.068387,3.9239242,3.775557,3.631094,3.4866312,3.3616903,3.232845,3.1039999,2.979059,2.8502135,3.2484627,3.6467118,4.041056,4.4393053,4.8375545,4.466636,4.0918136,3.7208953,3.3460727,2.9751544,3.1508527,3.330455,3.506153,3.6857557,3.8614538,3.5022488,3.1430438,2.7838387,2.4207294,2.0615244,1.9600099,1.8584955,1.7530766,1.6515622,1.5500476,2.8463092,4.1464753,5.4427366,6.7389984,8.039165,8.23048,8.421796,8.6131115,8.8083315,8.999647,10.241247,11.478943,12.720543,13.958238,15.199838,14.653222,14.11051,13.563893,13.021181,12.4745655,12.763491,13.056321,13.345247,13.634172,13.923099,12.728352,11.533605,10.338858,9.14411,7.9493628,7.4691215,6.984976,6.5008297,6.0205884,5.5364423,7.016211,8.492075,9.971844,11.447707,12.923572,17.49953,22.07549,26.65145,31.223505,35.799465,35.916595,36.03373,36.15086,36.271896,36.38903,40.312954,44.236877,48.1608,52.08863,56.012554,47.040237,38.06792,29.095606,20.12329,11.150972,11.533605,11.916236,12.298867,12.681499,13.06413,13.118792,13.173453,13.228115,13.282777,13.337439,13.25935,13.177358,13.09927,13.017277,12.939189,17.308216,21.677242,26.046267,30.419197,34.788223,36.287514,37.786804,39.286095,40.78929,42.28858,41.546745,40.801003,40.059166,39.31733,38.575493,39.977173,41.378857,42.78444,44.18612,45.5878,45.841587,46.099277,46.353065,46.60685,46.860638,46.81378,46.763027,46.71227,46.66151,46.610756,46.837208,47.063663,47.286217,47.512672,47.73913,47.58295,47.426773,47.2706,47.11833,46.96215,47.305737,47.65323,47.99682,48.344307,48.687897,46.09147,43.498947,40.90252,38.30609,35.713566,34.893642,34.07762,33.261604,32.441677,31.625658,32.07076,32.519768,32.968773,33.413876,33.86288,31.32502,28.787157,26.249296,23.711435,21.173573,19.39707,17.620567,15.844065,14.063657,12.287154,13.610746,14.934339,16.254026,17.57762,18.90121,19.07691,19.256512,19.43221,19.611813,19.78751,19.256512,18.729418,18.19842,17.66742,17.136421,16.058807,14.981192,13.903577,12.825961,11.748346,11.924045,12.099743,12.27544,12.4511385,12.626837,13.770826,14.918721,16.066616,17.21451,18.362404,18.108618,17.858736,17.60495,17.351164,17.101282,16.183748,15.270117,14.356487,13.438952,12.525322,12.306676,12.084125,11.8654785,11.6468315,11.424281,11.900618,12.380859,12.857197,13.333533,13.813775,12.583888,11.357906,10.128019,8.902037,7.676055,7.996216,8.320281,8.644346,8.964508,9.288573,9.753197,10.221725,10.690253,11.158782,11.623405,12.697116,13.770826,14.840633,15.914344,16.988054,17.265266,17.542479,17.819693,18.096905,18.374117,17.96806,17.565907,17.159847,16.75379,16.351637,16.71865,17.08957,17.460487,17.831406,18.19842,19.213564,20.228708,21.243853,22.258997,23.274141,22.551826,21.82561,21.09939,20.37317,19.650856,18.850454,18.05005,17.24965,16.449247,15.648844,15.0827055,14.516567,13.946525,13.380386,12.814248,11.955279,11.096312,10.241247,9.382278,8.52331,8.702912,8.878611,9.058213,9.2339115,9.413514,1.4992905,1.5110037,1.5266213,1.5383345,1.5500476,1.5617609,1.5500476,1.5383345,1.5266213,1.5110037,1.4992905,1.4992905,1.4992905,1.4992905,1.4992905,1.4992905,1.43682,1.3743496,1.3118792,1.2494087,1.1869383,1.2494087,1.3118792,1.3743496,1.43682,1.4992905,1.5617609,1.6242313,1.6867018,1.7491722,1.8116426,1.6515622,1.4875772,1.3235924,1.1635119,0.999527,4.5876727,8.175818,11.763964,15.348206,18.936352,15.875299,12.814248,9.749292,6.688241,3.6232853,3.5608149,3.4983444,3.435874,3.3734035,3.310933,2.8619268,2.4129205,1.9639144,1.5110037,1.0619974,0.999527,0.93705654,0.8745861,0.81211567,0.74964523,0.80040246,0.8511597,0.9019169,0.94876975,0.999527,0.81211567,0.62470436,0.43729305,0.24988174,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,1.3509232,2.639376,3.9239242,5.212377,6.5008297,6.1494336,5.801942,5.4505453,5.099149,4.7516575,4.548629,4.349504,4.1503797,3.951255,3.7482262,3.7638438,3.775557,3.78727,3.7989833,3.8106966,4.251894,4.689187,5.12648,5.563773,6.001066,5.911265,5.825368,5.735567,5.64967,5.563773,5.4115014,5.263134,5.1108627,4.9624953,4.814128,4.8765984,4.939069,5.001539,5.0640097,5.12648,4.814128,4.5017757,4.1894236,3.873167,3.5608149,4.0137253,4.462732,4.911738,5.3607445,5.813655,5.9620223,6.114294,6.262661,6.4110284,6.5633,7.137247,7.7111945,8.289046,8.862993,9.43694,9.124588,8.812236,8.499884,8.187531,7.8751793,7.988407,8.101635,8.210958,8.324185,8.437413,8.164105,7.8868923,7.6135845,7.336372,7.0630636,7.5003567,7.9376497,8.374943,8.812236,9.249529,10.561408,11.873287,13.189071,14.50095,15.812829,16.687416,17.562002,18.436588,19.311174,20.18576,19.974922,19.764084,19.549341,19.338505,19.123762,17.526861,15.926057,14.325252,12.724447,11.123642,10.487225,9.850807,9.21439,8.574067,7.9376497,8.312472,8.687295,9.062118,9.43694,9.811763,9.999174,10.186585,10.373997,10.561408,10.748819,11.186112,11.623405,12.0606985,12.501896,12.939189,12.400381,11.861574,11.326671,10.787864,10.249056,13.263254,16.273548,19.287746,22.301945,25.31224,26.175114,27.037985,27.900858,28.763731,29.626604,30.251308,30.876013,31.500717,32.125423,32.750126,32.898495,33.050766,33.19913,33.351402,33.49977,32.7267,31.949724,31.176653,30.399675,29.626604,29.411861,29.201025,28.986282,28.775444,28.560703,32.41435,36.264088,40.11383,43.96357,47.81331,46.064137,44.31106,42.56189,40.812717,39.063545,35.373886,31.68813,27.998468,24.312714,20.623053,20.81437,21.00178,21.189192,21.376602,21.564014,23.438128,25.31224,27.186354,29.064371,30.938484,28.099983,25.261482,22.422981,19.588387,16.749886,15.262308,13.774731,12.287154,10.799577,9.311999,8.648251,7.988407,7.3246584,6.66091,6.001066,5.938596,5.8761253,5.813655,5.7511845,5.688714,6.699954,7.7111945,8.726339,9.737579,10.748819,10.764437,10.77615,10.787864,10.799577,10.81129,11.924045,13.036799,14.149553,15.262308,16.375063,17.601046,18.823124,20.049105,21.275087,22.50107,21.724094,20.951023,20.174046,19.400974,18.623999,17.101282,15.57466,14.048039,12.525322,10.998701,11.225157,11.4516115,11.674163,11.900618,12.123169,14.700074,17.273075,19.849981,22.426888,24.999887,21.860748,18.725513,15.586374,12.4511385,9.311999,14.036326,18.760653,23.488884,28.213211,32.93754,27.998468,23.063305,18.124235,13.189071,8.250002,10.963562,13.673217,16.386776,19.100336,21.813896,23.063305,24.312714,25.562122,26.811531,28.06094,22.462027,16.863113,11.2642,5.661383,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.23816854,0.3513962,0.46071947,0.57394713,0.6871748,1.5266213,2.3621633,3.2016098,4.037152,4.8765984,4.73604,4.5993857,4.462732,4.3260775,4.1894236,4.037152,3.8887846,3.736513,3.5881457,3.435874,3.8380275,4.2362766,4.6384296,5.036679,5.4388323,4.985922,4.5369153,4.087909,3.638903,3.1859922,3.4007344,3.611572,3.8263142,4.037152,4.251894,3.7638438,3.2757936,2.787743,2.2996929,1.8116426,1.7491722,1.6867018,1.6242313,1.5617609,1.4992905,3.1000953,4.7009,6.3017054,7.898606,9.499411,9.80005,10.100689,10.401327,10.698062,10.998701,12.400381,13.798158,15.199838,16.601519,17.999294,17.163752,16.324306,15.488764,14.649317,13.813775,13.513136,13.212498,12.911859,12.611219,12.31058,11.139259,9.964035,8.78881,7.6135845,6.4383593,6.348558,6.262661,6.1767645,6.086963,6.001066,7.648724,9.300286,10.951848,12.599506,14.251068,19.350218,24.449368,29.548515,34.65157,39.75072,38.813663,37.876606,36.935646,35.99859,35.06153,39.78586,44.51409,49.23842,53.96274,58.68707,48.024147,37.361225,26.698303,16.039284,5.376362,6.8756523,8.374943,9.874233,11.373524,12.8767185,12.63855,12.400381,12.162213,11.924045,11.685876,12.525322,13.360865,14.200311,15.035853,15.875299,21.12672,26.374237,31.625658,36.873177,42.124596,43.08898,44.049465,45.013855,45.974335,46.938725,45.56047,44.18612,42.81177,41.43742,40.063072,41.61312,43.163166,44.713215,46.263264,47.81331,48.024147,48.23889,48.449726,48.660564,48.87531,48.52391,48.17642,47.825024,47.473625,47.126137,46.700554,46.274975,45.849396,45.423817,44.998238,45.349632,45.701027,46.04852,46.399918,46.751312,47.5361,48.324787,49.113476,49.898262,50.68695,47.63761,44.588272,41.538937,38.485695,35.436356,34.788223,34.13619,33.48806,32.83602,32.187893,32.613472,33.03905,33.460728,33.886307,34.311886,31.563189,28.81449,26.061886,23.313187,20.560583,18.58886,16.613232,14.637604,12.661977,10.686349,11.974802,13.263254,14.551707,15.836256,17.124708,17.86264,18.600573,19.338505,20.076437,20.81437,20.388788,19.96321,19.537628,19.11205,18.68647,17.437061,16.187653,14.938243,13.688834,12.439425,12.013845,11.588266,11.162686,10.737106,10.311526,11.924045,13.536563,15.14908,16.761599,18.374117,18.68647,18.998821,19.311174,19.623526,19.935879,18.448301,16.960724,15.473146,13.989473,12.501896,12.0606985,11.623405,11.186112,10.748819,10.311526,10.826907,11.338385,11.849861,12.361338,12.8767185,11.514082,10.151445,8.78881,7.426173,6.0635366,6.375889,6.688241,7.000593,7.3129454,7.6252975,7.898606,8.175818,8.449126,8.726339,8.999647,10.4637985,11.924045,13.388195,14.848442,16.312593,16.476578,16.636658,16.800642,16.960724,17.124708,16.749886,16.375063,16.00024,15.625418,15.250595,15.875299,16.500004,17.124708,17.749413,18.374117,19.36193,20.349745,21.337559,22.325373,23.313187,22.62601,21.938837,21.251661,20.564487,19.873407,19.276033,18.674755,18.073479,17.476105,16.874826,16.125181,15.375536,14.625891,13.8762455,13.1266,12.123169,11.123642,10.124115,9.124588,8.125061,8.437413,8.749765,9.062118,9.37447,9.686822,1.5110037,1.5266213,1.5383345,1.5500476,1.5617609,1.5734742,1.5734742,1.5734742,1.5734742,1.5734742,1.5734742,1.5734742,1.5695697,1.5656652,1.5656652,1.5617609,1.5188124,1.475864,1.43682,1.3938715,1.3509232,1.3938715,1.43682,1.475864,1.5188124,1.5617609,1.6281357,1.698415,1.7647898,1.8311646,1.901444,1.7530766,1.6086137,1.4641509,1.319688,1.175225,4.5993857,8.019642,11.443803,14.864059,18.28822,15.293544,12.302772,9.308095,6.3173227,3.3265507,3.2679846,3.2094188,3.1508527,3.096191,3.0376248,2.639376,2.2372224,1.8389735,1.43682,1.038571,0.97610056,0.91753453,0.8589685,0.79649806,0.737932,0.75745404,0.77697605,0.79649806,0.8160201,0.8394465,0.6910792,0.5466163,0.40215343,0.25769055,0.113227665,0.09761006,0.08199245,0.06637484,0.05075723,0.039044023,0.031235218,0.027330816,0.023426414,0.015617609,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.14446288,0.20302892,0.26159495,0.31625658,0.37482262,1.5969005,2.8189783,4.041056,5.263134,6.4891167,6.114294,5.735567,5.3607445,4.985922,4.6110992,4.4314966,4.2479897,4.0644827,3.8809757,3.7013733,3.7716527,3.8458362,3.9161155,3.9902992,4.0605783,4.415879,4.7672753,5.1186714,5.473972,5.825368,5.6848097,5.5442514,5.4036927,5.263134,5.12648,4.970304,4.814128,4.661856,4.50568,4.349504,4.4393053,4.5252023,4.6110992,4.7009,4.786797,4.4978714,4.2089458,3.9161155,3.6271896,3.338264,3.736513,4.1308575,4.5291066,4.927356,5.3256044,5.481781,5.6418614,5.7980375,5.9542136,6.114294,6.649197,7.1880045,7.726812,8.261715,8.800523,8.566258,8.32809,8.093826,7.859562,7.6252975,7.6643414,7.699481,7.7385254,7.773665,7.812709,7.6916723,7.5667315,7.445695,7.320754,7.1997175,7.918128,8.636538,9.351044,10.069453,10.787864,11.861574,12.93138,14.005091,15.078801,16.148607,16.88654,17.620567,18.354595,19.088623,19.826555,19.584482,19.346313,19.10424,18.866072,18.623999,17.1169,15.605896,14.0948925,12.583888,11.076789,10.670732,10.264673,9.858616,9.456462,9.050405,9.386183,9.718058,10.053836,10.389614,10.725393,10.944039,11.158782,11.377428,11.596075,11.810817,12.326198,12.837675,13.349152,13.860628,14.376009,13.919194,13.466284,13.009468,12.556558,12.099743,14.661031,17.226223,19.78751,22.348799,24.91399,25.917421,26.920853,27.92819,28.931622,29.938957,30.091228,30.2435,30.395771,30.548042,30.700315,30.672985,30.645653,30.618322,30.590992,30.563662,30.14589,29.732023,29.318157,28.90429,28.486519,28.361578,28.232733,28.103888,27.978947,27.850101,31.898966,35.943928,39.992794,44.041656,48.086617,46.212505,44.33839,42.46428,40.58626,38.712147,35.366077,32.023907,28.677835,25.331762,21.98569,22.430792,22.871988,23.313187,23.758287,24.199486,25.070168,25.94085,26.811531,27.678308,28.548988,25.991606,23.430319,20.86903,18.311647,15.750359,14.313539,12.8767185,11.435994,9.999174,8.562354,8.648251,8.734148,8.81614,8.902037,8.987934,8.55845,8.128965,7.6955767,7.266093,6.8366084,7.6370106,8.437413,9.237816,10.0382185,10.838621,10.61607,10.393518,10.170968,9.948417,9.725866,10.608261,11.490656,12.373051,13.2554455,14.13784,15.461433,16.78112,18.104713,19.428307,20.751898,20.423927,20.099863,19.775797,19.451733,19.123762,17.72989,16.33602,14.938243,13.544372,12.150499,12.353529,12.560462,12.763491,12.970425,13.173453,15.434102,17.690847,19.947592,22.204336,24.46108,21.485926,18.51077,15.535617,12.564366,9.589212,13.903577,18.217941,22.532305,26.84667,31.161034,27.10436,23.047686,18.991013,14.934339,10.87376,12.814248,14.750832,16.687416,18.623999,20.560583,21.111103,21.657719,22.204336,22.750952,23.301472,18.67085,14.040231,9.40961,4.7789884,0.14836729,0.13665408,0.12103647,0.10541886,0.08980125,0.07418364,0.08199245,0.08980125,0.09761006,0.10541886,0.113227665,0.30454338,0.4958591,0.6910792,0.8823949,1.0737107,1.7530766,2.4285383,3.1079042,3.7833657,4.462732,4.31046,4.1581883,4.0059166,3.853645,3.7013733,3.7052777,3.7091823,3.7130866,3.7208953,3.7247996,4.11524,4.50568,4.8961205,5.2865605,5.6730967,5.2318993,4.786797,4.3416953,3.8965936,3.4514916,3.8106966,4.169902,4.5291066,4.8883114,5.251421,5.0483923,4.8492675,4.650143,4.4510183,4.251894,4.154284,4.056674,3.959064,3.8614538,3.7638438,5.337318,6.910792,8.488171,10.061645,11.639023,11.799104,11.959184,12.119265,12.2793455,12.439425,13.274967,14.114414,14.949956,15.789403,16.624945,15.890917,15.160794,14.426766,13.696643,12.962616,12.603411,12.24811,11.888905,11.533605,11.174399,10.569217,9.96013,9.351044,8.745861,8.136774,7.7385254,7.336372,6.9381227,6.5359693,6.13772,8.94889,11.763964,14.575133,17.386303,20.201378,24.49622,28.794966,33.09371,37.388557,41.6873,39.746815,37.806328,35.86584,33.929256,31.988768,36.25628,40.527695,44.79911,49.066624,53.33804,43.838627,34.33922,24.835903,15.336493,5.8370814,7.5667315,9.296382,11.0260315,12.755682,14.489237,13.716166,12.943093,12.170022,11.39695,10.6238785,12.228588,13.829392,15.434102,17.034906,18.635712,22.321468,26.003319,29.685171,33.367023,37.048874,37.724335,38.399796,39.075256,39.75072,40.42618,39.090874,37.759476,36.428074,35.096672,33.761368,35.2099,36.658432,38.106964,39.551594,41.00013,41.351524,41.699017,42.05041,42.40181,42.749302,42.885956,43.026512,43.163166,43.29982,43.436474,42.905476,42.370575,41.839573,41.308575,40.773674,40.773674,40.773674,40.773674,40.773674,40.773674,41.61312,42.44866,43.28811,44.12365,44.963097,42.417427,39.871758,37.326084,34.78432,32.23865,32.094185,31.953629,31.809166,31.668606,31.524143,31.965342,32.40654,32.84383,33.28503,33.726227,30.895535,28.068748,25.24196,22.415173,19.588387,17.874353,16.164225,14.450192,12.73616,11.0260315,12.056794,13.091461,14.122223,15.152986,16.187653,16.792833,17.398016,18.003199,18.608381,19.213564,19.13157,19.045673,18.963682,18.88169,18.799696,17.554192,16.30869,15.063184,13.821584,12.576079,12.091934,11.611692,11.127546,10.6434,10.163159,11.314958,12.466757,13.618555,14.774258,15.926057,16.324306,16.71865,17.1169,17.515148,17.913397,16.988054,16.062712,15.137367,14.212025,13.286681,12.490183,11.693685,10.893282,10.096785,9.300286,9.882042,10.4637985,11.0494585,11.631214,12.212971,11.217348,10.221725,9.226103,8.234385,7.238762,7.8634663,8.492075,9.120684,9.749292,10.373997,10.557504,10.741011,10.920613,11.10412,11.287627,12.70102,14.114414,15.523903,16.937298,18.35069,18.401447,18.448301,18.499058,18.549814,18.600573,18.256985,17.913397,17.573715,17.230127,16.88654,17.26917,17.651802,18.034433,18.417065,18.799696,19.803127,20.80656,21.806087,22.809519,23.81295,23.05159,22.294136,21.532778,20.77142,20.013966,19.393166,18.77627,18.159374,17.542479,16.925583,16.55076,16.175938,15.801116,15.426293,15.051471,13.7474,12.44333,11.143164,9.839094,8.538928,8.683391,8.827853,8.972317,9.116779,9.261242,1.5266213,1.5383345,1.5500476,1.5617609,1.5734742,1.5890918,1.6008049,1.6125181,1.6242313,1.6359446,1.6515622,1.6437533,1.639849,1.6359446,1.6281357,1.6242313,1.6008049,1.5812829,1.5578566,1.53443,1.5110037,1.53443,1.5578566,1.5812829,1.6008049,1.6242313,1.698415,1.7686942,1.8428779,1.9131571,1.9873407,1.8584955,1.7335546,1.6047094,1.475864,1.3509232,4.607195,7.8634663,11.123642,14.379913,17.636185,14.7156925,11.791295,8.870802,5.9464045,3.0259118,2.97125,2.920493,2.8658314,2.815074,2.7643168,2.4129205,2.0615244,1.7140326,1.3626363,1.0112402,0.95657855,0.8980125,0.8394465,0.78088045,0.7262188,0.7145056,0.7066968,0.6949836,0.6832704,0.6754616,0.57394713,0.46852827,0.3670138,0.26549935,0.1639849,0.14446288,0.12884527,0.10932326,0.093705654,0.07418364,0.06637484,0.05466163,0.046852827,0.03513962,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.27721256,0.37872702,0.48414588,0.58566034,0.6871748,1.8467822,3.0024853,4.1581883,5.3177958,6.473499,6.0752497,5.6730967,5.2748475,4.8765984,4.474445,4.31046,4.1464753,3.978586,3.814601,3.6506162,3.7833657,3.9161155,4.0488653,4.181615,4.3143644,4.579864,4.8492675,5.114767,5.3841705,5.64967,5.4583545,5.263134,5.0718184,4.8805027,4.689187,4.5291066,4.369026,4.2089458,4.0488653,3.8887846,3.998108,4.1113358,4.224563,4.337791,4.4510183,4.181615,3.9161155,3.6467118,3.3812122,3.1118085,3.4593005,3.802888,4.1464753,4.493967,4.8375545,5.001539,5.169429,5.3334136,5.4973984,5.661383,6.1611466,6.66091,7.1606736,7.6643414,8.164105,8.0040245,7.8478484,7.6916723,7.531592,7.375416,7.336372,7.3012323,7.262188,7.223144,7.1880045,7.2192397,7.2465706,7.277806,7.309041,7.336372,8.335898,9.331521,10.331048,11.326671,12.326198,13.157836,13.989473,14.821111,15.656653,16.48829,17.08176,17.679134,18.272602,18.866072,19.463446,19.194042,18.928543,18.659138,18.393639,18.124235,16.706938,15.285735,13.864532,12.44333,11.0260315,10.8542385,10.67854,10.506746,10.334952,10.163159,10.455989,10.752724,11.0494585,11.342289,11.639023,11.885,12.130978,12.380859,12.626837,12.8767185,13.462379,14.051944,14.637604,15.223265,15.812829,15.441911,15.067088,14.69617,14.321347,13.950429,16.062712,18.174992,20.287273,22.399555,24.511837,25.65973,26.807627,27.95552,29.103415,30.251308,29.931149,29.610987,29.290825,28.970665,28.650503,28.443571,28.240541,28.033607,27.83058,27.623646,27.568985,27.514322,27.459661,27.404999,27.350338,27.30739,27.26444,27.221493,27.178545,27.135595,31.383585,35.62767,39.871758,44.11584,48.36383,46.360874,44.36182,42.362766,40.363712,38.360752,35.35827,32.35578,29.353296,26.350811,23.348326,24.047213,24.746101,25.441086,26.139973,26.838861,26.702208,26.569458,26.432804,26.296148,26.163399,23.879324,21.599154,19.315079,17.031002,14.750832,13.360865,11.974802,10.588739,9.198771,7.812709,8.644346,9.475985,10.311526,11.143164,11.974802,11.178304,10.381805,9.581403,8.784905,7.988407,8.574067,9.163632,9.749292,10.338858,10.924518,10.467703,10.010887,9.554072,9.093353,8.636538,9.288573,9.940608,10.596548,11.248583,11.900618,13.32182,14.739119,16.16032,17.581524,18.998821,19.123762,19.248703,19.373644,19.498585,19.623526,18.3585,17.093473,15.828446,14.56342,13.298394,13.4858055,13.6693125,13.856724,14.040231,14.223738,16.164225,18.104713,20.0452,21.98569,23.926178,21.111103,18.299932,15.488764,12.67369,9.86252,13.766922,17.671324,21.575727,25.484034,29.388435,26.210253,23.032068,19.853886,16.675701,13.501423,14.661031,15.824542,16.988054,18.151566,19.311174,19.158901,19.002726,18.84655,18.694279,18.538101,14.875772,11.217348,7.558923,3.8965936,0.23816854,0.20693332,0.1756981,0.14836729,0.11713207,0.08589685,0.08980125,0.093705654,0.093705654,0.09761006,0.10151446,0.3709182,0.6442264,0.91753453,1.1908426,1.4641509,1.979532,2.4988174,3.0141985,3.533484,4.0488653,3.8809757,3.7130866,3.5491016,3.3812122,3.213323,3.3734035,3.533484,3.6935644,3.853645,4.0137253,4.3924527,4.7711797,5.153811,5.532538,5.911265,5.473972,5.0327744,4.591577,4.154284,3.7130866,4.220659,4.728231,5.2358036,5.743376,6.250948,6.336845,6.426646,6.5125427,6.5984397,6.688241,6.5554914,6.422742,6.289992,6.1572423,6.0244927,7.57454,9.124588,10.674636,12.224684,13.774731,13.794253,13.813775,13.833297,13.856724,13.8762455,14.149553,14.426766,14.700074,14.973383,15.250595,14.621986,13.993378,13.368673,12.740065,12.111456,11.697589,11.283723,10.865952,10.452085,10.0382185,9.999174,9.956225,9.917182,9.878138,9.839094,9.124588,8.413987,7.699481,6.98888,6.2743745,10.249056,14.223738,18.19842,22.177006,26.151686,29.646126,33.140568,36.635006,40.129448,43.623886,40.683872,37.739952,34.796032,31.856018,28.912098,32.7267,36.5413,40.355904,44.174408,47.98901,39.649204,31.313307,22.973503,14.637604,6.3017054,8.261715,10.221725,12.181735,14.141745,16.101755,14.79378,13.4858055,12.177831,10.869856,9.561881,11.931853,14.297921,16.663988,19.03396,21.400028,23.516214,25.628496,27.744682,29.860868,31.97315,32.36359,32.750126,33.13666,33.523197,33.91364,32.62128,31.332829,30.04047,28.752018,27.463566,28.80668,30.153698,31.496813,32.84383,34.186947,34.674995,35.163048,35.651096,36.13915,36.623295,37.251904,37.876606,38.501312,39.126015,39.75072,39.110397,38.470074,37.829754,37.18943,36.54911,36.20162,35.85022,35.498825,35.151333,34.79994,35.686237,36.57644,37.462738,38.349037,39.239243,37.19724,35.15914,33.11714,31.079042,29.037039,29.404053,29.767162,30.134176,30.497286,30.8643,31.317211,31.774025,32.226936,32.68375,33.13666,30.231787,27.326912,24.422035,21.51716,18.612286,17.163752,15.711315,14.262781,12.814248,11.361811,12.138786,12.915763,13.696643,14.473619,15.250595,15.723028,16.195461,16.667892,17.140326,17.612759,17.874353,18.132044,18.393639,18.651329,18.912924,17.671324,16.43363,15.192029,13.954333,12.712734,12.173926,11.631214,11.092407,10.553599,10.010887,10.705871,11.39695,12.091934,12.783013,13.4740925,13.958238,14.438479,14.922626,15.406772,15.8870125,15.523903,15.160794,14.801589,14.438479,14.07537,12.915763,11.760059,10.604357,9.444749,8.289046,8.941081,9.593117,10.2451515,10.897186,11.549222,10.920613,10.295909,9.6673,9.0386915,8.413987,9.354948,10.295909,11.240774,12.181735,13.1266,13.216402,13.306203,13.396004,13.4858055,13.575606,14.938243,16.300879,17.663515,19.026152,20.388788,20.326319,20.263847,20.201378,20.138906,20.076437,19.764084,19.455637,19.143284,18.834837,18.526388,18.666946,18.8036,18.94416,19.084719,19.225277,20.244326,21.25947,22.278519,23.293663,24.312714,23.481075,22.645533,21.813896,20.982258,20.15062,19.514202,18.88169,18.245272,17.608854,16.976341,16.976341,16.976341,16.976341,16.976341,16.976341,15.371632,13.763018,12.158309,10.553599,8.94889,8.929368,8.905942,8.882515,8.859089,8.835662,1.5383345,1.5500476,1.5617609,1.5734742,1.5890918,1.6008049,1.6242313,1.6515622,1.6749885,1.698415,1.7257458,1.717937,1.7101282,1.7023194,1.6945106,1.6867018,1.6867018,1.6827974,1.678893,1.678893,1.6749885,1.678893,1.678893,1.6827974,1.6867018,1.6867018,1.7647898,1.8428779,1.9209659,1.999054,2.0732377,1.9639144,1.8545911,1.7452679,1.6359446,1.5266213,4.618908,7.7111945,10.803481,13.895767,16.988054,14.133936,11.283723,8.429605,5.579391,2.7252727,2.67842,2.631567,2.5808098,2.533957,2.4871042,2.1864653,1.8858263,1.5890918,1.2884527,0.9878138,0.93315214,0.8784905,0.8238289,0.76916724,0.7106012,0.6715572,0.63251317,0.59346914,0.5544251,0.5114767,0.45291066,0.39434463,0.3318742,0.27330816,0.21083772,0.19131571,0.1717937,0.15227169,0.13274968,0.113227665,0.09761006,0.08199245,0.06637484,0.05075723,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10541886,0.15617609,0.21083772,0.26159495,0.40996224,0.5583295,0.7066968,0.8511597,0.999527,2.0927596,3.1859922,4.279225,5.368553,6.461786,6.036206,5.610626,5.1889505,4.7633705,4.337791,4.1894236,4.041056,3.8965936,3.7482262,3.5998588,3.7911747,3.9863946,4.1777105,4.369026,4.564246,4.743849,4.927356,5.1108627,5.2943697,5.473972,5.2318993,4.985922,4.7399445,4.493967,4.251894,4.084005,3.9200199,3.7560349,3.5881457,3.4241607,3.5608149,3.7013733,3.8380275,3.9746814,4.1113358,3.8692627,3.6232853,3.377308,3.1313305,2.8892577,3.1781836,3.4710135,3.7638438,4.056674,4.349504,4.521298,4.6930914,4.8687897,5.040583,5.212377,5.6730967,6.13772,6.5984397,7.0630636,7.523783,7.445695,7.363703,7.2856145,7.2036223,7.125534,7.012306,6.899079,6.785851,6.676528,6.5633,6.746807,6.9264097,7.1099167,7.2934237,7.47693,8.75367,10.03041,11.307149,12.583888,13.860628,14.454097,15.047566,15.641035,16.2306,16.82407,17.280884,17.733795,18.19061,18.64352,19.100336,18.8036,18.51077,18.214037,17.921206,17.624472,16.296974,14.965574,13.634172,12.306676,10.975275,11.033841,11.096312,11.154878,11.213444,11.275913,11.5297,11.783486,12.041177,12.294963,12.548749,12.825961,13.103174,13.384291,13.661504,13.938716,14.59856,15.262308,15.926057,16.585901,17.24965,16.960724,16.671797,16.378967,16.090042,15.801116,17.464392,19.123762,20.787037,22.450314,24.113588,25.40204,26.694399,27.982851,29.271303,30.563662,29.771067,28.978474,28.18588,27.393286,26.600693,26.218061,25.83543,25.452799,25.070168,24.687536,24.992079,25.296621,25.601166,25.905708,26.214157,26.2532,26.296148,26.339098,26.382046,26.424995,30.868204,35.311413,39.75072,44.193928,48.63714,46.513145,44.38915,42.26125,40.137257,38.01326,35.354362,32.69156,30.032661,27.373764,24.710962,25.663635,26.61631,27.568985,28.521658,29.474333,28.334248,27.194162,26.054077,24.91399,23.773905,21.770947,19.764084,17.761126,15.754263,13.751305,12.412095,11.076789,9.737579,8.398369,7.0630636,8.644346,10.221725,11.803008,13.384291,14.96167,13.798158,12.630741,11.46723,10.303718,9.136301,9.511124,9.885946,10.260769,10.6355915,11.014318,10.319335,9.628256,8.933272,8.242193,7.551114,7.9727893,8.3944645,8.81614,9.24172,9.663396,11.178304,12.697116,14.215929,15.730837,17.24965,17.823597,18.401447,18.975395,19.549341,20.12329,18.991013,17.854832,16.71865,15.586374,14.450192,14.614178,14.778163,14.946052,15.110037,15.274021,16.898252,18.51858,20.14281,21.763138,23.38737,20.73628,18.089096,15.438006,12.786918,10.135828,13.634172,17.128613,20.623053,24.117493,27.611933,25.316145,23.01645,20.720663,18.420969,16.125181,16.511717,16.898252,17.288692,17.675228,18.061766,17.206701,16.347733,15.488764,14.633699,13.774731,11.084598,8.3944645,5.704332,3.0141985,0.3240654,0.28111696,0.23426414,0.19131571,0.14446288,0.10151446,0.09761006,0.093705654,0.093705654,0.08980125,0.08589685,0.44119745,0.79259366,1.1439898,1.4992905,1.8506867,2.2059872,2.5651922,2.9243972,3.279698,3.638903,3.455396,3.2718892,3.0883822,2.9087796,2.7252727,3.0415294,3.3538816,3.6701381,3.9863946,4.298747,4.6696653,5.040583,5.4115014,5.7785153,6.1494336,5.716045,5.278752,4.845363,4.40807,3.9746814,4.630621,5.2865605,5.938596,6.5945354,7.250475,7.6252975,8.00012,8.374943,8.749765,9.124588,8.956698,8.78881,8.62092,8.453031,8.289046,9.811763,11.338385,12.861101,14.387722,15.914344,15.793307,15.672271,15.551234,15.434102,15.313066,15.024139,14.739119,14.450192,14.161267,13.8762455,13.353056,12.829865,12.306676,11.783486,11.2642,10.791768,10.319335,9.846903,9.370565,8.898132,9.4291315,9.956225,10.48332,11.010414,11.537509,10.510651,9.487698,8.460839,7.437886,6.4110284,11.549222,16.687416,21.82561,26.963802,32.09809,34.79213,37.486168,40.1763,42.87034,45.564373,41.617023,37.673576,33.726227,29.78278,25.839334,29.19712,32.55881,35.916595,39.278286,42.636074,35.463684,28.287394,21.111103,13.938716,6.7624245,8.952794,11.143164,13.333533,15.523903,17.714273,15.871395,14.028518,12.185639,10.342762,8.499884,11.631214,14.766449,17.89778,21.02911,24.164345,24.710962,25.257578,25.804195,26.350811,26.90133,26.998941,27.100456,27.201971,27.29958,27.401094,26.151686,24.906181,23.656773,22.411268,21.16186,22.40346,23.648964,24.890564,26.132164,27.373764,27.998468,28.623173,29.251781,29.876486,30.50119,31.613945,32.7267,33.839455,34.948303,36.061058,35.31532,34.565674,33.81993,33.074192,32.324547,31.625658,30.926771,30.223978,29.52509,28.826202,29.763258,30.700315,31.637371,32.57443,33.511486,31.977055,30.442625,28.908194,27.373764,25.839334,26.710016,27.580698,28.455284,29.325966,30.200552,30.669079,31.141512,31.61004,32.078568,32.551003,29.568039,26.585075,23.602112,20.619148,17.636185,16.449247,15.262308,14.07537,12.888432,11.701493,12.220779,12.743969,13.2671585,13.790349,14.313539,14.653222,14.992905,15.332587,15.672271,16.011953,16.613232,17.218414,17.819693,18.420969,19.026152,17.788456,16.554665,15.320874,14.0831785,12.849388,12.252014,11.654641,11.057267,10.459893,9.86252,10.096785,10.327144,10.561408,10.791768,11.0260315,11.592171,12.158309,12.728352,13.29449,13.860628,14.063657,14.262781,14.461906,14.661031,14.864059,13.345247,11.826434,10.311526,8.792714,7.2739015,7.996216,8.718531,9.440845,10.163159,10.889378,10.627783,10.366188,10.108498,9.846903,9.589212,10.84643,12.103647,13.360865,14.618082,15.875299,15.871395,15.871395,15.867491,15.863586,15.863586,17.175465,18.487345,19.799223,21.111103,22.426888,22.251188,22.07549,21.899792,21.724094,21.548395,21.271183,20.99397,20.716759,20.439547,20.162333,20.06082,19.959305,19.853886,19.75237,19.650856,20.68162,21.716286,22.747047,23.781713,24.812477,23.906654,23.000834,22.098917,21.193096,20.287273,19.635239,18.983204,18.33117,17.679134,17.023193,17.40192,17.776743,18.151566,18.526388,18.90121,16.991959,15.086611,13.177358,11.272009,9.362757,9.171441,8.98403,8.792714,8.601398,8.413987,1.5500476,1.5617609,1.5734742,1.5890918,1.6008049,1.6125181,1.6515622,1.6867018,1.7257458,1.7608855,1.7999294,1.7882162,1.7804074,1.7686942,1.7608855,1.7491722,1.7686942,1.7843118,1.8038338,1.8194515,1.8389735,1.8194515,1.8038338,1.7843118,1.7686942,1.7491722,1.8311646,1.9131571,1.999054,2.0810463,2.1630387,2.069333,1.9756275,1.8858263,1.7921207,1.698415,4.6267166,7.5550184,10.48332,13.411622,16.33602,13.556085,10.772245,7.988407,5.2084727,2.4246337,2.3816853,2.338737,2.2957885,2.2567444,2.2137961,1.9639144,1.7140326,1.4641509,1.2142692,0.96438736,0.9097257,0.8589685,0.80430686,0.75354964,0.698888,0.62860876,0.5583295,0.48805028,0.42167544,0.3513962,0.3318742,0.31625658,0.29673457,0.28111696,0.26159495,0.23816854,0.21864653,0.19522011,0.1717937,0.14836729,0.12884527,0.10932326,0.08980125,0.07027924,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07027924,0.14055848,0.21083772,0.28111696,0.3513962,0.5427119,0.7340276,0.92924774,1.1205635,1.3118792,2.338737,3.3655949,4.396357,5.423215,6.4500723,6.001066,5.548156,5.099149,4.650143,4.2011366,4.068387,3.9395418,3.8106966,3.6818514,3.5491016,3.802888,4.056674,4.3065557,4.560342,4.814128,4.911738,5.009348,5.1030536,5.2006636,5.298274,5.001539,4.704805,4.40807,4.1113358,3.8106966,3.6428072,3.4710135,3.3031244,3.1313305,2.9634414,3.1235218,3.2875066,3.4514916,3.611572,3.775557,3.5530062,3.330455,3.1079042,2.8853533,2.6628022,2.900971,3.1430438,3.3812122,3.6232853,3.8614538,4.041056,4.220659,4.4041657,4.5837684,4.7633705,5.1889505,5.610626,6.036206,6.461786,6.8873653,6.883461,6.883461,6.8795567,6.8756523,6.8756523,6.688241,6.5008297,6.3134184,6.126007,5.938596,6.2743745,6.606249,6.942027,7.277806,7.6135845,9.171441,10.729298,12.28325,13.841106,15.398962,15.754263,16.10566,16.457056,16.808453,17.163752,17.476105,17.79236,18.108618,18.420969,18.737226,18.41316,18.093,17.768934,17.448774,17.124708,15.883108,14.645412,13.403813,12.166118,10.924518,11.217348,11.510178,11.803008,12.095839,12.388668,12.603411,12.818152,13.032895,13.247637,13.462379,13.770826,14.079274,14.383818,14.6922655,15.000713,15.738646,16.476578,17.210606,17.948538,18.68647,18.479536,18.272602,18.06567,17.858736,17.651802,18.862167,20.076437,21.2868,22.50107,23.711435,25.14435,26.577267,28.010181,29.443098,30.876013,29.610987,28.34596,27.080935,25.815908,24.55088,23.988647,23.430319,22.868084,22.309755,21.751425,22.415173,23.078922,23.746574,24.410322,25.074072,25.202917,25.331762,25.456703,25.585548,25.714394,30.352823,34.991253,39.633587,44.27202,48.914352,46.66151,44.412575,42.16364,39.9108,37.661865,35.346554,33.02734,30.708124,28.392813,26.073599,27.283962,28.490423,29.696884,30.903343,32.11371,29.966288,27.822771,25.679255,23.531832,21.388315,19.658665,17.93292,16.20327,14.477524,12.751778,11.4633255,10.174872,8.886419,7.601871,6.3134184,8.640442,10.967466,13.29449,15.621513,17.948538,16.41801,14.883581,13.353056,11.818625,10.2881,10.44818,10.612165,10.77615,10.936231,11.100216,10.170968,9.245625,8.316377,7.3910336,6.461786,6.6531014,6.8483214,7.039637,7.230953,7.426173,9.0386915,10.655114,12.271536,13.884054,15.500477,16.52343,17.550287,18.573242,19.6001,20.626957,19.619621,18.61619,17.608854,16.605423,15.598087,15.746454,15.890917,16.03538,16.179844,16.324306,17.628376,18.936352,20.240421,21.54449,22.848562,20.361458,17.874353,15.387249,12.900145,10.413041,13.497519,16.581997,19.666473,22.750952,25.839334,24.41813,23.000834,21.583536,20.166237,18.74894,18.362404,17.975868,17.589333,17.198893,16.812357,15.250595,13.692739,12.130978,10.573121,9.01136,7.2934237,5.571582,3.853645,2.1318035,0.41386664,0.3513962,0.29283017,0.23426414,0.1717937,0.113227665,0.10541886,0.09761006,0.08980125,0.08199245,0.07418364,0.5075723,0.94096094,1.3743496,1.8038338,2.2372224,2.436347,2.631567,2.8306916,3.0259118,3.2250361,3.0259118,2.8306916,2.631567,2.436347,2.2372224,2.7057507,3.1781836,3.6467118,4.1191444,4.5876727,4.9468775,5.3060827,5.6691923,6.028397,6.387602,5.958118,5.5286336,5.099149,4.6657605,4.2362766,5.040583,5.840986,6.6452928,7.445695,8.250002,8.913751,9.573594,10.237343,10.901091,11.560935,11.361811,11.158782,10.955752,10.752724,10.549695,12.0489855,13.548276,15.051471,16.55076,18.05005,17.788456,17.530766,17.26917,17.01148,16.749886,15.8987255,15.051471,14.200311,13.349152,12.501896,12.084125,11.666354,11.248583,10.8308115,10.413041,9.882042,9.351044,8.823949,8.292951,7.7619514,8.859089,9.952321,11.0494585,12.142691,13.235924,11.900618,10.561408,9.226103,7.8868923,6.551587,12.849388,19.151093,25.448895,31.750599,38.0484,39.942036,41.831764,43.721497,45.61123,47.500957,42.55408,37.6033,32.65642,27.709543,22.762665,25.66754,28.572416,31.477291,34.382168,37.28704,31.274261,25.261482,19.248703,13.235924,7.223144,9.643873,12.064603,14.4853325,16.906061,19.326792,16.94901,14.571229,12.193448,9.815667,7.437886,11.334479,15.231073,19.13157,23.028164,26.924759,25.905708,24.88666,23.863707,22.844658,21.82561,21.638197,21.450787,21.263374,21.075964,20.888552,19.682093,18.475632,17.273075,16.066616,14.864059,16.004145,17.14423,18.284315,19.420496,20.560583,21.325846,22.087204,22.848562,23.613825,24.375183,25.975988,27.576794,29.173695,30.774498,32.375305,31.520239,30.665174,29.810112,28.955048,28.099983,27.049698,25.999414,24.949131,23.898846,22.848562,23.836376,24.82419,25.812004,26.799816,27.78763,26.756868,25.726107,24.69925,23.668486,22.637724,24.015978,25.398136,26.77639,28.158548,29.536802,30.020948,30.508999,30.993145,31.477291,31.961437,28.900385,25.843239,22.782187,19.721136,16.663988,15.738646,14.813302,13.887959,12.962616,12.037272,12.306676,12.572175,12.841579,13.107079,13.376482,13.583415,13.790349,13.997282,14.204215,14.411149,15.356014,16.300879,17.245745,18.19061,19.13938,17.905588,16.675701,15.445815,14.215929,12.986042,12.334006,11.678067,11.022127,10.366188,9.714153,9.483793,9.257338,9.030883,8.804427,8.574067,9.226103,9.878138,10.534078,11.186112,11.838148,12.599506,13.360865,14.126127,14.8874855,15.648844,13.770826,11.896713,10.018696,8.140678,6.262661,7.055255,7.8478484,8.640442,9.433036,10.22563,10.331048,10.4403715,10.545791,10.655114,10.764437,12.334006,13.907481,15.480955,17.050524,18.623999,18.530293,18.436588,18.338978,18.245272,18.151566,19.412687,20.67381,21.938837,23.199959,24.46108,24.17606,23.887133,23.598207,23.313187,23.02426,22.778282,22.53621,22.290232,22.044254,21.798277,21.45469,21.111103,20.76361,20.420023,20.076437,21.122816,22.169195,23.21948,24.26586,25.31224,24.33614,23.356134,22.380033,21.403933,20.423927,19.756275,19.084719,18.41316,17.745508,17.073952,17.823597,18.573242,19.326792,20.076437,20.826082,18.61619,16.406298,14.196406,11.986515,9.776623,9.4174185,9.058213,8.702912,8.343708,7.988407,1.5617609,1.5734742,1.5890918,1.6008049,1.6125181,1.6242313,1.6749885,1.7257458,1.7765031,1.8233559,1.8741131,1.8623998,1.8506867,1.8389735,1.8233559,1.8116426,1.8506867,1.8858263,1.9248703,1.9639144,1.999054,1.9639144,1.9248703,1.8858263,1.8506867,1.8116426,1.901444,1.9873407,2.0732377,2.1630387,2.2489357,2.174752,2.1005683,2.0263848,1.9482968,1.8741131,4.6384296,7.3988423,10.163159,12.923572,15.687888,12.974329,10.260769,7.551114,4.8375545,2.1239948,2.0888553,2.0498111,2.0107672,1.9756275,1.9365835,1.737459,1.5383345,1.33921,1.1361811,0.93705654,0.8862993,0.8394465,0.78868926,0.737932,0.6871748,0.58566034,0.48805028,0.38653582,0.28892577,0.18741131,0.21083772,0.23816854,0.26159495,0.28892577,0.31235218,0.28892577,0.26159495,0.23816854,0.21083772,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.6754616,0.9136301,1.1517987,1.3860629,1.6242313,2.5886188,3.5491016,4.513489,5.473972,6.4383593,5.9620223,5.4856853,5.0132523,4.5369153,4.0605783,3.951255,3.8380275,3.7247996,3.611572,3.4983444,3.8106966,4.123049,4.4393053,4.7516575,5.0640097,5.0757227,5.087436,5.099149,5.1108627,5.12648,4.775084,4.423688,4.0761957,3.7247996,3.3734035,3.2016098,3.0259118,2.8502135,2.6745155,2.4988174,2.6862288,2.87364,3.0610514,3.2484627,3.435874,3.2367494,3.0376248,2.8385005,2.639376,2.436347,2.6237583,2.8111696,2.998581,3.1859922,3.3734035,3.5608149,3.7482262,3.9356375,4.126953,4.3143644,4.7009,5.087436,5.473972,5.8644123,6.250948,6.3251314,6.3993154,6.473499,6.551587,6.6257706,6.364176,6.098676,5.8370814,5.575486,5.3138914,5.801942,6.2860875,6.774138,7.262188,7.7502384,9.589212,11.424281,13.263254,15.098324,16.937298,17.050524,17.163752,17.273075,17.386303,17.49953,17.675228,17.850927,18.026625,18.19842,18.374117,18.026625,17.675228,17.323833,16.976341,16.624945,15.473146,14.325252,13.173453,12.025558,10.87376,11.400854,11.924045,12.4511385,12.974329,13.501423,13.673217,13.848915,14.024612,14.200311,14.376009,14.711788,15.051471,15.387249,15.726933,16.062712,16.874826,17.686943,18.499058,19.311174,20.12329,19.998348,19.873407,19.748466,19.623526,19.498585,20.263847,21.025206,21.786564,22.551826,23.313187,24.88666,26.464039,28.037512,29.610987,31.188366,29.450907,27.713448,25.975988,24.23853,22.50107,21.763138,21.025206,20.287273,19.549341,18.81141,19.838268,20.861221,21.888079,22.911032,23.937891,24.148727,24.36347,24.574308,24.78905,24.999887,29.837442,34.674995,39.51255,44.350105,49.18766,46.81378,44.436,42.062126,39.688248,37.314373,35.338745,33.363117,31.38749,29.411861,27.436235,28.900385,30.360632,31.824783,33.288933,34.74918,31.598328,28.45138,25.300526,22.149673,18.998821,17.550287,16.101755,14.649317,13.200784,11.748346,10.510651,9.276859,8.039165,6.801469,5.563773,8.636538,11.713207,14.785972,17.86264,20.93931,19.037865,17.136421,15.238882,13.337439,11.435994,11.389141,11.338385,11.287627,11.23687,11.186112,10.0265045,8.862993,7.699481,6.5359693,5.376362,5.337318,5.298274,5.263134,5.22409,5.1889505,6.899079,8.6131115,10.323239,12.037272,13.751305,15.223265,16.69913,18.174992,19.650856,21.12672,20.24823,19.373644,18.499058,17.624472,16.749886,16.874826,16.999767,17.124708,17.24965,17.37459,18.362404,19.350218,20.338032,21.325846,22.31366,19.986635,17.663515,15.336493,13.013372,10.686349,13.360865,16.039284,18.7138,21.388315,24.062832,23.524023,22.98912,22.450314,21.911505,21.376602,20.21309,19.049578,17.886066,16.72646,15.562947,13.298394,11.037745,8.773191,6.5125427,4.251894,3.4983444,2.7486992,1.999054,1.2494087,0.4997635,0.42557985,0.3513962,0.27330816,0.19912452,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.57394713,1.0893283,1.6008049,2.1122816,2.6237583,2.6628022,2.7018464,2.736986,2.77603,2.8111696,2.6003318,2.3855898,2.174752,1.9639144,1.7491722,2.3738766,2.998581,3.6232853,4.251894,4.8765984,5.22409,5.575486,5.9268827,6.2743745,6.6257706,6.2001905,5.774611,5.349031,4.9234514,4.5017757,5.4505453,6.3993154,7.348085,8.300759,9.249529,10.198298,11.150972,12.099743,13.048512,14.001186,13.763018,13.524849,13.286681,13.048512,12.814248,14.286208,15.762072,17.237936,18.7138,20.18576,19.78751,19.389261,18.987108,18.58886,18.186707,16.773312,15.363823,13.950429,12.537036,11.123642,10.81129,10.498938,10.186585,9.874233,9.561881,8.976221,8.386656,7.800996,7.211431,6.6257706,8.289046,9.948417,11.611692,13.274967,14.938243,13.286681,11.639023,9.987461,8.335898,6.688241,14.149553,21.610867,29.076084,36.537395,43.99871,45.088036,46.173462,47.26279,48.348213,49.437542,43.487232,37.536922,31.586615,25.636305,19.685997,22.13796,24.586021,27.037985,29.486046,31.938011,27.088743,22.239475,17.386303,12.537036,7.687768,10.338858,12.986042,15.637131,18.28822,20.93931,18.026625,15.113941,12.201257,9.288573,6.375889,11.037745,15.699601,20.361458,25.023314,29.689075,27.100456,24.511837,21.923218,19.338505,16.749886,16.273548,15.801116,15.324779,14.848442,14.376009,13.212498,12.0489855,10.889378,9.725866,8.562354,9.600925,10.6355915,11.674163,12.712734,13.751305,14.649317,15.551234,16.449247,17.351164,18.249176,20.338032,22.426888,24.511837,26.600693,28.685644,27.72516,26.760773,25.80029,24.835903,23.87542,22.47374,21.075964,19.674282,18.276506,16.874826,17.913397,18.948065,19.986635,21.025206,22.063778,21.536682,21.013493,20.486399,19.96321,19.436115,21.325846,23.211672,25.101402,26.987228,28.873055,29.376722,29.876486,30.37625,30.876013,31.375776,28.236637,25.101402,21.962263,18.823124,15.687888,15.024139,14.364296,13.700547,13.036799,12.373051,12.388668,12.400381,12.412095,12.423808,12.439425,12.513609,12.587793,12.661977,12.73616,12.814248,14.098797,15.387249,16.675701,17.964155,19.248703,18.026625,16.800642,15.57466,14.348679,13.1266,12.412095,11.701493,10.986988,10.276386,9.561881,8.874706,8.187531,7.5003567,6.813182,6.126007,6.8639393,7.601871,8.335898,9.073831,9.811763,11.139259,12.4628525,13.786445,15.113941,16.437534,14.200311,11.963089,9.725866,7.4886436,5.251421,6.114294,6.9732623,7.8361354,8.699008,9.561881,10.0382185,10.510651,10.986988,11.4633255,11.935758,13.825488,15.711315,17.601046,19.486872,21.376602,21.189192,21.00178,20.81437,20.626957,20.435642,21.64991,22.86418,24.074545,25.288813,26.499178,26.10093,25.698776,25.300526,24.898373,24.500124,24.289286,24.074545,23.863707,23.648964,23.438128,22.848562,22.262901,21.673336,21.087677,20.498112,21.564014,22.62601,23.68801,24.750006,25.812004,24.761719,23.711435,22.66115,21.610867,20.560583,19.873407,19.186234,18.499058,17.811884,17.124708,18.249176,19.373644,20.498112,21.626484,22.750952,20.236517,17.725986,15.211552,12.70102,10.186585,9.663396,9.136301,8.6131115,8.086017,7.562827,1.5383345,1.5539521,1.5656652,1.5812829,1.5969005,1.6125181,1.6593709,1.7023194,1.7491722,1.7921207,1.8389735,1.8428779,1.8467822,1.8506867,1.8584955,1.8623998,1.8975395,1.9326792,1.9678187,2.0029583,2.0380979,2.0107672,1.9834363,1.9561055,1.9287747,1.901444,1.9717231,2.0380979,2.1083772,2.1786566,2.2489357,2.4012074,2.5534792,2.7057507,2.8619268,3.0141985,5.1577153,7.3012323,9.448653,11.592171,13.735687,11.377428,9.019169,6.657006,4.298747,1.9365835,1.8897307,1.8428779,1.796025,1.7491722,1.698415,1.5305257,1.358732,1.1908426,1.0190489,0.8511597,0.80430686,0.75354964,0.7066968,0.659844,0.61299115,0.5270943,0.44119745,0.359205,0.27330816,0.18741131,0.20302892,0.21864653,0.23426414,0.24597734,0.26159495,0.24207294,0.22255093,0.20302892,0.1835069,0.1639849,0.14055848,0.12103647,0.10151446,0.08199245,0.062470436,0.058566034,0.05075723,0.046852827,0.042948425,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14446288,0.21864653,0.28892577,0.3631094,0.61689556,0.8667773,1.1205635,1.3743496,1.6242313,2.4441557,3.260176,4.0761957,4.8961205,5.7121406,5.3334136,4.958591,4.579864,4.2011366,3.8263142,3.7443218,3.6662338,3.5842414,3.506153,3.4241607,3.6935644,3.959064,4.2284675,4.493967,4.7633705,4.7633705,4.7672753,4.7711797,4.7711797,4.775084,4.447114,4.1191444,3.7911747,3.4632049,3.1391394,3.0805733,3.0220075,2.9634414,2.9087796,2.8502135,2.900971,2.951728,2.998581,3.049338,3.1000953,3.0805733,3.0649557,3.049338,3.0298162,3.0141985,3.0883822,3.1664703,3.2445583,3.3226464,3.4007344,3.6076677,3.814601,4.0215344,4.2284675,4.4393053,4.6540475,4.872694,5.0913405,5.3060827,5.5247293,5.5871997,5.64967,5.7121406,5.774611,5.8370814,5.645766,5.45445,5.2592297,5.067914,4.8765984,5.290465,5.704332,6.1181984,6.5359693,6.949836,8.581876,10.213917,11.845957,13.481901,15.113941,15.531713,15.953387,16.371159,16.792833,17.210606,17.218414,17.226223,17.234032,17.24184,17.24965,16.792833,16.33602,15.879204,15.418485,14.96167,13.985569,13.013372,12.037272,11.061172,10.088976,10.686349,11.287627,11.888905,12.486279,13.087557,13.25935,13.431144,13.606842,13.778636,13.950429,14.379913,14.809398,15.238882,15.668366,16.101755,16.730364,17.358973,17.991486,18.620094,19.248703,19.268225,19.283842,19.303364,19.318983,19.338505,19.85779,20.377075,20.89636,21.415646,21.938837,23.035973,24.137014,25.238056,26.339098,27.436235,25.901804,24.367374,22.832945,21.298513,19.764084,19.604004,19.447828,19.29165,19.13157,18.975395,20.072533,21.169668,22.266806,23.363943,24.46108,24.98427,25.503555,26.02284,26.542126,27.061413,31.446056,35.8307,40.219246,44.60389,48.988537,47.73132,46.4741,45.21688,43.95576,42.698544,40.820526,38.938602,37.060585,35.178665,33.300648,34.038578,34.780415,35.51835,36.260185,36.998116,32.960964,28.919907,24.87885,20.8417,16.800642,15.637131,14.473619,13.314012,12.150499,10.986988,10.6434,10.295909,9.952321,9.608734,9.261242,11.584361,13.903577,16.222792,18.542006,20.861221,18.787983,16.710842,14.637604,12.564366,10.487225,10.569217,10.647305,10.729298,10.807385,10.889378,9.749292,8.609207,7.4691215,6.329036,5.1889505,5.263134,5.3412223,5.4193106,5.4973984,5.575486,7.094299,8.609207,10.128019,11.6468315,13.16174,14.746927,16.332115,17.917301,19.50249,21.087677,20.50592,19.924164,19.338505,18.756748,18.174992,18.276506,18.381926,18.48344,18.584955,18.68647,19.190138,19.693806,20.19357,20.697237,21.200905,20.021774,18.84655,17.66742,16.48829,15.313066,16.933393,18.557625,20.181856,21.802181,23.426414,22.481548,21.536682,20.591818,19.643047,18.698183,18.534197,18.370213,18.206228,18.038338,17.874353,15.344301,12.810344,10.276386,7.746334,5.212377,4.290938,3.3734035,2.4519646,1.53443,0.61299115,0.5192855,0.42557985,0.3357786,0.24207294,0.14836729,0.12884527,0.10932326,0.08980125,0.07027924,0.05075723,0.5349031,1.0190489,1.5031948,1.9912452,2.475391,2.5612879,2.6432803,2.7291772,2.815074,2.900971,2.6276627,2.3543546,2.0810463,1.8116426,1.5383345,2.1396124,2.7408905,3.3460727,3.9473507,4.548629,4.83365,5.114767,5.395884,5.6809053,5.9620223,5.6965227,5.4310236,5.169429,4.903929,4.6384296,5.434928,6.2314262,7.0318284,7.8283267,8.624825,9.343235,10.061645,10.77615,11.49456,12.212971,12.189544,12.166118,12.146595,12.123169,12.099743,13.177358,14.254972,15.332587,16.410202,17.487818,17.280884,17.077856,16.870922,16.667892,16.46096,15.324779,14.188598,13.048512,11.912332,10.77615,10.436467,10.100689,9.761005,9.425227,9.089449,8.531119,7.9727893,7.4144597,6.8561306,6.3017054,7.6135845,8.929368,10.2451515,11.560935,12.8767185,12.447234,12.021654,11.592171,11.166591,10.737106,17.234032,23.727053,30.223978,36.717,43.213924,43.061653,42.90938,42.753204,42.600933,42.44866,37.92346,33.394352,28.86915,24.340044,19.810938,21.895887,23.980839,26.06579,28.15074,30.235691,26.132164,22.028637,17.921206,13.817679,9.714153,11.639023,13.567798,15.4965725,17.421442,19.350218,16.652275,13.954333,11.256392,8.55845,5.8644123,11.088503,16.312593,21.536682,26.760773,31.988768,28.34596,24.707058,21.068155,17.429253,13.786445,13.638077,13.4858055,13.337439,13.189071,13.036799,11.900618,10.768341,9.63216,8.495979,7.363703,8.097731,8.831758,9.565785,10.303718,11.037745,11.760059,12.482374,13.204688,13.927003,14.649317,16.410202,18.171087,19.931974,21.688955,23.44984,22.684578,21.919313,21.15405,20.388788,19.623526,18.592764,17.558098,16.527334,15.4965725,14.461906,15.398962,16.33602,17.273075,18.214037,19.151093,19.041769,18.928543,18.81922,18.709896,18.600573,20.033487,21.470308,22.903223,24.340044,25.776863,25.979893,26.186827,26.389854,26.596788,26.799816,24.546976,22.294136,20.041296,17.788456,15.535617,15.043662,14.551707,14.059752,13.567798,13.075843,12.90405,12.73616,12.564366,12.396477,12.224684,12.185639,12.150499,12.111456,12.076316,12.037272,13.06413,14.090988,15.12175,16.148607,17.175465,16.222792,15.270117,14.317443,13.364769,12.412095,11.8537655,11.29934,10.741011,10.182681,9.6243515,8.85128,8.078208,7.309041,6.5359693,5.7628975,6.3407493,6.9225054,7.504261,8.082112,8.663869,9.796145,10.932326,12.068507,13.200784,14.336966,13.040704,11.744442,10.444276,9.148014,7.8517528,8.531119,9.2104845,9.889851,10.569217,11.248583,12.029464,12.810344,13.591225,14.3682,15.14908,16.359446,17.56981,18.780174,19.99054,21.200905,20.853413,20.50592,20.158428,19.810938,19.463446,20.34584,21.228235,22.11063,22.993025,23.87542,23.887133,23.898846,23.910559,23.926178,23.937891,23.789522,23.641155,23.496693,23.348326,23.199959,22.53621,21.868557,21.20481,20.54106,19.873407,20.93931,22.00521,23.071114,24.13311,25.199013,24.36347,23.531832,22.696291,21.860748,21.025206,20.19357,19.365835,18.534197,17.706465,16.874826,17.917301,18.959778,20.002253,21.044727,22.087204,19.818747,17.550287,15.285735,13.017277,10.748819,10.311526,9.874233,9.43694,8.999647,8.562354,1.5110037,1.5305257,1.5461433,1.5656652,1.5812829,1.6008049,1.639849,1.678893,1.7218413,1.7608855,1.7999294,1.8233559,1.8467822,1.8663043,1.8897307,1.9131571,1.9443923,1.9756275,2.0107672,2.0420024,2.0732377,2.05762,2.0380979,2.0224805,2.0068626,1.9873407,2.0380979,2.0927596,2.1435168,2.1981785,2.2489357,2.631567,3.0102942,3.3890212,3.7716527,4.1503797,5.677001,7.2036223,8.734148,10.260769,11.787391,9.780528,7.773665,5.7668023,3.7560349,1.7491722,1.6906061,1.6359446,1.5773785,1.5188124,1.4641509,1.3235924,1.183034,1.0424755,0.9019169,0.76135844,0.71841,0.6715572,0.62860876,0.58175594,0.5388075,0.46852827,0.39824903,0.3279698,0.25769055,0.18741131,0.19131571,0.19912452,0.20302892,0.20693332,0.21083772,0.19912452,0.1835069,0.1678893,0.15227169,0.13665408,0.12103647,0.10932326,0.093705654,0.078088045,0.062470436,0.06637484,0.06637484,0.07027924,0.07418364,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.113227665,0.1717937,0.23035973,0.28892577,0.5544251,0.8238289,1.0893283,1.358732,1.6242313,2.2957885,2.97125,3.6428072,4.3143644,4.985922,4.7087092,4.4275923,4.1464753,3.8692627,3.5881457,3.541293,3.49444,3.4436827,3.39683,3.349977,3.5725281,3.795079,4.01763,4.240181,4.462732,4.454923,4.447114,4.4393053,4.4314966,4.423688,4.1191444,3.814601,3.5100577,3.2055142,2.900971,2.959537,3.018103,3.0805733,3.1391394,3.2016098,3.1118085,3.0259118,2.9361105,2.8502135,2.7643168,2.9283018,3.0922866,3.2562714,3.4241607,3.5881457,3.5569105,3.521771,3.4905357,3.4593005,3.4241607,3.6506162,3.8809757,4.1074314,4.3338866,4.564246,4.6110992,4.657952,4.704805,4.7516575,4.7985106,4.8492675,4.900025,4.950782,5.001539,5.0483923,4.927356,4.806319,4.6813784,4.560342,4.4393053,4.7789884,5.1225758,5.466163,5.805846,6.1494336,7.578445,9.0035515,10.432563,11.861574,13.286681,14.016804,14.743023,15.469242,16.199366,16.925583,16.765503,16.605423,16.445343,16.285261,16.125181,15.559043,14.996809,14.430671,13.864532,13.298394,12.501896,11.701493,10.901091,10.100689,9.300286,9.975748,10.651209,11.326671,11.998228,12.67369,12.845484,13.013372,13.185166,13.353056,13.524849,14.048039,14.571229,15.0944195,15.613705,16.136894,16.585901,17.031002,17.48001,17.929016,18.374117,18.534197,18.694279,18.854359,19.014439,19.174519,19.451733,19.728945,20.006157,20.28337,20.560583,21.189192,21.813896,22.4386,23.063305,23.68801,22.356607,21.021301,19.689901,18.3585,17.023193,17.448774,17.87045,18.292124,18.7138,19.13938,20.306797,21.478117,22.649437,23.816854,24.988174,25.815908,26.64364,27.471375,28.299107,29.12684,33.058575,36.990307,40.92204,44.853775,48.78941,48.648853,48.508293,48.367737,48.227177,48.086617,46.302307,44.517994,42.733685,40.94937,39.161156,39.180676,39.196293,39.215816,39.231434,39.250957,34.319695,29.388435,24.46108,19.52982,14.59856,13.723974,12.849388,11.974802,11.100216,10.22563,10.772245,11.318862,11.869383,12.415999,12.962616,14.528281,16.093946,17.655706,19.221373,20.787037,18.538101,16.289165,14.036326,11.787391,9.538455,9.749292,9.956225,10.167064,10.377901,10.588739,9.468176,8.351517,7.2348576,6.1181984,5.001539,5.192855,5.3841705,5.579391,5.7707067,5.9620223,7.2856145,8.609207,9.928895,11.252487,12.576079,14.27059,15.965101,17.65961,19.354122,21.048632,20.759706,20.470781,20.181856,19.889025,19.6001,19.678188,19.76018,19.838268,19.92026,19.998348,20.01787,20.033487,20.053009,20.068628,20.08815,20.056915,20.025679,19.998348,19.967113,19.935879,20.50592,21.075964,21.646006,22.21605,22.78609,21.43517,20.084246,18.729418,17.378494,16.023666,16.85921,17.690847,18.522484,19.354122,20.18576,17.386303,14.582942,11.779582,8.976221,6.1767645,5.083532,3.9942036,2.9048753,1.815547,0.7262188,0.61689556,0.5036679,0.39434463,0.28502136,0.1756981,0.14836729,0.12103647,0.093705654,0.06637484,0.039044023,0.4958591,0.95267415,1.4094892,1.8663043,2.3231194,2.455869,2.5886188,2.7213683,2.854118,2.9868677,2.6549935,2.3231194,1.9912452,1.6593709,1.3235924,1.9053483,2.4831998,3.0649557,3.6467118,4.224563,4.4393053,4.6540475,4.8687897,5.083532,5.298274,5.196759,5.0913405,4.985922,4.8805027,4.775084,5.4193106,6.0635366,6.7116675,7.355894,8.00012,8.484266,8.968412,9.456462,9.940608,10.424754,10.61607,10.81129,11.002605,11.193921,11.389141,12.068507,12.747873,13.427239,14.106606,14.785972,14.778163,14.766449,14.75864,14.746927,14.739119,13.8762455,13.013372,12.150499,11.287627,10.424754,10.061645,9.698535,9.339331,8.976221,8.6131115,8.086017,7.558923,7.0318284,6.5008297,5.9737353,6.942027,7.910319,8.878611,9.846903,10.81129,11.607788,12.404286,13.196879,13.993378,14.785972,20.314606,25.843239,31.371872,36.896603,42.425236,41.031364,39.641396,38.247524,36.853653,35.463684,32.35578,29.251781,26.147781,23.043781,19.935879,21.657719,23.375656,25.097498,26.81934,28.537275,25.175587,21.8178,18.45611,15.098324,11.736633,12.943093,14.145649,15.35211,16.55857,17.761126,15.277926,12.798631,10.315431,7.832231,5.349031,11.139259,16.925583,22.711908,28.498232,34.28846,29.59537,24.902277,20.209187,15.516094,10.826907,10.998701,11.174399,11.350098,11.525795,11.701493,10.592644,9.483793,8.378847,7.269997,6.1611466,6.5945354,7.027924,7.461313,7.890797,8.324185,8.870802,9.413514,9.96013,10.506746,11.0494585,12.482374,13.91529,15.348206,16.78112,18.214037,17.643993,17.077856,16.511717,15.941674,15.375536,14.711788,14.044135,13.380386,12.716639,12.0489855,12.888432,13.723974,14.56342,15.398962,16.238409,16.542952,16.847496,17.152039,17.456583,17.761126,18.745035,19.728945,20.70895,21.69286,22.67677,22.583063,22.493261,22.40346,22.31366,22.223858,20.857317,19.490776,18.124235,16.75379,15.387249,15.063184,14.743023,14.418958,14.098797,13.774731,13.423335,13.0719385,12.716639,12.365242,12.013845,11.861574,11.713207,11.560935,11.412568,11.2642,12.029464,12.798631,13.563893,14.33306,15.098324,14.418958,13.739592,13.0602255,12.380859,11.701493,11.29934,10.893282,10.491129,10.088976,9.686822,8.831758,7.9727893,7.113821,6.2587566,5.3997884,5.8214636,6.2431393,6.6687193,7.0903945,7.5120697,8.456935,9.4018,10.346666,11.291532,12.236397,11.881096,11.521891,11.166591,10.807385,10.44818,10.947944,11.443803,11.943566,12.439425,12.939189,14.020708,15.1061325,16.191557,17.27698,18.362404,18.893402,19.428307,19.959305,20.494207,21.025206,20.517633,20.010061,19.50249,18.994917,18.487345,19.041769,19.59229,20.146715,20.697237,21.251661,21.673336,22.098917,22.524496,22.950077,23.375656,23.293663,23.211672,23.125774,23.043781,22.96179,22.219954,21.478117,20.73628,19.994444,19.248703,20.31851,21.38441,22.454218,23.520119,24.586021,23.969126,23.348326,22.727526,22.106726,21.485926,20.51373,19.541533,18.569338,17.597141,16.624945,17.585428,18.54591,19.506393,20.466877,21.423454,19.400974,17.378494,15.356014,13.333533,11.311053,10.963562,10.612165,10.260769,9.913278,9.561881,1.4875772,1.5070993,1.5266213,1.5461433,1.5656652,1.5890918,1.6242313,1.6593709,1.6906061,1.7257458,1.7608855,1.8038338,1.8428779,1.8819219,1.9209659,1.9639144,1.9912452,2.0224805,2.0537157,2.0810463,2.1122816,2.1044729,2.096664,2.0888553,2.0810463,2.0732377,2.1083772,2.1435168,2.1786566,2.2137961,2.2489357,2.8580225,3.4632049,4.0722914,4.6813784,5.2865605,6.196286,7.1060123,8.015738,8.929368,9.839094,8.183627,6.5281606,4.872694,3.2172275,1.5617609,1.4953861,1.4290112,1.358732,1.2923572,1.2259823,1.116659,1.0034313,0.8941081,0.78478485,0.6754616,0.63251317,0.58956474,0.5466163,0.5036679,0.46071947,0.40605783,0.3513962,0.29673457,0.24207294,0.18741131,0.1835069,0.1756981,0.1717937,0.1678893,0.1639849,0.15227169,0.14055848,0.13274968,0.12103647,0.113227665,0.10151446,0.093705654,0.08199245,0.07418364,0.062470436,0.07418364,0.08199245,0.093705654,0.10151446,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.042948425,0.08589685,0.12884527,0.1717937,0.21083772,0.4958591,0.77697605,1.0580931,1.3431144,1.6242313,2.1513257,2.67842,3.2094188,3.736513,4.263607,4.0801005,3.8965936,3.7130866,3.533484,3.349977,3.3343596,3.3187418,3.3031244,3.2914112,3.2757936,3.4514916,3.631094,3.8067923,3.9863946,4.1620927,4.1464753,4.126953,4.1113358,4.0918136,4.0761957,3.7911747,3.5100577,3.2289407,2.9439192,2.6628022,2.8385005,3.018103,3.193801,3.3734035,3.5491016,3.3265507,3.1000953,2.87364,2.6510892,2.4246337,2.7721257,3.1196175,3.4671092,3.814601,4.1620927,4.0215344,3.8770714,3.736513,3.59205,3.4514916,3.697469,3.9434462,4.193328,4.4393053,4.689187,4.564246,4.4432096,4.318269,4.1972322,4.0761957,4.1113358,4.1503797,4.1894236,4.224563,4.263607,4.2089458,4.1581883,4.1035266,4.0527697,3.998108,4.271416,4.5408196,4.8102236,5.0796275,5.349031,6.571109,7.793187,9.019169,10.241247,11.4633255,12.497992,13.532659,14.567325,15.601992,16.636658,16.30869,15.980719,15.656653,15.328683,15.000713,14.329156,13.653695,12.982138,12.31058,11.639023,11.014318,10.38571,9.761005,9.136301,8.511597,9.261242,10.010887,10.764437,11.514082,12.263727,12.431617,12.595602,12.763491,12.93138,13.09927,13.716166,14.329156,14.946052,15.559043,16.175938,16.441439,16.706938,16.968533,17.234032,17.49953,17.804073,18.104713,18.409256,18.709896,19.014439,19.045673,19.080814,19.115953,19.151093,19.186234,19.338505,19.486872,19.639143,19.78751,19.935879,18.807507,17.679134,16.546856,15.418485,14.286208,15.289639,16.29307,17.296501,18.296028,19.29946,20.54106,21.786564,23.028164,24.269764,25.511364,26.647545,27.783726,28.916002,30.052185,31.188366,34.667187,38.14601,41.62874,45.10756,48.58638,49.566387,50.54249,51.51859,52.498592,53.474693,51.78409,50.09348,48.40678,46.71617,45.025566,44.31887,43.616077,42.90938,42.20659,41.499893,35.67843,29.860868,24.039404,18.221846,12.400381,11.810817,11.225157,10.6355915,10.049932,9.464272,10.901091,12.341816,13.78254,15.223265,16.663988,17.4722,18.284315,19.092527,19.900738,20.712854,18.28822,15.863586,13.438952,11.014318,8.58578,8.929368,9.269051,9.608734,9.948417,10.2881,9.190963,8.097731,7.000593,5.9073606,4.814128,5.1186714,5.4271193,5.735567,6.044015,6.348558,7.47693,8.605303,9.733675,10.858143,11.986515,13.794253,15.598087,17.40192,19.205755,21.013493,21.013493,21.017397,21.021301,21.021301,21.025206,21.083773,21.138433,21.197,21.255566,21.314133,20.845604,20.377075,19.908546,19.443924,18.975395,20.092054,21.208714,22.329277,23.445936,24.562595,24.07845,23.598207,23.114061,22.63382,22.149673,20.388788,18.631807,16.870922,15.110037,13.349152,15.180316,17.01148,18.838741,20.669905,22.50107,19.428307,16.355541,13.282777,10.2100115,7.137247,5.8761253,4.618908,3.357786,2.096664,0.8394465,0.7106012,0.58175594,0.45681506,0.3279698,0.19912452,0.1639849,0.12884527,0.093705654,0.058566034,0.023426414,0.45681506,0.8862993,1.3157835,1.7452679,2.174752,2.3543546,2.533957,2.7135596,2.893162,3.076669,2.6823244,2.2918842,1.8975395,1.5031948,1.1127546,1.6710842,2.2294137,2.7838387,3.3421683,3.900498,4.0488653,4.193328,4.3416953,4.4900627,4.6384296,4.6930914,4.747753,4.802415,4.8570766,4.911738,5.4036927,5.8956475,6.3915067,6.883461,7.375416,7.629202,7.8790836,8.13287,8.386656,8.636538,9.0465,9.452558,9.858616,10.268578,10.674636,10.955752,11.240774,11.521891,11.806912,12.08803,12.271536,12.458947,12.642454,12.825961,13.013372,12.423808,11.838148,11.248583,10.662923,10.073358,9.686822,9.300286,8.913751,8.52331,8.136774,7.6409154,7.141152,6.6452928,6.1494336,5.64967,6.27047,6.89127,7.5081654,8.128965,8.749765,10.768341,12.783013,14.801589,16.820166,18.838741,23.399082,27.95552,32.51586,37.076202,41.636547,39.00498,36.373413,33.741844,31.106373,28.474806,26.792007,25.109211,23.426414,21.743616,20.06082,21.415646,22.774378,24.129206,25.484034,26.838861,24.222912,21.606962,18.991013,16.378967,13.763018,14.243259,14.727406,15.211552,15.6917925,16.175938,13.907481,11.639023,9.370565,7.1060123,4.8375545,11.186112,17.538574,23.887133,30.235691,36.588154,30.840874,25.097498,19.354122,13.606842,7.8634663,8.36323,8.862993,9.362757,9.86252,10.362284,9.280765,8.203149,7.1216297,6.044015,4.9624953,5.0913405,5.22409,5.3529353,5.481781,5.610626,5.9815445,6.348558,6.715572,7.082586,7.4495993,8.554545,9.659492,10.764437,11.869383,12.974329,12.603411,12.236397,11.8654785,11.49456,11.123642,10.826907,10.530173,10.2334385,9.936704,9.636065,10.373997,11.111929,11.849861,12.587793,13.325725,14.044135,14.766449,15.484859,16.20327,16.925583,17.456583,17.983677,18.514675,19.045673,19.576674,19.190138,18.8036,18.420969,18.034433,17.651802,17.167656,16.683512,16.20327,15.719124,15.238882,15.086611,14.934339,14.778163,14.625891,14.473619,13.938716,13.403813,12.86891,12.334006,11.799104,11.537509,11.275913,11.014318,10.748819,10.487225,10.994797,11.502369,12.009941,12.517513,13.025085,12.619028,12.209065,11.803008,11.39695,10.986988,10.741011,10.491129,10.2451515,9.999174,9.749292,8.8083315,7.8634663,6.9225054,5.9815445,5.036679,5.3021784,5.5676775,5.833177,6.098676,6.364176,7.1177254,7.871275,8.628729,9.382278,10.135828,10.721489,11.303245,11.885,12.466757,13.048512,13.364769,13.6810255,13.993378,14.309634,14.625891,16.015858,17.405825,18.795792,20.18576,21.575727,21.431265,21.2868,21.138433,20.99397,20.849508,20.181856,19.514202,18.84655,18.178898,17.511244,17.733795,17.956347,18.178898,18.401447,18.623999,19.463446,20.298986,21.138433,21.973976,22.813423,22.7939,22.778282,22.75876,22.743143,22.723621,21.903696,21.083773,20.263847,19.443924,18.623999,19.693806,20.76361,21.833418,22.903223,23.976934,23.570877,23.164818,22.75876,22.356607,21.95055,20.83389,19.721136,18.604477,17.491722,16.375063,17.253553,18.132044,19.00663,19.88512,20.76361,18.983204,17.206701,15.430198,13.653695,11.873287,11.611692,11.350098,11.088503,10.826907,10.561408,1.4641509,1.4836729,1.5070993,1.5305257,1.5539521,1.5734742,1.6047094,1.6359446,1.6632754,1.6945106,1.7257458,1.7843118,1.8389735,1.8975395,1.9561055,2.0107672,2.0380979,2.069333,2.096664,2.1239948,2.1513257,2.1513257,2.15523,2.1591344,2.1591344,2.1630387,2.1786566,2.1981785,2.2137961,2.233318,2.2489357,3.084478,3.9200199,4.755562,5.591104,6.426646,6.715572,7.008402,7.3012323,7.5940623,7.8868923,6.5867267,5.282656,3.978586,2.67842,1.3743496,1.2962615,1.2181735,1.1439898,1.0659018,0.9878138,0.9058213,0.8277333,0.74574083,0.6676528,0.58566034,0.5466163,0.5075723,0.46852827,0.42557985,0.38653582,0.3474918,0.30844778,0.26940376,0.22645533,0.18741131,0.1717937,0.15617609,0.14055848,0.12884527,0.113227665,0.10932326,0.10151446,0.09761006,0.093705654,0.08589685,0.08199245,0.078088045,0.07418364,0.06637484,0.062470436,0.078088045,0.09761006,0.113227665,0.13274968,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.43338865,0.7340276,1.0307622,1.3274968,1.6242313,2.0068626,2.3894942,2.7721257,3.154757,3.5373883,3.4514916,3.3655949,3.2836022,3.1977055,3.1118085,3.1313305,3.1469483,3.1664703,3.182088,3.2016098,3.3343596,3.4632049,3.5959544,3.7287042,3.8614538,3.8341231,3.8067923,3.7794614,3.7521305,3.7247996,3.4632049,3.2055142,2.9439192,2.6862288,2.4246337,2.7213683,3.0141985,3.310933,3.6037633,3.900498,3.5373883,3.174279,2.8111696,2.4480603,2.0888553,2.6159496,3.1469483,3.677947,4.2089458,4.73604,4.4861584,4.2323723,3.978586,3.7287042,3.474918,3.7443218,4.009821,4.279225,4.5447245,4.814128,4.521298,4.2284675,3.9356375,3.6428072,3.349977,3.3734035,3.4007344,3.4241607,3.4514916,3.474918,3.49444,3.5100577,3.5256753,3.5451972,3.5608149,3.7599394,3.959064,4.154284,4.3534083,4.548629,5.5676775,6.5867267,7.601871,8.62092,9.636065,10.979179,12.322293,13.665408,15.008522,16.351637,15.855778,15.359919,14.864059,14.3682,13.8762455,13.095366,12.314485,11.533605,10.756628,9.975748,9.526741,9.073831,8.624825,8.175818,7.726812,8.550641,9.37447,10.198298,11.0260315,11.849861,12.013845,12.181735,12.34572,12.509705,12.67369,13.384291,14.090988,14.797685,15.504381,16.211079,16.29307,16.378967,16.46096,16.542952,16.624945,17.070047,17.515148,17.96025,18.405352,18.850454,18.64352,18.436588,18.22575,18.018816,17.811884,17.487818,17.163752,16.835783,16.511717,16.187653,15.258404,14.33306,13.403813,12.47847,11.549222,13.130505,14.7156925,16.296974,17.878258,19.463446,20.779228,22.091108,23.40689,24.722675,26.038458,27.479183,28.923813,30.364536,31.809166,33.24989,36.275803,39.30562,42.331528,45.361347,48.387257,50.48392,52.57668,54.673344,56.766106,58.86277,57.26587,55.67287,54.07597,52.482975,50.886074,49.460968,48.031956,46.60685,45.177837,43.74883,37.041065,30.329397,23.621634,16.909966,10.198298,9.901564,9.600925,9.300286,8.999647,8.699008,11.033841,13.364769,15.695697,18.030529,20.361458,20.416119,20.470781,20.529346,20.58401,20.63867,18.038338,15.438006,12.837675,10.237343,7.6370106,8.105539,8.577971,9.0465,9.518932,9.987461,8.913751,7.843944,6.7702336,5.6965227,4.6267166,5.0483923,5.4700675,5.891743,6.3134184,6.7389984,7.6682463,8.601398,9.534551,10.467703,11.400854,13.314012,15.231073,17.14423,19.061293,20.97445,21.271183,21.564014,21.860748,22.153578,22.450314,22.485453,22.520592,22.555733,22.590872,22.62601,21.673336,20.720663,19.767988,18.815315,17.86264,20.127193,22.391747,24.6563,26.920853,29.189312,27.650976,26.116547,24.582117,23.047686,21.513256,19.346313,17.17937,15.008522,12.841579,10.674636,13.501423,16.32821,19.158901,21.98569,24.812477,21.470308,18.12814,14.785972,11.443803,8.101635,6.6687193,5.239708,3.8106966,2.3816853,0.94876975,0.80430686,0.659844,0.5153811,0.3709182,0.22645533,0.1835069,0.14055848,0.09761006,0.05466163,0.011713207,0.41386664,0.8160201,1.2181735,1.6242313,2.0263848,2.25284,2.4792955,2.7057507,2.9361105,3.1625657,2.7096553,2.2567444,1.8038338,1.3509232,0.9019169,1.43682,1.9717231,2.5066261,3.0415294,3.5764325,3.6545205,3.736513,3.814601,3.8965936,3.9746814,4.1894236,4.4041657,4.618908,4.83365,5.0483923,5.388075,5.7316628,6.0713453,6.4110284,6.7507114,6.7702336,6.7897553,6.8092775,6.8287997,6.8483214,7.473026,8.093826,8.718531,9.339331,9.964035,9.846903,9.733675,9.616543,9.503315,9.386183,9.768814,10.147541,10.526268,10.9089,11.287627,10.975275,10.662923,10.350571,10.0382185,9.725866,9.311999,8.898132,8.488171,8.074304,7.6643414,7.195813,6.727285,6.2587566,5.794133,5.3256044,5.5989127,5.8683167,6.141625,6.4149327,6.688241,9.928895,13.165645,16.406298,19.646952,22.887606,26.479656,30.071707,33.663757,37.255806,40.85176,36.978592,33.105427,29.23226,25.359093,21.485926,21.228235,20.96664,20.70895,20.447355,20.18576,21.177479,22.169195,23.15701,24.148727,25.136541,23.266333,21.396124,19.525915,17.655706,15.789403,15.54733,15.309161,15.067088,14.828919,14.586847,12.533132,10.48332,8.429605,6.375889,4.3260775,11.23687,18.151566,25.062359,31.977055,38.887848,32.090282,25.292717,18.495153,11.697589,4.900025,5.7238536,6.551587,7.375416,8.1992445,9.023073,7.9727893,6.918601,5.8683167,4.814128,3.7638438,3.5881457,3.416352,3.2445583,3.0727646,2.900971,3.0883822,3.279698,3.4710135,3.6584249,3.8497405,4.6267166,5.4036927,6.180669,6.9615493,7.7385254,7.5667315,7.3910336,7.2192397,7.0474463,6.8756523,6.9459314,7.016211,7.08649,7.1567693,7.223144,7.8634663,8.499884,9.136301,9.776623,10.413041,11.549222,12.681499,13.817679,14.95386,16.086138,16.164225,16.242313,16.320402,16.398489,16.476578,15.793307,15.113941,14.434575,13.755209,13.075843,13.477997,13.88015,14.282304,14.684457,15.086611,15.1061325,15.12175,15.141272,15.15689,15.176412,14.458001,13.739592,13.021181,12.306676,11.588266,11.213444,10.838621,10.4637985,10.088976,9.714153,9.96013,10.206107,10.455989,10.701966,10.951848,10.815194,10.67854,10.545791,10.409137,10.276386,10.182681,10.088976,9.999174,9.905469,9.811763,8.784905,7.758047,6.7311897,5.704332,4.6735697,4.7828927,4.8883114,4.997635,5.1030536,5.212377,5.7785153,6.3407493,6.9068875,7.473026,8.039165,9.561881,11.080693,12.603411,14.126127,15.648844,15.781594,15.914344,16.047092,16.179844,16.312593,18.007103,19.701614,21.396124,23.090635,24.78905,23.965221,23.141392,22.321468,21.497639,20.67381,19.846077,19.018343,18.19061,17.366781,16.539047,16.429726,16.324306,16.214983,16.10566,16.00024,17.24965,18.499058,19.748466,21.00178,22.251188,22.29804,22.344894,22.391747,22.4386,22.489357,21.591345,20.693333,19.795319,18.897306,17.999294,19.073006,20.146715,21.216522,22.290232,23.363943,23.172626,22.981312,22.7939,22.602585,22.411268,21.15405,19.896833,18.639616,17.382399,16.125181,16.921679,17.714273,18.51077,19.303364,20.099863,18.569338,17.034906,15.504381,13.969952,12.439425,12.263727,12.08803,11.912332,11.736633,11.560935,1.43682,1.4641509,1.4875772,1.5110037,1.5383345,1.5617609,1.5890918,1.6125181,1.6359446,1.6632754,1.6867018,1.7608855,1.8389735,1.9131571,1.9873407,2.0615244,2.0888553,2.1122816,2.135708,2.1630387,2.1864653,2.1981785,2.2137961,2.2255092,2.2372224,2.2489357,2.2489357,2.2489357,2.2489357,2.2489357,2.2489357,3.310933,4.376835,5.4388323,6.5008297,7.562827,7.238762,6.910792,6.5867267,6.262661,5.938596,4.985922,4.037152,3.0883822,2.135708,1.1869383,1.1010414,1.0112402,0.92534333,0.8394465,0.74964523,0.698888,0.6481308,0.60127795,0.5505207,0.4997635,0.46071947,0.42557985,0.38653582,0.3513962,0.31235218,0.28892577,0.26159495,0.23816854,0.21083772,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.37482262,0.6871748,0.999527,1.3118792,1.6242313,1.8623998,2.1005683,2.338737,2.5769055,2.8111696,2.8267872,2.8385005,2.8502135,2.8619268,2.87364,2.9243972,2.9751544,3.0259118,3.076669,3.1235218,3.213323,3.2992198,3.3890212,3.474918,3.5608149,3.5256753,3.4866312,3.4514916,3.4124475,3.3734035,3.1391394,2.900971,2.6628022,2.4246337,2.1864653,2.6003318,3.0141985,3.4241607,3.8380275,4.251894,3.7482262,3.2484627,2.7486992,2.2489357,1.7491722,2.463678,3.174279,3.8887846,4.5993857,5.3138914,4.950782,4.5876727,4.224563,3.8614538,3.4983444,3.78727,4.0761957,4.3612175,4.650143,4.939069,4.474445,4.0137253,3.5491016,3.0883822,2.6237583,2.639376,2.6510892,2.6628022,2.6745155,2.6862288,2.77603,2.8619268,2.951728,3.0376248,3.1235218,3.2484627,3.3734035,3.4983444,3.6232853,3.7482262,4.564246,5.376362,6.1884775,7.000593,7.812709,9.464272,11.111929,12.763491,14.411149,16.062712,15.398962,14.739119,14.07537,13.411622,12.751778,11.861574,10.975275,10.088976,9.198771,8.312472,8.039165,7.7619514,7.4886436,7.211431,6.9381227,7.8361354,8.738052,9.636065,10.537982,11.435994,11.599979,11.763964,11.924045,12.08803,12.24811,13.048512,13.848915,14.649317,15.449719,16.250122,16.148607,16.050997,15.949483,15.851873,15.750359,16.33602,16.925583,17.511244,18.10081,18.68647,18.237463,17.788456,17.335546,16.88654,16.437534,15.637131,14.836729,14.036326,13.235924,12.439425,11.713207,10.986988,10.260769,9.538455,8.812236,10.975275,13.138313,15.3013525,17.464392,19.623526,21.013493,22.399555,23.785618,25.175587,26.56165,28.310822,30.063898,31.81307,33.56224,35.311413,37.88832,40.46132,43.038227,45.61123,48.188133,51.401455,54.610874,57.824196,61.03752,64.25085,62.751553,61.24836,59.74907,58.24978,56.75049,54.59916,52.45174,50.300415,48.14909,46.001667,38.399796,30.80183,23.199959,15.598087,8.00012,7.988407,7.9766936,7.9610763,7.9493628,7.9376497,11.162686,14.387722,17.612759,20.837795,24.062832,23.363943,22.66115,21.962263,21.263374,20.560583,17.788456,15.012426,12.236397,9.464272,6.688241,7.2856145,7.8868923,8.488171,9.089449,9.686822,8.636538,7.5862536,6.5359693,5.4856853,4.4393053,4.9742084,5.5130157,6.0518236,6.5867267,7.125534,7.8634663,8.601398,9.339331,10.073358,10.81129,12.837675,14.864059,16.88654,18.912924,20.93931,21.52497,22.11063,22.700195,23.285854,23.87542,23.887133,23.898846,23.910559,23.926178,23.937891,22.50107,21.06425,19.623526,18.186707,16.749886,20.162333,23.574781,26.987228,30.399675,33.812122,31.223505,28.63879,26.05017,23.461554,20.876839,18.299932,15.726933,13.150026,10.573121,8.00012,11.826434,15.648844,19.475159,23.301472,27.123882,23.51231,19.900738,16.289165,12.67369,9.062118,7.461313,5.8644123,4.263607,2.6628022,1.0619974,0.9019169,0.737932,0.57394713,0.41386664,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.37482262,0.74964523,1.1244678,1.4992905,1.8741131,2.1513257,2.4246337,2.7018464,2.9751544,3.2484627,2.736986,2.2255092,1.7140326,1.1986516,0.6871748,1.1986516,1.7140326,2.2255092,2.736986,3.2484627,3.2640803,3.2757936,3.2875066,3.2992198,3.310933,3.6857557,4.0605783,4.4393053,4.814128,5.1889505,5.376362,5.563773,5.7511845,5.938596,6.126007,5.911265,5.700427,5.4856853,5.2748475,5.0640097,5.899552,6.7389984,7.57454,8.413987,9.249529,8.738052,8.226576,7.7111945,7.1997175,6.688241,7.262188,7.8361354,8.413987,8.987934,9.561881,9.526741,9.487698,9.448653,9.413514,9.37447,8.937177,8.499884,8.062591,7.6252975,7.1880045,6.7507114,6.3134184,5.8761253,5.4388323,5.001539,4.9234514,4.8492675,4.775084,4.7009,4.6267166,9.089449,13.548276,18.011007,22.47374,26.936472,29.564135,32.187893,34.81165,37.439312,40.063072,34.948303,29.837442,24.72658,19.611813,14.50095,15.664462,16.82407,17.987581,19.151093,20.310701,20.93931,21.564014,22.188719,22.813423,23.438128,22.31366,21.189192,20.06082,18.936352,17.811884,16.8514,15.8870125,14.92653,13.962143,13.001659,11.162686,9.323712,7.4886436,5.64967,3.8106966,11.287627,18.760653,26.237583,33.71451,41.18754,33.335785,25.487938,17.636185,9.788337,1.9365835,3.0883822,4.2362766,5.388075,6.5359693,7.687768,6.66091,5.6379566,4.6110992,3.5881457,2.5612879,2.0888553,1.6125181,1.1361811,0.6637484,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,0.698888,1.1517987,1.6008049,2.0498111,2.4988174,2.5261483,2.5495746,2.5769055,2.6003318,2.6237583,3.0610514,3.4983444,3.9356375,4.376835,4.814128,5.349031,5.8878384,6.426646,6.9615493,7.5003567,9.050405,10.600452,12.150499,13.700547,15.250595,14.875772,14.50095,14.126127,13.751305,13.376482,12.400381,11.424281,10.44818,9.475985,8.499884,9.788337,11.076789,12.361338,13.64979,14.938243,15.125654,15.313066,15.500477,15.687888,15.875299,14.973383,14.07537,13.173453,12.27544,11.373524,10.889378,10.401327,9.913278,9.425227,8.937177,8.925464,8.913751,8.898132,8.886419,8.874706,9.01136,9.151918,9.288573,9.425227,9.561881,9.6243515,9.686822,9.749292,9.811763,9.874233,8.761478,7.648724,6.5359693,5.423215,4.3143644,4.263607,4.21285,4.1620927,4.1113358,4.0605783,4.4393053,4.814128,5.1889505,5.563773,5.938596,8.398369,10.862047,13.325725,15.785499,18.249176,18.19842,18.151566,18.10081,18.05005,17.999294,19.998348,22.001307,24.00036,25.999414,27.998468,26.499178,24.999887,23.500597,22.001307,20.498112,19.514202,18.526388,17.538574,16.55076,15.562947,15.125654,14.688361,14.251068,13.813775,13.376482,15.035853,16.69913,18.362404,20.025679,21.688955,21.798277,21.911505,22.024733,22.13796,22.251188,21.275087,20.298986,19.326792,18.35069,17.37459,18.448301,19.525915,20.599627,21.673336,22.750952,22.774378,22.801708,22.825136,22.848562,22.875893,21.474213,20.076437,18.674755,17.27698,15.875299,16.585901,17.300406,18.011007,18.725513,19.436115,18.151566,16.863113,15.57466,14.286208,13.001659,12.911859,12.825961,12.73616,12.650263,12.564366,1.4251068,1.4485333,1.475864,1.4992905,1.5266213,1.5500476,1.5812829,1.6164225,1.6476578,1.678893,1.7140326,1.7882162,1.8663043,1.9443923,2.0224805,2.1005683,2.135708,2.1708477,2.2059872,2.241127,2.2762666,2.2840753,2.2957885,2.3035975,2.3153105,2.3231194,2.3035975,2.280171,2.2567444,2.233318,2.2137961,3.4514916,4.6930914,5.930787,7.172387,8.413987,7.816613,7.2192397,6.621866,6.0205884,5.423215,4.5681505,3.7091823,2.854118,1.9951496,1.1361811,1.0541886,0.96829176,0.8823949,0.79649806,0.7106012,0.6715572,0.63251317,0.59346914,0.5544251,0.5114767,0.47633708,0.43729305,0.39824903,0.3631094,0.3240654,0.29673457,0.26549935,0.23426414,0.20693332,0.1756981,0.15227169,0.12884527,0.10932326,0.08589685,0.062470436,0.06637484,0.06637484,0.07027924,0.07418364,0.07418364,0.078088045,0.08589685,0.08980125,0.093705654,0.10151446,0.113227665,0.12884527,0.14446288,0.16008049,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.25769055,0.21474212,0.1717937,0.12884527,0.08589685,0.3435874,0.59737355,0.8511597,1.1088502,1.3626363,1.542239,1.7218413,1.901444,2.0810463,2.260649,2.2762666,2.2879796,2.2996929,2.3114061,2.3231194,2.4012074,2.4792955,2.5573835,2.6354716,2.7135596,2.7565079,2.803361,2.8463092,2.893162,2.9361105,2.9048753,2.87364,2.8385005,2.8072653,2.77603,2.6354716,2.494913,2.3543546,2.2137961,2.0732377,2.3816853,2.6862288,2.9907722,3.2953155,3.5998588,3.213323,2.8267872,2.436347,2.0498111,1.6632754,2.3270237,2.9907722,3.6584249,4.322173,4.985922,4.786797,4.5837684,4.380739,4.1777105,3.9746814,4.1581883,4.3416953,4.521298,4.704805,4.8883114,4.4393053,3.9863946,3.5373883,3.0883822,2.639376,2.6549935,2.6706111,2.690133,2.7057507,2.7252727,2.7643168,2.803361,2.8463092,2.8853533,2.9243972,3.232845,3.541293,3.8458362,4.154284,4.462732,5.12648,5.794133,6.4578815,7.1216297,7.7892823,9.17925,10.569217,11.959184,13.349152,14.739119,14.239355,13.735687,13.235924,12.73616,12.236397,11.39695,10.553599,9.710248,8.866898,8.023546,7.746334,7.4691215,7.191909,6.914696,6.6374836,7.519879,8.402273,9.284669,10.167064,11.0494585,11.381332,11.709302,12.041177,12.369146,12.70102,13.25935,13.813775,14.372105,14.930434,15.488764,15.141272,14.79378,14.446288,14.098797,13.751305,14.727406,15.7035055,16.683512,17.65961,18.635712,18.151566,17.663515,17.175465,16.687416,16.199366,15.395058,14.590752,13.786445,12.978233,12.173926,12.24811,12.326198,12.400381,12.4745655,12.548749,14.317443,16.086138,17.850927,19.619621,21.388315,22.47374,23.563068,24.64849,25.73782,26.823244,28.42405,30.024853,31.625658,33.226463,34.823364,37.575966,40.32857,43.081173,45.83378,48.58638,52.170624,55.75096,59.3352,62.91944,66.49978,64.81308,63.126377,61.43577,59.74907,58.062366,55.153587,52.240902,49.332123,46.423344,43.51066,36.8068,30.099037,23.391273,16.683512,9.975748,10.061645,10.143637,10.229534,10.315431,10.401327,12.6463585,14.89139,17.136421,19.381453,21.626484,23.84809,26.069695,28.291298,30.516808,32.738415,28.338152,23.937891,19.537628,15.137367,10.737106,10.295909,9.850807,9.40961,8.968412,8.52331,8.113348,7.703386,7.2934237,6.883461,6.473499,7.0786815,7.6799593,8.281238,8.886419,9.487698,10.491129,11.490656,12.494087,13.497519,14.50095,16.296974,18.089096,19.88512,21.681147,23.473267,24.316618,25.159967,26.003319,26.84667,27.686117,27.666594,27.647072,27.62755,27.608028,27.588507,25.761246,23.937891,22.11063,20.287273,18.463919,20.74409,23.02426,25.304432,27.580698,29.860868,27.350338,24.835903,22.325373,19.810938,17.300406,15.14908,12.993851,10.8425255,8.691199,6.5359693,9.6243515,12.708829,15.793307,18.877785,21.962263,19.053482,16.140799,13.232019,10.323239,7.4105554,6.1064854,4.802415,3.4983444,2.194274,0.8862993,1.1791295,1.4719596,1.7647898,2.05762,2.35045,1.9951496,1.639849,1.2845483,0.92924774,0.57394713,0.8589685,1.1400855,1.4212024,1.7062237,1.9873407,2.1981785,2.4090161,2.6159496,2.8267872,3.0376248,2.5964274,2.1591344,1.717937,1.2767396,0.8394465,1.2650263,1.6906061,2.1200905,2.5456703,2.9751544,3.0259118,3.076669,3.1235218,3.174279,3.2250361,3.49444,3.7638438,4.0332475,4.3065557,4.575959,4.759466,4.9468775,5.1303844,5.3138914,5.5013027,5.364649,5.2318993,5.095245,4.958591,4.825841,5.5832953,6.3407493,7.098203,7.8556576,8.6131115,8.156297,7.703386,7.2465706,6.79366,6.336845,6.7663293,7.191909,7.621393,8.046973,8.476458,8.429605,8.386656,8.339804,8.296855,8.250002,7.968885,7.6838636,7.4027467,7.1216297,6.8366084,6.4188375,6.001066,5.5832953,5.169429,4.7516575,4.6540475,4.560342,4.466636,4.369026,4.2753205,8.644346,13.009468,17.378494,21.743616,26.112642,27.775917,29.439194,31.098564,32.76184,34.425114,30.356728,26.28834,22.223858,18.15547,14.087084,15.402867,16.71865,18.034433,19.346313,20.662096,21.177479,21.69286,22.20824,22.723621,23.239002,22.130152,21.021301,19.916355,18.807507,17.698656,16.835783,15.976814,15.113941,14.251068,13.388195,12.150499,10.912805,9.675109,8.437413,7.1997175,12.494087,17.784552,23.078922,28.369387,33.663757,28.892576,24.121397,19.354122,14.582942,9.811763,9.448653,9.089449,8.726339,8.36323,8.00012,7.0708723,6.141625,5.2084727,4.279225,3.349977,2.7096553,2.069333,1.4290112,0.78868926,0.14836729,0.16008049,0.1717937,0.1796025,0.19131571,0.19912452,0.5583295,0.92143893,1.2806439,1.639849,1.999054,2.018576,2.0380979,2.0615244,2.0810463,2.1005683,2.4519646,2.7994564,3.1508527,3.4983444,3.8497405,4.283129,4.716518,5.1460023,5.579391,6.012779,7.2543793,8.492075,9.733675,10.971371,12.212971,11.912332,11.611692,11.311053,11.014318,10.71368,9.952321,9.190963,8.433509,7.6721506,6.910792,8.265619,9.616543,10.971371,12.322293,13.673217,14.157363,14.641508,15.12175,15.605896,16.086138,15.176412,14.262781,13.349152,12.439425,11.525795,11.447707,11.369619,11.291532,11.213444,11.139259,11.100216,11.061172,11.0260315,10.986988,10.951848,10.795672,10.639496,10.48332,10.331048,10.174872,10.2100115,10.2451515,10.280292,10.315431,10.350571,9.499411,8.648251,7.800996,6.949836,6.098676,6.153338,6.2040954,6.2587566,6.309514,6.364176,6.688241,7.012306,7.336372,7.6643414,7.988407,10.0265045,12.068507,14.106606,16.148607,18.186707,18.10081,18.011007,17.92511,17.839214,17.749413,19.178425,20.60353,22.032541,23.461554,24.88666,23.531832,22.177006,20.822178,19.46735,18.112522,17.206701,16.300879,15.398962,14.493141,13.58732,13.306203,13.028991,12.747873,12.466757,12.185639,13.837202,15.488764,17.136421,18.787983,20.435642,20.509825,20.58401,20.654287,20.728472,20.79875,20.021774,19.240894,18.460014,17.679134,16.898252,18.011007,19.123762,20.236517,21.349272,22.462027,22.668959,22.871988,23.078922,23.28195,23.488884,22.27071,21.052536,19.834364,18.61619,17.40192,18.073479,18.74894,19.4244,20.099863,20.775324,19.326792,17.878258,16.43363,14.985096,13.536563,13.196879,12.857197,12.517513,12.177831,11.838148,1.4133936,1.43682,1.4641509,1.4875772,1.5110037,1.5383345,1.5773785,1.6164225,1.6593709,1.698415,1.737459,1.815547,1.8975395,1.9756275,2.05762,2.135708,2.182561,2.2294137,2.2723622,2.3192148,2.3621633,2.3699722,2.377781,2.3855898,2.3933985,2.4012074,2.3543546,2.3114061,2.2645533,2.2216048,2.174752,3.59205,5.009348,6.426646,7.843944,9.261242,8.3944645,7.523783,6.6531014,5.7824197,4.911738,4.1464753,3.3812122,2.6159496,1.8506867,1.0893283,1.0034313,0.92143893,0.8394465,0.75745404,0.6754616,0.6442264,0.61689556,0.58566034,0.5544251,0.5231899,0.48805028,0.44900626,0.41386664,0.37482262,0.3357786,0.30063897,0.26940376,0.23426414,0.19912452,0.1639849,0.14055848,0.12103647,0.10151446,0.08199245,0.062470436,0.06637484,0.07418364,0.078088045,0.08199245,0.08589685,0.09761006,0.10932326,0.11713207,0.12884527,0.13665408,0.14055848,0.14836729,0.15227169,0.15617609,0.1639849,0.12884527,0.09761006,0.06637484,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12103647,0.23816854,0.359205,0.48024148,0.60127795,0.5036679,0.40605783,0.30844778,0.21083772,0.113227665,0.30844778,0.5075723,0.7066968,0.9019169,1.1010414,1.2220778,1.3431144,1.4680552,1.5890918,1.7140326,1.7257458,1.737459,1.7491722,1.7608855,1.7765031,1.8819219,1.9834363,2.0888553,2.194274,2.2996929,2.3035975,2.3035975,2.3075018,2.3114061,2.3114061,2.2840753,2.2567444,2.2294137,2.2020829,2.174752,2.1318035,2.0888553,2.0459068,2.0068626,1.9639144,2.1591344,2.358259,2.5534792,2.7526035,2.951728,2.6745155,2.4012074,2.1239948,1.8506867,1.5734742,2.194274,2.8111696,3.4280653,4.044961,4.661856,4.618908,4.575959,4.5369153,4.493967,4.4510183,4.5291066,4.60329,4.6813784,4.759466,4.8375545,4.4002614,3.9629683,3.5256753,3.0883822,2.6510892,2.6706111,2.6940374,2.717464,2.7408905,2.7643168,2.7565079,2.7486992,2.7408905,2.7330816,2.7252727,3.213323,3.7052777,4.193328,4.6852827,5.173333,5.6926184,6.211904,6.727285,7.2465706,7.7619514,8.894228,10.0226,11.150972,12.28325,13.411622,13.075843,12.73616,12.400381,12.0606985,11.72492,10.928422,10.131924,9.331521,8.535024,7.7385254,7.4574084,7.1762915,6.899079,6.617962,6.336845,7.2036223,8.066495,8.933272,9.796145,10.662923,11.158782,11.6585455,12.154405,12.654168,13.150026,13.466284,13.778636,14.0948925,14.411149,14.723501,14.130032,13.536563,12.939189,12.34572,11.748346,13.118792,14.4853325,15.851873,17.218414,18.58886,18.061766,17.538574,17.01148,16.48829,15.961197,15.152986,14.34087,13.532659,12.720543,11.912332,12.786918,13.661504,14.53609,15.410676,16.289165,17.65961,19.03396,20.404406,21.778755,23.1492,23.937891,24.72658,25.511364,26.300053,27.088743,28.537275,29.98581,31.438248,32.88678,34.33922,37.26752,40.19582,43.12803,46.056328,48.988537,52.93979,56.891045,60.846207,64.79746,68.74872,66.8746,65.00049,63.126377,61.24836,59.374245,55.704105,52.03397,48.36383,44.69369,41.023556,35.2099,29.396244,23.578686,17.76503,11.951375,12.130978,12.314485,12.497992,12.681499,12.861101,14.126127,15.391153,16.65618,17.921206,19.186234,24.332235,29.478237,34.62424,39.76634,44.91234,38.887848,32.863354,26.838861,20.81437,14.785972,13.302299,11.818625,10.331048,8.847376,7.363703,7.5940623,7.824422,8.050878,8.281238,8.511597,9.17925,9.846903,10.514555,11.182208,11.849861,13.118792,14.383818,15.652749,16.921679,18.186707,19.75237,21.318037,22.883701,24.449368,26.011127,27.108265,28.209307,29.306444,30.40358,31.500717,31.446056,31.395298,31.340637,31.289879,31.239122,29.025326,26.811531,24.601639,22.387842,20.174046,21.321941,22.469835,23.61773,24.765623,25.913517,23.473267,21.036919,18.600573,16.164225,13.723974,11.994324,10.264673,8.535024,6.805373,5.0757227,7.4183645,9.76491,12.111456,14.454097,16.800642,14.590752,12.384764,10.178777,7.968885,5.7628975,4.7516575,3.7443218,2.7330816,1.7218413,0.7106012,1.4602464,2.2059872,2.9556324,3.7013733,4.4510183,3.7911747,3.1313305,2.4714866,1.8116426,1.1517987,1.33921,1.5305257,1.7218413,1.9092526,2.1005683,2.2450314,2.3894942,2.533957,2.67842,2.8267872,2.455869,2.0888553,1.7218413,1.3548276,0.9878138,1.3314011,1.6710842,2.0146716,2.358259,2.7018464,2.787743,2.87364,2.9634414,3.049338,3.1391394,3.3031244,3.4671092,3.631094,3.7989833,3.9629683,4.1464753,4.3260775,4.5095844,4.6930914,4.8765984,4.8180323,4.759466,4.7009,4.646239,4.5876727,5.263134,5.9425,6.621866,7.297328,7.9766936,7.578445,7.180196,6.7819467,6.3836975,5.989353,6.266566,6.547683,6.8287997,7.1060123,7.387129,7.336372,7.28171,7.230953,7.1762915,7.125534,6.996689,6.871748,6.7429028,6.6140575,6.4891167,6.0908675,5.6926184,5.2943697,4.8961205,4.5017757,4.3846436,4.271416,4.154284,4.041056,3.9239242,8.1992445,12.470661,16.742077,21.013493,25.288813,25.987701,26.68659,27.389381,28.08827,28.787157,25.76515,22.743143,19.721136,16.69913,13.673217,15.141272,16.609327,18.077383,19.545437,21.013493,21.415646,21.821705,22.227762,22.63382,23.035973,21.946646,20.857317,19.767988,18.678661,17.589333,16.82407,16.062712,15.3013525,14.53609,13.774731,13.138313,12.501896,11.861574,11.225157,10.588739,13.696643,16.808453,19.916355,23.028164,26.136068,24.445463,22.75876,21.068155,19.377548,17.686943,15.812829,13.938716,12.0606985,10.186585,8.312472,7.47693,6.6413884,5.805846,4.9742084,4.138666,3.3343596,2.5261483,1.7218413,0.91753453,0.113227665,0.12103647,0.12884527,0.13665408,0.14055848,0.14836729,0.42167544,0.6910792,0.96048295,1.2298868,1.4992905,1.5149081,1.5305257,1.5461433,1.5617609,1.5734742,1.8389735,2.1005683,2.3621633,2.6237583,2.8892577,3.213323,3.541293,3.8692627,4.1972322,4.5252023,5.45445,6.3836975,7.3168497,8.246098,9.175345,8.94889,8.726339,8.499884,8.273428,8.050878,7.504261,6.9615493,6.4149327,5.8683167,5.3256044,6.7429028,8.160201,9.577498,10.994797,12.412095,13.189071,13.966047,14.746927,15.523903,16.300879,15.375536,14.450192,13.524849,12.599506,11.674163,12.006037,12.341816,12.67369,13.005564,13.337439,13.274967,13.212498,13.150026,13.087557,13.025085,12.576079,12.130978,11.681972,11.23687,10.787864,10.795672,10.803481,10.81129,10.819098,10.826907,10.237343,9.651682,9.062118,8.476458,7.8868923,8.043069,8.1992445,8.351517,8.507692,8.663869,8.937177,9.21439,9.487698,9.761005,10.0382185,11.654641,13.271063,14.89139,16.507812,18.124235,17.999294,17.874353,17.749413,17.624472,17.49953,18.354595,19.20966,20.064724,20.919786,21.77485,20.564487,19.354122,18.143757,16.933393,15.726933,14.903104,14.079274,13.25935,12.435521,11.611692,11.490656,11.365715,11.2446785,11.123642,10.998701,12.63855,14.274494,15.914344,17.550287,19.186234,19.221373,19.252607,19.283842,19.318983,19.350218,18.764557,18.178898,17.593237,17.01148,16.42582,17.573715,18.725513,19.873407,21.025206,22.1731,22.559637,22.946173,23.328804,23.71534,24.101875,23.063305,22.028637,20.99397,19.959305,18.924637,19.561056,20.201378,20.837795,21.474213,22.11063,20.50592,18.897306,17.288692,15.683984,14.07537,13.481901,12.888432,12.298867,11.705398,11.111929,1.4016805,1.4251068,1.4485333,1.475864,1.4992905,1.5266213,1.5734742,1.620327,1.6671798,1.7140326,1.7608855,1.8467822,1.9287747,2.0107672,2.0927596,2.174752,2.2294137,2.2840753,2.338737,2.3933985,2.4480603,2.455869,2.4597735,2.463678,2.4714866,2.475391,2.4090161,2.338737,2.2723622,2.2059872,2.135708,3.7326086,5.3256044,6.9225054,8.519405,10.112402,8.968412,7.8283267,6.6843367,5.5442514,4.4002614,3.7287042,3.0532427,2.3816853,1.7101282,1.038571,0.95657855,0.8784905,0.79649806,0.71841,0.63641757,0.61689556,0.59737355,0.57785153,0.5583295,0.5388075,0.4997635,0.46071947,0.42557985,0.38653582,0.3513962,0.30844778,0.26940376,0.23035973,0.19131571,0.14836729,0.13274968,0.113227665,0.09761006,0.078088045,0.062470436,0.07027924,0.078088045,0.08589685,0.093705654,0.10151446,0.113227665,0.12884527,0.14446288,0.16008049,0.1756981,0.1717937,0.1639849,0.16008049,0.15617609,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1796025,0.359205,0.5388075,0.71841,0.9019169,0.74574083,0.59346914,0.44119745,0.28892577,0.13665408,0.27721256,0.41777104,0.5583295,0.698888,0.8394465,0.9019169,0.96829176,1.0307622,1.097137,1.1635119,1.175225,1.1869383,1.1986516,1.2142692,1.2259823,1.358732,1.4914817,1.6242313,1.7530766,1.8858263,1.8467822,1.8077383,1.7686942,1.7257458,1.6867018,1.6632754,1.6437533,1.620327,1.5969005,1.5734742,1.6281357,1.6867018,1.7413634,1.796025,1.8506867,1.9404879,2.0302892,2.1200905,2.2098918,2.2996929,2.135708,1.9756275,1.8116426,1.6515622,1.4875772,2.05762,2.6276627,3.1977055,3.767748,4.337791,4.454923,4.572055,4.689187,4.806319,4.9234514,4.8961205,4.8687897,4.841459,4.814128,4.786797,4.3612175,3.9356375,3.513962,3.0883822,2.6628022,2.690133,2.717464,2.7447948,2.7721257,2.7994564,2.7447948,2.690133,2.6354716,2.5808098,2.5261483,3.1977055,3.8692627,4.5408196,5.2162814,5.8878384,6.2587566,6.6257706,6.996689,7.367607,7.7385254,8.609207,9.475985,10.346666,11.217348,12.08803,11.912332,11.736633,11.560935,11.389141,11.213444,10.459893,9.706344,8.956698,8.203149,7.4495993,7.168483,6.883461,6.602344,6.321227,6.036206,6.883461,7.7307167,8.581876,9.4291315,10.276386,10.940135,11.603884,12.271536,12.935285,13.599033,13.673217,13.743496,13.817679,13.891863,13.962143,13.118792,12.2793455,11.435994,10.592644,9.749292,11.506273,13.263254,15.024139,16.78112,18.538101,17.975868,17.413633,16.8514,16.289165,15.726933,14.9109125,14.0948925,13.2788725,12.466757,11.650736,13.325725,15.000713,16.675701,18.35069,20.025679,21.00178,21.981785,22.957886,23.933987,24.91399,25.398136,25.886187,26.374237,26.862288,27.350338,28.650503,29.95067,31.250835,32.551003,33.851166,36.959072,40.063072,43.170975,46.27888,49.386784,53.708958,58.03113,62.353306,66.67938,71.00156,68.93613,66.8746,64.81308,62.751553,60.686123,56.258533,51.827034,47.39554,42.967945,38.53645,33.616905,28.693453,23.77,18.84655,13.923099,14.204215,14.4853325,14.766449,15.043662,15.324779,15.6098,15.894821,16.179844,16.464865,16.749886,24.816381,32.882877,40.953274,49.01977,57.086266,49.437542,41.78882,34.13619,26.487465,18.838741,16.30869,13.78254,11.256392,8.726339,6.2001905,7.0708723,7.941554,8.8083315,9.679013,10.549695,11.283723,12.013845,12.747873,13.481901,14.212025,15.746454,17.27698,18.81141,20.341936,21.876366,23.211672,24.543072,25.878378,27.213684,28.548988,29.903816,31.25474,32.605663,33.96049,35.311413,35.22942,35.143524,35.05763,34.97173,34.885834,32.285503,29.689075,27.088743,24.48841,21.888079,21.903696,21.919313,21.931028,21.946646,21.962263,19.6001,17.237936,14.875772,12.513609,10.151445,8.843472,7.535496,6.2275214,4.919547,3.611572,5.2162814,6.8209906,8.4257,10.034314,11.639023,10.131924,8.628729,7.1216297,5.618435,4.1113358,3.39683,2.6823244,1.9678187,1.2533131,0.5388075,1.7413634,2.9439192,4.1464753,5.349031,6.551587,5.5832953,4.618908,3.6545205,2.690133,1.7257458,1.8233559,1.9209659,2.018576,2.1161861,2.2137961,2.2918842,2.3738766,2.4519646,2.533957,2.612045,2.3192148,2.0224805,1.7257458,1.4329157,1.1361811,1.3938715,1.6515622,1.9092526,2.1669433,2.4246337,2.5495746,2.6745155,2.7994564,2.9243972,3.049338,3.1118085,3.1703746,3.2289407,3.2914112,3.349977,3.5295796,3.7091823,3.8887846,4.068387,4.251894,4.271416,4.290938,4.31046,4.3299823,4.349504,4.9468775,5.5442514,6.141625,6.7389984,7.336372,6.996689,6.657006,6.3173227,5.9776397,5.6379566,5.7707067,5.903456,6.036206,6.168956,6.3017054,6.239235,6.180669,6.1181984,6.0596323,6.001066,6.028397,6.055728,6.083059,6.1103897,6.13772,5.758993,5.3841705,5.0054436,4.6267166,4.251894,4.11524,3.978586,3.8458362,3.7091823,3.5764325,7.7541428,11.927949,16.109564,20.28337,24.46108,24.199486,23.937891,23.676296,23.410795,23.1492,21.173573,19.194042,17.218414,15.238882,13.263254,14.883581,16.503908,18.124235,19.740658,21.360985,21.657719,21.95055,22.247284,22.544018,22.83685,21.763138,20.693333,19.619621,18.54591,17.476105,16.812357,16.148607,15.488764,14.825015,14.161267,14.126127,14.087084,14.051944,14.012899,13.973856,14.903104,15.828446,16.757694,17.683039,18.612286,20.002253,21.39222,22.782187,24.172153,25.562122,22.1731,18.787983,15.398962,12.013845,8.624825,7.8868923,7.1450562,6.4032197,5.6652875,4.9234514,3.9551594,2.9868677,2.0146716,1.0463798,0.07418364,0.078088045,0.08589685,0.08980125,0.093705654,0.10151446,0.28111696,0.46071947,0.64032197,0.8199245,0.999527,1.0112402,1.0190489,1.0307622,1.038571,1.0502841,1.2259823,1.4016805,1.5734742,1.7491722,1.9248703,2.1474214,2.3699722,2.592523,2.815074,3.0376248,3.6584249,4.279225,4.8961205,5.5169206,6.13772,5.989353,5.8370814,5.688714,5.5364423,5.388075,5.056201,4.728231,4.396357,4.068387,3.736513,5.2201858,6.703859,8.183627,9.6673,11.150972,12.220779,13.29449,14.3682,15.438006,16.511717,15.57466,14.637604,13.700547,12.763491,11.826434,12.568271,13.310107,14.051944,14.79378,15.535617,15.449719,15.363823,15.274021,15.188125,15.098324,14.360392,13.618555,12.880623,12.138786,11.400854,11.381332,11.361811,11.338385,11.318862,11.29934,10.975275,10.651209,10.323239,9.999174,9.675109,9.932799,10.19049,10.44818,10.705871,10.963562,11.186112,11.412568,11.639023,11.861574,12.08803,13.282777,14.477524,15.672271,16.867018,18.061766,17.901684,17.7377,17.573715,17.413633,17.24965,17.530766,17.815788,18.096905,18.378021,18.663042,17.597141,16.531239,15.469242,14.40334,13.337439,12.595602,11.85767,11.115833,10.377901,9.636065,9.671205,9.706344,9.741484,9.776623,9.811763,11.435994,13.06413,14.688361,16.312593,17.936825,17.929016,17.921206,17.913397,17.905588,17.901684,17.511244,17.120804,16.730364,16.339924,15.949483,17.136421,18.32336,19.514202,20.701141,21.888079,22.454218,23.01645,23.58259,24.148727,24.710962,23.859802,23.008642,22.153578,21.302418,20.45126,21.048632,21.64991,22.251188,22.848562,23.44984,21.681147,19.916355,18.147661,16.378967,14.614178,13.766922,12.923572,12.076316,11.232965,10.38571,1.3860629,1.4133936,1.43682,1.4641509,1.4875772,1.5110037,1.5656652,1.6242313,1.678893,1.7335546,1.7882162,1.8741131,1.9561055,2.0420024,2.1278992,2.2137961,2.2762666,2.3426414,2.4090161,2.4714866,2.5378613,2.541766,2.541766,2.5456703,2.5456703,2.5495746,2.4597735,2.3699722,2.280171,2.1903696,2.1005683,3.873167,5.645766,7.4183645,9.190963,10.963562,9.546264,8.13287,6.715572,5.3021784,3.8887846,3.3070288,2.7291772,2.1474214,1.5656652,0.9878138,0.9097257,0.8316377,0.75354964,0.679366,0.60127795,0.58956474,0.58175594,0.5700427,0.5583295,0.5505207,0.5114767,0.47633708,0.43729305,0.39824903,0.3631094,0.31625658,0.27330816,0.22645533,0.1835069,0.13665408,0.12103647,0.10932326,0.093705654,0.078088045,0.062470436,0.07418364,0.08199245,0.093705654,0.10151446,0.113227665,0.13274968,0.15227169,0.1717937,0.19131571,0.21083772,0.19912452,0.1835069,0.1678893,0.15227169,0.13665408,0.10932326,0.08199245,0.05466163,0.027330816,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23816854,0.48024148,0.71841,0.96048295,1.1986516,0.9917182,0.78478485,0.57785153,0.3709182,0.1639849,0.24597734,0.3279698,0.40996224,0.49195468,0.57394713,0.58175594,0.58956474,0.59737355,0.60518235,0.61299115,0.62470436,0.63641757,0.6481308,0.6637484,0.6754616,0.8355421,0.9956226,1.1557031,1.3157835,1.475864,1.3938715,1.3118792,1.2259823,1.1439898,1.0619974,1.0463798,1.0268579,1.0112402,0.9917182,0.97610056,1.1283722,1.2806439,1.4329157,1.5851873,1.737459,1.7218413,1.7023194,1.6867018,1.6671798,1.6515622,1.6008049,1.5500476,1.4992905,1.4485333,1.4016805,1.9209659,2.4441557,2.9673457,3.4905357,4.0137253,4.290938,4.5681505,4.845363,5.1225758,5.3997884,5.267039,5.134289,5.001539,4.8687897,4.73604,4.3260775,3.912211,3.4983444,3.0883822,2.6745155,2.7057507,2.7408905,2.7721257,2.803361,2.8385005,2.7330816,2.631567,2.5300527,2.4285383,2.3231194,3.1781836,4.0332475,4.8883114,5.743376,6.5984397,6.8209906,7.043542,7.266093,7.4886436,7.7111945,8.324185,8.933272,9.542359,10.151445,10.764437,10.748819,10.737106,10.725393,10.71368,10.698062,9.991365,9.284669,8.577971,7.871275,7.1606736,6.8756523,6.590631,6.3056097,6.0205884,5.735567,6.5672045,7.3988423,8.226576,9.058213,9.885946,10.721489,11.553126,12.384764,13.216402,14.051944,13.88015,13.708356,13.540467,13.368673,13.200784,12.111456,11.018223,9.928895,8.839567,7.7502384,9.897659,12.045081,14.192502,16.339924,18.487345,17.886066,17.288692,16.687416,16.086138,15.488764,14.668839,13.848915,13.028991,12.209065,11.389141,13.860628,16.33602,18.81141,21.2868,23.762192,24.343948,24.925705,25.511364,26.09312,26.674877,26.862288,27.049698,27.23711,27.424522,27.611933,28.763731,29.911625,31.063425,32.21132,33.363117,36.64672,39.934227,43.217827,46.50143,49.788937,54.478127,59.171215,63.864307,68.557396,73.25049,71.00156,68.74872,66.49978,64.25085,62.001907,56.80905,51.620102,46.431152,41.238297,36.049347,32.020004,27.99066,23.961317,19.92807,15.8987255,16.277452,16.65618,17.031002,17.409729,17.788456,17.093473,16.398489,15.7035055,15.008522,14.313539,25.300526,36.29142,47.28231,58.273205,69.2641,59.987236,50.71428,41.43742,32.16056,22.887606,19.318983,15.746454,12.177831,8.609207,5.036679,6.547683,8.058686,9.565785,11.076789,12.587793,13.384291,14.180789,14.981192,15.77769,16.574188,18.374117,20.170141,21.966167,23.766096,25.562122,26.667067,27.772013,28.876959,29.981905,31.086851,32.695465,34.304077,35.908787,37.517403,39.126015,39.008884,38.89175,38.770714,38.653584,38.53645,35.549583,32.562714,29.575848,26.58898,23.598207,22.481548,21.36489,20.24823,19.13157,18.011007,15.723028,13.438952,11.150972,8.862993,6.575013,5.688714,4.806319,3.9200199,3.0337205,2.1513257,3.0141985,3.8809757,4.743849,5.610626,6.473499,5.6730967,4.8687897,4.068387,3.2640803,2.463678,2.0420024,1.6242313,1.2025559,0.78088045,0.3631094,2.018576,3.677947,5.3334136,6.9927845,8.648251,7.37932,6.1103897,4.841459,3.5686235,2.2996929,2.3035975,2.3114061,2.3153105,2.3192148,2.3231194,2.338737,2.3543546,2.3699722,2.3855898,2.4012074,2.1786566,1.9561055,1.7335546,1.5110037,1.2884527,1.4602464,1.6320401,1.8038338,1.9756275,2.1513257,2.3114061,2.475391,2.639376,2.7994564,2.9634414,2.9165885,2.87364,2.8267872,2.7838387,2.736986,2.9165885,3.0922866,3.2718892,3.4475873,3.6232853,3.7208953,3.8185053,3.9161155,4.0137253,4.1113358,4.630621,5.1460023,5.6652875,6.180669,6.699954,6.4188375,6.133816,5.852699,5.571582,5.2865605,5.270943,5.2592297,5.2436123,5.2279944,5.212377,5.1460023,5.0757227,5.009348,4.942973,4.8765984,5.056201,5.239708,5.423215,5.606722,5.786324,5.4310236,5.0718184,4.716518,4.357313,3.998108,3.8458362,3.68966,3.533484,3.3812122,3.2250361,7.309041,11.389141,15.473146,19.553246,23.63725,22.411268,21.189192,19.96321,18.737226,17.511244,16.578093,15.648844,14.7156925,13.78254,12.849388,14.621986,16.394585,18.167183,19.939783,21.712381,21.895887,22.0833,22.266806,22.454218,22.637724,21.583536,20.529346,19.471254,18.417065,17.362877,16.800642,16.238409,15.676175,15.113941,14.551707,15.113941,15.676175,16.238409,16.800642,17.362877,16.10566,14.852346,13.599033,12.341816,11.088503,15.559043,20.025679,24.49622,28.96676,33.4373,28.537275,23.63725,18.737226,13.837202,8.937177,8.292951,7.648724,7.000593,6.356367,5.7121406,4.575959,3.4436827,2.3075018,1.1713207,0.039044023,0.039044023,0.042948425,0.046852827,0.046852827,0.05075723,0.14055848,0.23035973,0.32016098,0.40996224,0.4997635,0.5036679,0.5114767,0.5153811,0.5192855,0.5231899,0.61299115,0.698888,0.78868926,0.8745861,0.96438736,1.0815194,1.1986516,1.3157835,1.4329157,1.5500476,1.8584955,2.1708477,2.4792955,2.7916477,3.1000953,3.0259118,2.951728,2.87364,2.7994564,2.7252727,2.6081407,2.494913,2.3816853,2.2645533,2.1513257,3.697469,5.2436123,6.79366,8.339804,9.885946,11.256392,12.622932,13.989473,15.356014,16.72646,15.773785,14.825015,13.8762455,12.923572,11.974802,13.1266,14.278399,15.434102,16.585901,17.7377,17.624472,17.511244,17.40192,17.288692,17.175465,16.140799,15.110037,14.079274,13.044608,12.013845,11.963089,11.916236,11.869383,11.82253,11.775677,11.713207,11.650736,11.588266,11.525795,11.4633255,11.82253,12.181735,12.54094,12.90405,13.263254,13.438952,13.610746,13.786445,13.962143,14.13784,14.9109125,15.683984,16.453152,17.226223,17.999294,17.800169,17.601046,17.40192,17.198893,16.999767,16.710842,16.421915,16.129086,15.84016,15.551234,14.629795,13.708356,12.790822,11.869383,10.951848,10.292005,9.636065,8.976221,8.320281,7.6643414,7.8556576,8.046973,8.238289,8.433509,8.624825,10.237343,11.849861,13.462379,15.074897,16.687416,16.640562,16.59371,16.546856,16.4961,16.449247,16.254026,16.058807,15.863586,15.668366,15.473146,16.69913,17.92511,19.151093,20.37317,21.599154,22.344894,23.090635,23.836376,24.578213,25.323954,24.6563,23.984743,23.313187,22.645533,21.973976,22.53621,23.098444,23.660677,24.226816,24.78905,22.860275,20.931501,19.00663,17.077856,15.14908,14.051944,12.954806,11.85767,10.760532,9.663396,1.3743496,1.4016805,1.4251068,1.4485333,1.475864,1.4992905,1.5617609,1.6242313,1.6867018,1.7491722,1.8116426,1.901444,1.9873407,2.0732377,2.1630387,2.2489357,2.3231194,2.4012074,2.475391,2.5495746,2.6237583,2.6237583,2.6237583,2.6237583,2.6237583,2.6237583,2.514435,2.4012074,2.2879796,2.174752,2.0615244,4.0137253,5.9620223,7.914223,9.86252,11.810817,10.124115,8.437413,6.7507114,5.0640097,3.3734035,2.8892577,2.4012074,1.9131571,1.4251068,0.93705654,0.8628729,0.78868926,0.7106012,0.63641757,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.5231899,0.48805028,0.44900626,0.41386664,0.37482262,0.3240654,0.27330816,0.22645533,0.1756981,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.14836729,0.1756981,0.19912452,0.22645533,0.24988174,0.22645533,0.19912452,0.1756981,0.14836729,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.30063897,0.60127795,0.9019169,1.1986516,1.4992905,1.2376955,0.97610056,0.7106012,0.44900626,0.18741131,0.21083772,0.23816854,0.26159495,0.28892577,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.31235218,0.4997635,0.6871748,0.8745861,1.0619974,0.93705654,0.81211567,0.6871748,0.5622339,0.43729305,0.42557985,0.41386664,0.39824903,0.38653582,0.37482262,0.62470436,0.8745861,1.1244678,1.3743496,1.6242313,1.4992905,1.3743496,1.2494087,1.1244678,0.999527,1.0619974,1.1244678,1.1869383,1.2494087,1.3118792,1.7882162,2.260649,2.736986,3.213323,3.6857557,4.123049,4.564246,5.001539,5.4388323,5.8761253,5.6379566,5.3997884,5.1616197,4.9234514,4.689187,4.2870336,3.8887846,3.4866312,3.0883822,2.6862288,2.7252727,2.7643168,2.7994564,2.8385005,2.87364,2.7252727,2.5769055,2.4246337,2.2762666,2.1239948,3.1625657,4.2011366,5.2358036,6.2743745,7.3129454,7.387129,7.461313,7.5394006,7.6135845,7.687768,8.039165,8.386656,8.738052,9.089449,9.43694,9.589212,9.737579,9.885946,10.0382185,10.186585,9.526741,8.862993,8.1992445,7.5394006,6.8756523,6.5867267,6.3017054,6.012779,5.7238536,5.4388323,6.250948,7.0630636,7.8751793,8.687295,9.499411,10.498938,11.498465,12.501896,13.501423,14.50095,14.087084,13.673217,13.263254,12.849388,12.439425,11.100216,9.761005,8.4257,7.08649,5.7511845,8.289046,10.823003,13.360865,15.8987255,18.436588,17.800169,17.163752,16.52343,15.8870125,15.250595,14.426766,13.599033,12.775204,11.951375,11.123642,14.399435,17.675228,20.951023,24.226816,27.498705,27.686117,27.873528,28.06094,28.24835,28.435762,28.326439,28.213211,28.099983,27.986755,27.873528,28.873055,29.876486,30.876013,31.87554,32.87507,36.338272,39.801476,43.260777,46.72398,50.187187,55.251198,60.311302,65.37531,70.43932,75.49943,73.06308,70.62673,68.18648,65.75014,63.313786,57.36348,51.41317,45.46286,39.51255,33.56224,30.423103,27.287867,24.148727,21.013493,17.874353,18.35069,18.823124,19.29946,19.775797,20.24823,18.573242,16.898252,15.223265,13.548276,11.873287,25.788576,39.699963,53.611347,67.526634,81.43802,70.536934,59.639744,48.738655,37.837563,26.936472,22.325373,17.714273,13.09927,8.488171,3.873167,6.0244927,8.175818,10.323239,12.4745655,14.625891,15.488764,16.351637,17.210606,18.073479,18.936352,21.00178,23.063305,25.124828,27.186354,29.251781,30.126368,31.000954,31.87554,32.750126,33.624714,35.487114,37.34951,39.21191,41.07431,42.93671,42.788345,42.636074,42.487705,42.339336,42.187065,38.813663,35.436356,32.06295,28.685644,25.31224,23.063305,20.81437,18.56153,16.312593,14.063657,11.849861,9.636065,7.426173,5.212377,2.998581,2.5378613,2.0732377,1.6125181,1.1517987,0.6871748,0.81211567,0.93705654,1.0619974,1.1869383,1.3118792,1.2142692,1.1127546,1.0112402,0.9136301,0.81211567,0.6871748,0.5622339,0.43729305,0.31235218,0.18741131,2.2996929,4.4119744,6.524256,8.636538,10.748819,9.175345,7.601871,6.0244927,4.4510183,2.87364,2.787743,2.7018464,2.612045,2.5261483,2.436347,2.3855898,2.338737,2.2879796,2.2372224,2.1864653,2.0380979,1.8858263,1.737459,1.5890918,1.43682,1.5266213,1.6125181,1.698415,1.7882162,1.8741131,2.0732377,2.2762666,2.475391,2.6745155,2.87364,2.7252727,2.5769055,2.4246337,2.2762666,2.1239948,2.2996929,2.475391,2.6510892,2.8267872,2.998581,3.174279,3.349977,3.5256753,3.7013733,3.873167,4.3143644,4.7516575,5.1889505,5.6262436,6.0635366,5.8370814,5.610626,5.388075,5.1616197,4.939069,4.775084,4.6110992,4.4510183,4.2870336,4.123049,4.0488653,3.9746814,3.900498,3.8263142,3.7482262,4.087909,4.423688,4.7633705,5.099149,5.4388323,5.099149,4.7633705,4.423688,4.087909,3.7482262,3.5764325,3.4007344,3.2250361,3.049338,2.87364,6.8639393,10.850334,14.836729,18.823124,22.813423,20.623053,18.436588,16.250122,14.063657,11.873287,11.986515,12.099743,12.212971,12.326198,12.439425,14.364296,16.289165,18.214037,20.138906,22.063778,22.13796,22.212145,22.286327,22.364416,22.4386,21.400028,20.361458,19.326792,18.28822,17.24965,16.788929,16.324306,15.863586,15.398962,14.938243,16.101755,17.261362,18.424873,19.588387,20.751898,17.31212,13.8762455,10.436467,7.000593,3.5608149,11.111929,18.663042,26.214157,33.761368,41.31248,34.90145,28.486519,22.07549,15.660558,9.249529,8.699008,8.148487,7.601871,7.0513506,6.5008297,5.2006636,3.900498,2.6003318,1.3001659,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.1639849,0.26159495,0.3631094,0.46071947,0.5622339,2.174752,3.78727,5.3997884,7.012306,8.624825,10.2881,11.951375,13.610746,15.274021,16.937298,15.976814,15.012426,14.048039,13.087557,12.123169,13.688834,15.250595,16.812357,18.374117,19.935879,19.799223,19.662569,19.525915,19.389261,19.248703,17.92511,16.601519,15.274021,13.950429,12.626837,12.548749,12.4745655,12.400381,12.326198,12.24811,12.4511385,12.650263,12.849388,13.048512,13.251541,13.712261,14.176885,14.637604,15.098324,15.562947,15.687888,15.812829,15.93777,16.062712,16.187653,16.539047,16.88654,17.237936,17.589333,17.936825,17.698656,17.464392,17.226223,16.988054,16.749886,15.8870125,15.024139,14.161267,13.298394,12.439425,11.66245,10.885473,10.112402,9.339331,8.562354,7.988407,7.4105554,6.8366084,6.262661,5.688714,6.036206,6.387602,6.7389984,7.08649,7.437886,9.0386915,10.639496,12.236397,13.837202,15.438006,15.348206,15.262308,15.176412,15.086611,15.000713,15.000713,15.000713,15.000713,15.000713,15.000713,16.261835,17.526861,18.787983,20.049105,21.314133,22.239475,23.160913,24.086258,25.0116,25.936945,25.448895,24.960844,24.476698,23.988647,23.500597,24.023787,24.55088,25.074072,25.601166,26.124355,24.0355,21.95055,19.861694,17.776743,15.687888,14.336966,12.986042,11.639023,10.2881,8.937177,1.3509232,1.3821584,1.4133936,1.4485333,1.4797685,1.5110037,1.5890918,1.6632754,1.737459,1.8116426,1.8858263,1.9678187,2.0459068,2.1278992,2.2059872,2.2879796,2.3465457,2.4090161,2.4675822,2.5261483,2.5886188,2.612045,2.639376,2.6628022,2.6862288,2.7135596,2.5808098,2.4519646,2.3231194,2.194274,2.0615244,4.0761957,6.086963,8.101635,10.112402,12.123169,10.307622,8.488171,6.6726236,4.853172,3.0376248,2.619854,2.2020829,1.7843118,1.3665408,0.94876975,0.8628729,0.77307165,0.6871748,0.60127795,0.5114767,0.5075723,0.5036679,0.4958591,0.49195468,0.48805028,0.45291066,0.41777104,0.38263142,0.3474918,0.31235218,0.27330816,0.23426414,0.19131571,0.15227169,0.113227665,0.10932326,0.10932326,0.10541886,0.10151446,0.10151446,0.12884527,0.15617609,0.1835069,0.21083772,0.23816854,0.24988174,0.26159495,0.27330816,0.28892577,0.30063897,0.26159495,0.22645533,0.18741131,0.14836729,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.19912452,0.3631094,0.5231899,0.6871748,0.8511597,0.92143893,0.9917182,1.0580931,1.1283722,1.1986516,0.9917182,0.78088045,0.5700427,0.359205,0.14836729,0.1717937,0.19522011,0.21864653,0.23816854,0.26159495,0.26159495,0.25769055,0.25378615,0.25378615,0.24988174,0.23426414,0.21864653,0.20693332,0.19131571,0.1756981,0.30844778,0.44510186,0.58175594,0.7145056,0.8511597,0.74964523,0.6481308,0.5505207,0.44900626,0.3513962,0.339683,0.3318742,0.32016098,0.30844778,0.30063897,0.5309987,0.76135844,0.9917182,1.2181735,1.4485333,1.33921,1.2259823,1.1127546,0.999527,0.8862993,1.0659018,1.2494087,1.4290112,1.6086137,1.7882162,2.194274,2.6042364,3.0102942,3.416352,3.8263142,4.2167544,4.6110992,5.001539,5.395884,5.786324,5.4973984,5.2084727,4.9156423,4.6267166,4.337791,3.9863946,3.638903,3.2875066,2.9361105,2.5886188,2.6081407,2.6276627,2.6471848,2.6667068,2.6862288,2.5378613,2.3855898,2.2372224,2.0888553,1.9365835,3.0610514,4.181615,5.3060827,6.426646,7.551114,7.6252975,7.699481,7.773665,7.8517528,7.9259367,8.078208,8.23048,8.382751,8.535024,8.687295,8.855185,9.023073,9.190963,9.358852,9.526741,9.030883,8.535024,8.039165,7.5433054,7.0513506,6.6843367,6.321227,5.9542136,5.591104,5.22409,5.9776397,6.7311897,7.480835,8.234385,8.987934,9.866425,10.748819,11.62731,12.5058,13.388195,12.712734,12.037272,11.361811,10.686349,10.010887,9.132397,8.253906,7.3715115,6.493021,5.610626,8.152391,10.694158,13.232019,15.773785,18.311647,18.233559,18.151566,18.073479,17.991486,17.913397,16.613232,15.31697,14.020708,12.720543,11.424281,14.383818,17.343355,20.306797,23.266333,26.22587,26.674877,27.123882,27.576794,28.025799,28.474806,28.525562,28.580225,28.630981,28.685644,28.7364,29.919434,31.102468,32.285503,33.468536,34.65157,37.767284,40.882996,44.002613,47.11833,50.237946,54.380516,58.52699,62.673466,66.81603,70.96251,67.4056,63.84869,60.29178,56.730965,53.174053,48.195942,43.213924,38.235813,33.253796,28.27568,25.796385,23.320995,20.8417,18.366308,15.8870125,16.531239,17.17937,17.823597,18.467823,19.11205,17.718178,16.324306,14.92653,13.532659,12.138786,23.984743,35.8307,47.68056,59.526516,71.37638,61.990196,52.60401,43.217827,33.83555,24.449368,20.783133,17.1169,13.446761,9.780528,6.114294,7.9493628,9.788337,11.623405,13.462379,15.3013525,16.168129,17.03881,17.909492,18.780174,19.650856,21.411741,23.168722,24.92961,26.690495,28.45138,29.607082,30.76669,31.922394,33.078094,34.237705,35.752613,37.26752,38.78243,40.297337,41.812244,41.538937,41.26563,40.996223,40.722916,40.449608,38.735577,37.025448,35.311413,33.601284,31.887253,28.810585,25.73782,22.66115,19.588387,16.511717,13.88015,11.248583,8.6131115,5.9815445,3.349977,3.084478,2.8189783,2.5534792,2.2918842,2.0263848,1.9912452,1.9600099,1.9287747,1.893635,1.8623998,1.7765031,1.6906061,1.6086137,1.5227169,1.43682,1.2337911,1.0268579,0.8238289,0.61689556,0.41386664,2.3192148,4.220659,6.126007,8.031356,9.936704,8.628729,7.320754,6.016684,4.7087092,3.4007344,3.2367494,3.06886,2.9048753,2.7408905,2.5769055,2.541766,2.5105307,2.4792955,2.4441557,2.4129205,2.233318,2.0537157,1.8741131,1.6906061,1.5110037,1.5929961,1.6710842,1.7530766,1.8311646,1.9131571,2.0341935,2.1591344,2.280171,2.4012074,2.5261483,2.4792955,2.436347,2.3894942,2.3465457,2.2996929,2.4285383,2.5612879,2.690133,2.8189783,2.951728,3.2094188,3.4632049,3.7208953,3.978586,4.2362766,4.607195,4.9781127,5.349031,5.716045,6.086963,5.6965227,5.3021784,4.911738,4.5173936,4.123049,4.041056,3.959064,3.8770714,3.795079,3.7130866,3.6467118,3.5764325,3.5100577,3.4436827,3.3734035,3.6271896,3.8809757,4.1308575,4.3846436,4.6384296,4.4197836,4.2011366,3.9863946,3.767748,3.5491016,3.49444,3.4397783,3.3851168,3.330455,3.2757936,6.735094,10.194394,13.653695,17.1169,20.5762,18.631807,16.69132,14.746927,12.806439,10.862047,10.9089,10.955752,11.00651,11.053363,11.100216,12.786918,14.473619,16.164225,17.850927,19.537628,19.78751,20.037392,20.287273,20.537155,20.787037,20.15062,19.518106,18.88169,18.249176,17.612759,16.98415,16.351637,15.723028,15.0944195,14.461906,18.299932,22.13796,25.975988,29.814016,33.64814,27.846197,22.04035,16.234505,10.4286585,4.6267166,10.557504,16.48829,22.422981,28.35377,34.28846,29.361105,24.43375,19.506393,14.579038,9.651682,8.878611,8.105539,7.3324676,6.559396,5.786324,4.630621,3.4710135,2.3153105,1.1557031,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.015617609,0.015617609,0.019522011,0.023426414,0.023426414,0.03513962,0.046852827,0.05466163,0.06637484,0.07418364,0.07418364,0.07027924,0.06637484,0.06637484,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.14836729,0.23426414,0.31625658,0.40215343,0.48805028,1.815547,3.1430438,4.4705405,5.7980375,7.125534,8.421796,9.714153,11.010414,12.306676,13.599033,12.822057,12.045081,11.268105,10.491129,9.714153,11.182208,12.654168,14.122223,15.594183,17.062239,17.066143,17.073952,17.077856,17.08176,17.085665,16.008049,14.92653,13.848915,12.767395,11.685876,11.592171,11.498465,11.400854,11.307149,11.213444,11.377428,11.541413,11.709302,11.873287,12.037272,12.591698,13.142218,13.696643,14.247164,14.801589,14.809398,14.813302,14.821111,14.828919,14.836729,15.172507,15.5082855,15.844065,16.175938,16.511717,16.261835,16.008049,15.754263,15.504381,15.250595,14.621986,13.993378,13.368673,12.740065,12.111456,11.545318,10.979179,10.409137,9.8429985,9.276859,8.894228,8.515501,8.136774,7.7541428,7.375416,7.6135845,7.8517528,8.086017,8.324185,8.562354,9.854712,11.147068,12.439425,13.731783,15.024139,15.016331,15.008522,15.000713,14.996809,14.989,14.981192,14.977287,14.973383,14.965574,14.96167,15.965101,16.968533,17.971964,18.97149,19.974922,20.986162,22.001307,23.012547,24.023787,25.03893,24.46889,23.898846,23.328804,22.75876,22.188719,22.938364,23.691914,24.445463,25.199013,25.948658,24.297094,22.645533,20.99397,19.338505,17.686943,16.168129,14.645412,13.1266,11.607788,10.088976,1.3235924,1.3665408,1.4055848,1.4446288,1.4836729,1.5266213,1.6125181,1.698415,1.7882162,1.8741131,1.9639144,2.0341935,2.1083772,2.1786566,2.25284,2.3231194,2.3699722,2.416825,2.4597735,2.5066261,2.5495746,2.6003318,2.6510892,2.7018464,2.7486992,2.7994564,2.6510892,2.5066261,2.358259,2.2098918,2.0615244,4.138666,6.211904,8.289046,10.362284,12.439425,10.491129,8.542832,6.5945354,4.646239,2.7018464,2.3543546,2.0068626,1.6593709,1.3118792,0.96438736,0.8628729,0.76135844,0.6637484,0.5622339,0.46071947,0.45291066,0.44119745,0.43338865,0.42167544,0.41386664,0.37872702,0.3474918,0.31625658,0.28111696,0.24988174,0.21864653,0.19131571,0.16008049,0.12884527,0.10151446,0.10932326,0.113227665,0.12103647,0.12884527,0.13665408,0.1796025,0.22255093,0.26549935,0.30844778,0.3513962,0.3513962,0.3513962,0.3513962,0.3513962,0.3513962,0.30063897,0.24988174,0.19912452,0.14836729,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.39824903,0.7262188,1.0502841,1.3743496,1.698415,1.5383345,1.3782539,1.2181735,1.0580931,0.9019169,0.7418364,0.58566034,0.42557985,0.26940376,0.113227665,0.13274968,0.15227169,0.1717937,0.19131571,0.21083772,0.25769055,0.30063897,0.3474918,0.39434463,0.43729305,0.39434463,0.3513962,0.30844778,0.26940376,0.22645533,0.30844778,0.39044023,0.47243267,0.5544251,0.63641757,0.5622339,0.48805028,0.41386664,0.3357786,0.26159495,0.25378615,0.24597734,0.23816854,0.23426414,0.22645533,0.43338865,0.6442264,0.8550641,1.0659018,1.2767396,1.175225,1.0737107,0.97610056,0.8745861,0.77307165,1.0737107,1.3704453,1.6671798,1.9639144,2.260649,2.6042364,2.9439192,3.2836022,3.6232853,3.9629683,4.31046,4.657952,5.0054436,5.3529353,5.700427,5.35684,5.0132523,4.6735697,4.3299823,3.9863946,3.6857557,3.3890212,3.0883822,2.787743,2.4871042,2.4910088,2.4910088,2.494913,2.4988174,2.4988174,2.35045,2.1981785,2.0498111,1.901444,1.7491722,2.9556324,4.165997,5.3724575,6.578918,7.7892823,7.8634663,7.9376497,8.011833,8.086017,8.164105,8.117252,8.074304,8.027451,7.9805984,7.9376497,8.121157,8.308568,8.492075,8.675582,8.862993,8.535024,8.207053,7.8790836,7.551114,7.223144,6.7819467,6.3407493,5.8956475,5.45445,5.0132523,5.704332,6.3993154,7.0903945,7.7814736,8.476458,9.2339115,9.99527,10.756628,11.514082,12.27544,11.338385,10.401327,9.464272,8.52331,7.5862536,7.164578,6.7429028,6.321227,5.8956475,5.473972,8.015738,10.561408,13.103174,15.644939,18.186707,18.666946,19.143284,19.619621,20.095959,20.5762,18.8036,17.034906,15.266212,13.493614,11.72492,14.3682,17.015385,19.658665,22.305851,24.949131,25.663635,26.374237,27.088743,27.799343,28.51385,28.728592,28.947239,29.165884,29.380627,29.599274,30.965815,32.32845,33.694992,35.06153,36.424168,39.196293,41.96842,44.74445,47.516575,50.2887,53.513737,56.74268,59.97162,63.196655,66.4256,61.748123,57.07065,52.393173,47.7157,43.038227,39.028404,35.018585,31.008762,26.998941,22.98912,21.169668,19.354122,17.53467,15.719124,13.899672,14.7156925,15.531713,16.343828,17.159847,17.975868,16.85921,15.746454,14.629795,13.513136,12.400381,22.18091,31.965342,41.74587,51.5303,61.31083,53.44346,45.57218,37.70091,29.833538,21.962263,19.240894,16.519526,13.794253,11.072885,8.351517,9.874233,11.400854,12.923572,14.450192,15.976814,16.8514,17.72989,18.608381,19.486872,20.361458,21.821705,23.278046,24.734388,26.190731,27.650976,29.091702,30.52852,31.969246,33.40997,34.850693,36.018112,37.185528,38.352943,39.52036,40.687775,40.29343,39.899086,39.50084,39.10649,38.712147,38.661392,38.610634,38.56378,38.513023,38.462265,34.561768,30.66127,26.760773,22.86418,18.963682,15.9104395,12.857197,9.803954,6.7507114,3.7013733,3.631094,3.5647192,3.4983444,3.4280653,3.3616903,3.174279,2.9829633,2.7916477,2.6042364,2.4129205,2.3426414,2.2723622,2.2020829,2.1318035,2.0615244,1.7765031,1.4914817,1.2064602,0.92143893,0.63641757,2.3348327,4.0332475,5.7316628,7.426173,9.124588,8.086017,7.043542,6.0049706,4.9663997,3.9239242,3.6818514,3.4397783,3.1977055,2.9556324,2.7135596,2.697942,2.6823244,2.6667068,2.6510892,2.639376,2.4285383,2.2177005,2.0068626,1.796025,1.5890918,1.6593709,1.7335546,1.8038338,1.8780174,1.9482968,1.9951496,2.0380979,2.084951,2.1318035,2.174752,2.233318,2.2957885,2.3543546,2.416825,2.475391,2.5612879,2.6432803,2.7291772,2.815074,2.900971,3.240654,3.5803368,3.9200199,4.2597027,4.5993857,4.903929,5.2045684,5.5091114,5.8097506,6.114294,5.55206,4.9937305,4.4314966,3.873167,3.310933,3.310933,3.3070288,3.3031244,3.3031244,3.2992198,3.240654,3.1781836,3.1196175,3.0610514,2.998581,3.1664703,3.3343596,3.5022488,3.6701381,3.8380275,3.7404175,3.6428072,3.5451972,3.4475873,3.349977,3.416352,3.4788225,3.5451972,3.611572,3.6740425,6.606249,9.538455,12.470661,15.406772,18.338978,16.640562,14.942147,13.243732,11.549222,9.850807,9.8312845,9.815667,9.796145,9.780528,9.761005,11.213444,12.661977,14.114414,15.562947,17.01148,17.437061,17.86264,18.28822,18.7138,19.13938,18.905115,18.67085,18.440493,18.206228,17.975868,17.17937,16.378967,15.582469,14.785972,13.985569,20.502016,27.010654,33.527103,40.03574,46.548283,38.37637,30.204456,22.032541,13.860628,5.688714,10.003078,14.317443,18.631807,22.946173,27.260536,23.820759,20.377075,16.933393,13.493614,10.049932,9.054309,8.058686,7.0630636,6.0713453,5.0757227,4.0605783,3.0454338,2.0302892,1.0151446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.031235218,0.03513962,0.039044023,0.046852827,0.05075723,0.058566034,0.06637484,0.07418364,0.078088045,0.08589685,0.08199245,0.078088045,0.07418364,0.06637484,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.13274968,0.20302892,0.27330816,0.3435874,0.41386664,1.456342,2.4988174,3.541293,4.5837684,5.6262436,6.551587,7.480835,8.406178,9.335425,10.260769,9.671205,9.077735,8.484266,7.890797,7.3012323,8.679486,10.053836,11.43209,12.810344,14.188598,14.33306,14.481428,14.629795,14.778163,14.92653,14.090988,13.2554455,12.419904,11.584361,10.748819,10.6355915,10.518459,10.405232,10.2881,10.174872,10.303718,10.436467,10.565312,10.694158,10.826907,11.46723,12.111456,12.751778,13.396004,14.036326,13.927003,13.817679,13.708356,13.599033,13.4858055,13.805966,14.126127,14.446288,14.766449,15.086611,14.821111,14.551707,14.286208,14.016804,13.751305,13.35696,12.96652,12.572175,12.181735,11.787391,11.428185,11.06898,10.705871,10.346666,9.987461,9.803954,9.616543,9.433036,9.245625,9.062118,9.187058,9.311999,9.43694,9.561881,9.686822,10.670732,11.6585455,12.642454,13.626364,14.614178,14.684457,14.75864,14.828919,14.903104,14.973383,14.965574,14.95386,14.946052,14.934339,14.92653,15.668366,16.410202,17.152039,17.893875,18.635712,19.736753,20.837795,21.938837,23.035973,24.137014,23.48498,22.832945,22.18091,21.528873,20.876839,21.856844,22.83685,23.816854,24.796858,25.776863,24.558691,23.340517,22.122343,20.90417,19.685997,17.999294,16.30869,14.618082,12.927476,11.23687,1.3001659,1.3470187,1.3938715,1.4407244,1.4914817,1.5383345,1.6359446,1.737459,1.8389735,1.9365835,2.0380979,2.1005683,2.1669433,2.233318,2.2957885,2.3621633,2.3933985,2.4207294,2.4519646,2.4831998,2.514435,2.5886188,2.6628022,2.736986,2.8111696,2.8892577,2.7213683,2.5573835,2.3933985,2.2294137,2.0615244,4.2011366,6.336845,8.476458,10.612165,12.751778,10.670732,8.59359,6.5164475,4.4393053,2.3621633,2.084951,1.8077383,1.5305257,1.2533131,0.97610056,0.8628729,0.74964523,0.63641757,0.5231899,0.41386664,0.39824903,0.38263142,0.3670138,0.3513962,0.3357786,0.30844778,0.27721256,0.24597734,0.21864653,0.18741131,0.1678893,0.14836729,0.12884527,0.10932326,0.08589685,0.10541886,0.12103647,0.14055848,0.15617609,0.1756981,0.23426414,0.28892577,0.3474918,0.40605783,0.46071947,0.44900626,0.43729305,0.42557985,0.41386664,0.39824903,0.3357786,0.27330816,0.21083772,0.14836729,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.60127795,1.0893283,1.5734742,2.0615244,2.5495746,2.1591344,1.7686942,1.3782539,0.9917182,0.60127795,0.4958591,0.39044023,0.28502136,0.1796025,0.07418364,0.093705654,0.10932326,0.12884527,0.14446288,0.1639849,0.25378615,0.3474918,0.44119745,0.5309987,0.62470436,0.5544251,0.48414588,0.41386664,0.3435874,0.27330816,0.30454338,0.3357786,0.3631094,0.39434463,0.42557985,0.37482262,0.3240654,0.27330816,0.22645533,0.1756981,0.1717937,0.1639849,0.16008049,0.15617609,0.14836729,0.339683,0.5309987,0.71841,0.9097257,1.1010414,1.0112402,0.92534333,0.8394465,0.74964523,0.6637484,1.077615,1.4914817,1.9092526,2.3231194,2.736986,3.0102942,3.2836022,3.5569105,3.8263142,4.0996222,4.4041657,4.704805,5.009348,5.309987,5.610626,5.2162814,4.8219366,4.4275923,4.0332475,3.638903,3.3890212,3.1391394,2.8892577,2.639376,2.3855898,2.3738766,2.358259,2.3426414,2.3270237,2.3114061,2.1630387,2.0107672,1.8623998,1.7140326,1.5617609,2.854118,4.1464753,5.4388323,6.7311897,8.023546,8.101635,8.175818,8.250002,8.324185,8.398369,8.156297,7.914223,7.6721506,7.4300776,7.1880045,7.3910336,7.5940623,7.793187,7.996216,8.1992445,8.039165,7.8790836,7.719003,7.558923,7.3988423,6.8795567,6.3602715,5.840986,5.3217,4.7985106,5.4310236,6.0635366,6.6960497,7.328563,7.9610763,8.601398,9.24172,9.882042,10.522364,11.162686,9.964035,8.761478,7.562827,6.364176,5.1616197,5.196759,5.2318993,5.267039,5.3021784,5.337318,7.882988,10.4286585,12.974329,15.516094,18.061766,19.096432,20.131098,21.165764,22.204336,23.239002,20.99397,18.752844,16.511717,14.2666855,12.025558,14.356487,16.683512,19.014439,21.345367,23.676296,24.64849,25.624592,26.600693,27.576794,28.548988,28.931622,29.314253,29.696884,30.079515,30.462147,32.00829,33.55834,35.10448,36.650623,38.200672,40.62921,43.053844,45.482384,47.91092,50.335552,52.64696,54.958366,57.26587,59.577274,61.88868,56.09064,50.292606,44.494568,38.69653,32.898495,29.860868,26.81934,23.781713,20.740185,17.698656,16.542952,15.383345,14.227642,13.068034,11.912332,12.89624,13.884054,14.867964,15.851873,16.835783,16.004145,15.168603,14.33306,13.497519,12.661977,20.38098,28.096079,35.815083,43.534084,51.249184,44.89672,38.540356,32.183987,25.831526,19.475159,17.698656,15.918248,14.141745,12.365242,10.588739,11.799104,13.013372,14.223738,15.438006,16.64837,17.53467,18.420969,19.303364,20.189665,21.075964,22.231667,23.383465,24.539167,25.694872,26.850574,28.572416,30.294256,32.016098,33.741844,35.463684,36.28361,37.103535,37.92346,38.743385,39.56331,39.04402,38.52864,38.009357,37.493977,36.97469,38.587208,40.199726,41.812244,43.424763,45.03728,40.312954,35.588627,30.8643,26.136068,21.411741,17.94073,14.465811,10.994797,7.523783,4.0488653,4.181615,4.31046,4.4393053,4.5681505,4.7009,4.3534083,4.0059166,3.6584249,3.310933,2.9634414,2.9087796,2.854118,2.7994564,2.7408905,2.6862288,2.3231194,1.9561055,1.5929961,1.2259823,0.8628729,2.3543546,3.8419318,5.3334136,6.8209906,8.312472,7.5394006,6.7663293,5.9932575,5.22409,4.4510183,4.1308575,3.8106966,3.4905357,3.1703746,2.8502135,2.854118,2.854118,2.8580225,2.8619268,2.8619268,2.6237583,2.3816853,2.1435168,1.901444,1.6632754,1.7257458,1.7921207,1.8584955,1.9209659,1.9873407,1.9561055,1.9209659,1.8897307,1.8584955,1.8233559,1.9912452,2.15523,2.3192148,2.4831998,2.6510892,2.690133,2.7291772,2.7682211,2.8111696,2.8502135,3.2718892,3.6935644,4.1191444,4.5408196,4.9624953,5.196759,5.4310236,5.6691923,5.903456,6.13772,5.4115014,4.6813784,3.9551594,3.2289407,2.4988174,2.5769055,2.6549935,2.7330816,2.8111696,2.8892577,2.8345962,2.7838387,2.7291772,2.67842,2.6237583,2.7057507,2.7916477,2.87364,2.9556324,3.0376248,3.0610514,3.0805733,3.1039999,3.1274261,3.1508527,3.3343596,3.521771,3.7052777,3.8887846,4.0761957,6.481308,8.886419,11.291532,13.696643,16.101755,14.649317,13.196879,11.740538,10.2881,8.835662,8.75367,8.671678,8.589685,8.507692,8.4257,9.636065,10.850334,12.0606985,13.274967,14.489237,15.086611,15.687888,16.289165,16.88654,17.487818,17.655706,17.827501,17.999294,18.167183,18.338978,17.370686,16.406298,15.441911,14.477524,13.513136,22.700195,31.887253,41.07431,50.26137,59.44843,48.910446,38.36856,27.83058,17.288692,6.7507114,9.448653,12.146595,14.840633,17.538574,20.236517,18.28041,16.324306,14.364296,12.408191,10.44818,9.2339115,8.015738,6.7975645,5.579391,4.3612175,3.4905357,2.6159496,1.7452679,0.8706817,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.046852827,0.05075723,0.058566034,0.06637484,0.07418364,0.078088045,0.08589685,0.08980125,0.093705654,0.10151446,0.093705654,0.08589685,0.078088045,0.07027924,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.11713207,0.1717937,0.22645533,0.28111696,0.3357786,1.0932326,1.8506867,2.6081407,3.3655949,4.123049,4.6852827,5.2436123,5.805846,6.364176,6.9264097,6.5164475,6.1103897,5.704332,5.2943697,4.8883114,6.17286,7.4574084,8.741957,10.0265045,11.311053,11.603884,11.892809,12.181735,12.470661,12.763491,12.173926,11.584361,10.990892,10.401327,9.811763,9.679013,9.542359,9.405705,9.272955,9.136301,9.2339115,9.327617,9.421323,9.518932,9.612638,10.346666,11.076789,11.810817,12.54094,13.274967,13.048512,12.818152,12.591698,12.365242,12.138786,12.44333,12.747873,13.052417,13.35696,13.661504,13.380386,13.09927,12.814248,12.533132,12.24811,12.091934,11.935758,11.775677,11.619501,11.4633255,11.311053,11.158782,11.00651,10.8542385,10.698062,10.709775,10.721489,10.729298,10.741011,10.748819,10.764437,10.77615,10.787864,10.799577,10.81129,11.490656,12.166118,12.845484,13.520945,14.200311,14.352583,14.504854,14.657126,14.809398,14.96167,14.946052,14.934339,14.918721,14.903104,14.8874855,15.371632,15.851873,16.33602,16.816261,17.300406,18.487345,19.674282,20.861221,22.048159,23.239002,22.50107,21.767042,21.033014,20.298986,19.561056,20.77142,21.97788,23.184341,24.3908,25.601166,24.816381,24.0355,23.250715,22.469835,21.688955,19.826555,17.96806,16.10566,14.247164,12.388668,1.2767396,1.3314011,1.3860629,1.4407244,1.4953861,1.5500476,1.6632754,1.7765031,1.8858263,1.999054,2.1122816,2.1708477,2.2294137,2.2840753,2.3426414,2.4012074,2.416825,2.4285383,2.4441557,2.4597735,2.475391,2.5769055,2.6745155,2.77603,2.87364,2.9751544,2.7916477,2.6081407,2.4285383,2.2450314,2.0615244,4.263607,6.461786,8.663869,10.862047,13.06413,10.8542385,8.648251,6.4383593,4.2323723,2.0263848,1.8194515,1.6086137,1.4016805,1.1947471,0.9878138,0.8628729,0.737932,0.61299115,0.48805028,0.3631094,0.3435874,0.3240654,0.30063897,0.28111696,0.26159495,0.23426414,0.20693332,0.1796025,0.15227169,0.12494087,0.113227665,0.10541886,0.093705654,0.08589685,0.07418364,0.10151446,0.12884527,0.15617609,0.1835069,0.21083772,0.28502136,0.359205,0.42948425,0.5036679,0.57394713,0.5505207,0.5231899,0.4997635,0.47633708,0.44900626,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.80040246,1.4485333,2.1005683,2.7486992,3.4007344,2.7799344,2.1591344,1.5383345,0.92143893,0.30063897,0.24597734,0.19522011,0.14055848,0.08980125,0.039044023,0.05075723,0.06637484,0.08199245,0.09761006,0.113227665,0.25378615,0.39434463,0.5309987,0.6715572,0.81211567,0.7145056,0.61689556,0.5192855,0.42167544,0.3240654,0.30063897,0.28111696,0.25769055,0.23426414,0.21083772,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.08589685,0.08199245,0.078088045,0.078088045,0.07418364,0.24597734,0.41386664,0.58566034,0.75354964,0.92534333,0.8511597,0.77307165,0.698888,0.62470436,0.5505207,1.0815194,1.6164225,2.1474214,2.67842,3.213323,3.416352,3.6232853,3.8263142,4.0332475,4.2362766,4.493967,4.7516575,5.009348,5.267039,5.5247293,5.0757227,4.630621,4.181615,3.736513,3.2875066,3.0883822,2.8892577,2.6862288,2.4871042,2.2879796,2.2567444,2.2216048,2.1903696,2.1591344,2.1239948,1.9756275,1.8233559,1.6749885,1.5266213,1.3743496,2.7526035,4.1308575,5.5091114,6.883461,8.261715,8.335898,8.413987,8.488171,8.562354,8.636538,8.1992445,7.758047,7.3168497,6.8756523,6.4383593,6.657006,6.8756523,7.098203,7.3168497,7.5394006,7.5433054,7.551114,7.558923,7.5667315,7.57454,6.9771667,6.379793,5.7824197,5.185046,4.5876727,5.1616197,5.7316628,6.3056097,6.8756523,7.4495993,7.968885,8.488171,9.01136,9.530646,10.049932,8.58578,7.125534,5.661383,4.2011366,2.736986,3.2289407,3.7208953,4.2167544,4.7087092,5.2006636,7.746334,10.295909,12.841579,15.391153,17.936825,19.52982,21.122816,22.715813,24.30881,25.901804,23.184341,20.470781,17.753317,15.039758,12.326198,14.34087,16.355541,18.370213,20.384884,22.399555,23.63725,24.874947,26.112642,27.350338,28.588034,29.13465,29.681267,30.231787,30.778402,31.32502,33.05467,34.78432,36.51397,38.24362,39.97327,42.05822,44.139267,46.224216,48.305264,50.38631,51.78018,53.174053,54.564022,55.957893,57.351765,50.433163,43.514565,36.595963,29.681267,22.762665,20.693333,18.623999,16.55076,14.481428,12.412095,11.916236,11.416472,10.920613,10.42085,9.924991,11.080693,12.236397,13.388195,14.543899,15.699601,15.145176,14.590752,14.036326,13.481901,12.923572,18.577147,24.23072,29.884295,35.533966,41.18754,36.34608,31.508526,26.667067,21.82561,16.988054,16.156416,15.320874,14.489237,13.657599,12.825961,13.723974,14.625891,15.523903,16.42582,17.323833,18.217941,19.108145,20.002253,20.89636,21.786564,22.641628,23.492788,24.343948,25.199013,26.05017,28.057035,30.059994,32.066856,34.069813,36.076675,36.54911,37.02154,37.493977,37.966408,38.43884,37.79852,37.158195,36.517876,35.877552,35.237232,38.513023,41.78882,45.060707,48.3365,51.612293,46.060234,40.512077,34.96392,29.411861,23.863707,19.971018,16.07833,12.185639,8.292951,4.4002614,4.728231,5.056201,5.3841705,5.708236,6.036206,5.532538,5.02887,4.521298,4.01763,3.513962,3.4710135,3.4319696,3.3929255,3.3538816,3.310933,2.8658314,2.4207294,1.9756275,1.53443,1.0893283,2.3699722,3.6506162,4.9351645,6.2158084,7.5003567,6.996689,6.4891167,5.985449,5.481781,4.9742084,4.575959,4.181615,3.7833657,3.3851168,2.9868677,3.0063896,3.0259118,3.049338,3.06886,3.0883822,2.8189783,2.5456703,2.2762666,2.0068626,1.737459,1.796025,1.8506867,1.9092526,1.9678187,2.0263848,1.9131571,1.8038338,1.6945106,1.5851873,1.475864,1.7452679,2.0146716,2.2840753,2.5534792,2.8267872,2.8189783,2.815074,2.8111696,2.803361,2.7994564,3.3031244,3.8106966,4.3143644,4.8219366,5.3256044,5.493494,5.661383,5.8292727,5.9932575,6.1611466,5.267039,4.3729305,3.4788225,2.5808098,1.6867018,1.8467822,2.0029583,2.1591344,2.3192148,2.475391,2.4285383,2.3855898,2.338737,2.2957885,2.2489357,2.2489357,2.2450314,2.241127,2.241127,2.2372224,2.3816853,2.522244,2.6667068,2.8072653,2.951728,3.2562714,3.5608149,3.8653584,4.169902,4.474445,6.3524623,8.23048,10.108498,11.986515,13.860628,12.654168,11.447707,10.241247,9.030883,7.824422,7.676055,7.531592,7.3832245,7.2348576,7.08649,8.062591,9.0386915,10.010887,10.986988,11.963089,12.73616,13.513136,14.286208,15.063184,15.836256,16.410202,16.98415,17.554192,18.12814,18.698183,17.565907,16.43363,15.3013525,14.169076,13.036799,24.902277,36.76385,48.625427,60.487,72.34857,59.44062,46.53657,33.628616,20.720663,7.812709,8.894228,9.971844,11.053363,12.130978,13.212498,12.740065,12.267632,11.795199,11.322766,10.850334,9.40961,7.968885,6.5281606,5.0913405,3.6506162,2.920493,2.1903696,1.4602464,0.7301232,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.058566034,0.07027924,0.078088045,0.08980125,0.10151446,0.10151446,0.10541886,0.10932326,0.10932326,0.113227665,0.10151446,0.093705654,0.08199245,0.07418364,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.10151446,0.14055848,0.1835069,0.22255093,0.26159495,0.7340276,1.2064602,1.678893,2.1513257,2.6237583,2.8189783,3.0102942,3.2016098,3.39683,3.5881457,3.3655949,3.1430438,2.920493,2.697942,2.475391,3.6662338,4.860981,6.0518236,7.2465706,8.437413,8.870802,9.304191,9.733675,10.167064,10.600452,10.256865,9.909373,9.565785,9.218294,8.874706,8.718531,8.566258,8.410083,8.253906,8.101635,8.160201,8.218767,8.281238,8.339804,8.398369,9.2221985,10.046027,10.865952,11.68978,12.513609,12.166118,11.82253,11.478943,11.131451,10.787864,11.076789,11.365715,11.6585455,11.947471,12.236397,11.939662,11.642927,11.346193,11.0494585,10.748819,10.826907,10.904996,10.983084,11.061172,11.139259,11.193921,11.248583,11.303245,11.357906,11.412568,11.615597,11.82253,12.025558,12.232492,12.439425,12.337912,12.236397,12.138786,12.037272,11.935758,12.306676,12.677594,13.048512,13.415526,13.786445,14.020708,14.251068,14.4853325,14.7156925,14.949956,14.930434,14.9109125,14.89139,14.871868,14.848442,15.070992,15.293544,15.516094,15.738646,15.961197,17.237936,18.51077,19.78751,21.06425,22.337086,21.521065,20.701141,19.88512,19.069101,18.249176,19.685997,21.118912,22.555733,23.988647,25.425468,25.077976,24.730484,24.382992,24.0355,23.68801,21.657719,19.62743,17.597141,15.566852,13.536563,1.2494087,1.3118792,1.3743496,1.43682,1.4992905,1.5617609,1.6867018,1.8116426,1.9365835,2.0615244,2.1864653,2.2372224,2.2879796,2.338737,2.3855898,2.436347,2.436347,2.436347,2.436347,2.436347,2.436347,2.5612879,2.6862288,2.8111696,2.9361105,3.0610514,2.8619268,2.6628022,2.463678,2.260649,2.0615244,4.3260775,6.5867267,8.85128,11.111929,13.376482,11.037745,8.699008,6.364176,4.025439,1.6867018,1.5500476,1.4133936,1.2767396,1.1361811,0.999527,0.8628729,0.7262188,0.58566034,0.44900626,0.31235218,0.28892577,0.26159495,0.23816854,0.21083772,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.10151446,0.13665408,0.1756981,0.21083772,0.24988174,0.3357786,0.42557985,0.5114767,0.60127795,0.6871748,0.6481308,0.61299115,0.57394713,0.5388075,0.4997635,0.41386664,0.3240654,0.23816854,0.14836729,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.999527,1.8116426,2.6237583,3.435874,4.251894,3.4007344,2.5495746,1.698415,0.8511597,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.24988174,0.43729305,0.62470436,0.81211567,0.999527,0.8745861,0.74964523,0.62470436,0.4997635,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14836729,0.30063897,0.44900626,0.60127795,0.74964523,0.6871748,0.62470436,0.5622339,0.4997635,0.43729305,1.0893283,1.737459,2.3855898,3.0376248,3.6857557,3.8263142,3.9629683,4.0996222,4.2362766,4.376835,4.5876727,4.7985106,5.0132523,5.22409,5.4388323,4.939069,4.4393053,3.9356375,3.435874,2.9361105,2.787743,2.639376,2.4871042,2.338737,2.1864653,2.135708,2.0888553,2.0380979,1.9873407,1.9365835,1.7882162,1.6359446,1.4875772,1.33921,1.1869383,2.6510892,4.1113358,5.575486,7.0357327,8.499884,8.574067,8.648251,8.726339,8.800523,8.874706,8.238289,7.601871,6.9615493,6.3251314,5.688714,5.9268827,6.1611466,6.3993154,6.6374836,6.8756523,7.0513506,7.223144,7.3988423,7.57454,7.7502384,7.0747766,6.3993154,5.7238536,5.0483923,4.376835,4.8883114,5.3997884,5.911265,6.426646,6.9381227,7.336372,7.7385254,8.136774,8.538928,8.937177,7.211431,5.4856853,3.7638438,2.0380979,0.31235218,1.261122,2.2137961,3.1625657,4.1113358,5.0640097,7.6135845,10.163159,12.712734,15.262308,17.811884,19.96321,22.11063,24.261955,26.41328,28.560703,25.37471,22.188719,18.998821,15.812829,12.626837,14.325252,16.023666,17.725986,19.4244,21.12672,22.62601,24.125301,25.624592,27.123882,28.623173,29.337679,30.048279,30.762785,31.473387,32.187893,34.101048,36.014206,37.92346,39.836617,41.749775,43.487232,45.22469,46.96215,48.699608,50.43707,50.913406,51.385838,51.862175,52.338512,52.810944,44.775684,36.736523,28.701262,20.662096,12.626837,11.525795,10.424754,9.323712,8.226576,7.125534,7.2856145,7.4495993,7.6135845,7.773665,7.9376497,9.261242,10.588739,11.912332,13.235924,14.56342,14.286208,14.012899,13.735687,13.462379,13.189071,16.773312,20.361458,23.949604,27.537748,31.125895,27.799343,24.476698,21.150146,17.823597,14.50095,14.614178,14.723501,14.836729,14.949956,15.063184,15.648844,16.238409,16.82407,17.413633,17.999294,18.90121,19.799223,20.701141,21.599154,22.50107,23.05159,23.598207,24.148727,24.69925,25.24977,27.537748,29.82573,32.11371,34.401688,36.685764,36.810703,36.935646,37.060585,37.18943,37.314373,36.54911,35.78775,35.026394,34.26113,33.49977,38.43884,43.374004,48.313072,53.248238,58.187305,51.811417,45.439434,39.063545,32.687656,26.311768,22.001307,17.686943,13.376482,9.062118,4.7516575,5.2748475,5.7980375,6.3251314,6.8483214,7.375416,6.7116675,6.0518236,5.388075,4.7243266,4.0605783,4.037152,4.0137253,3.9863946,3.9629683,3.9356375,3.4124475,2.8892577,2.3621633,1.8389735,1.3118792,2.3894942,3.4632049,4.5369153,5.610626,6.688241,6.4500723,6.211904,5.9737353,5.735567,5.5013027,5.024966,4.548629,4.0761957,3.5998588,3.1235218,3.1625657,3.2016098,3.2367494,3.2757936,3.310933,3.0141985,2.7135596,2.4129205,2.1122816,1.8116426,1.8623998,1.9131571,1.9639144,2.0107672,2.0615244,1.8741131,1.6867018,1.4992905,1.3118792,1.1244678,1.4992905,1.8741131,2.2489357,2.6237583,2.998581,2.951728,2.900971,2.8502135,2.7994564,2.7486992,3.338264,3.9239242,4.513489,5.099149,5.688714,5.786324,5.8878384,5.989353,6.086963,6.1884775,5.12648,4.0644827,2.998581,1.9365835,0.8745861,1.1127546,1.3509232,1.5890918,1.8233559,2.0615244,2.0263848,1.9873407,1.9482968,1.9131571,1.8741131,1.7882162,1.698415,1.6125181,1.5266213,1.43682,1.698415,1.9639144,2.2255092,2.4871042,2.7486992,3.174279,3.5998588,4.025439,4.4510183,4.8765984,6.223617,7.57454,8.925464,10.276386,11.623405,10.662923,9.698535,8.738052,7.773665,6.813182,6.5984397,6.387602,6.1767645,5.9620223,5.7511845,6.4891167,7.223144,7.9610763,8.699008,9.43694,10.38571,11.338385,12.287154,13.235924,14.188598,15.160794,16.136894,17.112995,18.089096,19.061293,17.761126,16.46096,15.160794,13.860628,12.564366,27.100456,41.636547,56.17654,70.71263,85.24872,69.9747,54.700676,39.42275,24.148727,8.874706,8.335898,7.800996,7.262188,6.7233806,6.1884775,7.1997175,8.210958,9.226103,10.237343,11.248583,9.589212,7.9259367,6.262661,4.5993857,2.9361105,2.35045,1.7608855,1.175225,0.58566034,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.37482262,0.5622339,0.74964523,0.93705654,1.1244678,0.94876975,0.77307165,0.60127795,0.42557985,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,1.1635119,2.260649,3.3616903,4.462732,5.563773,6.13772,6.7116675,7.2856145,7.8634663,8.437413,8.335898,8.238289,8.136774,8.039165,7.9376497,7.7619514,7.5862536,7.4105554,7.238762,7.0630636,7.08649,7.113821,7.137247,7.1606736,7.1880045,8.101635,9.01136,9.924991,10.838621,11.748346,11.287627,10.826907,10.362284,9.901564,9.43694,9.714153,9.987461,10.260769,10.537982,10.81129,10.498938,10.186585,9.874233,9.561881,9.249529,9.561881,9.874233,10.186585,10.498938,10.81129,11.076789,11.338385,11.599979,11.861574,12.123169,12.525322,12.923572,13.325725,13.723974,14.126127,13.911386,13.700547,13.4858055,13.274967,13.06413,13.1266,13.189071,13.251541,13.314012,13.376482,13.688834,14.001186,14.313539,14.625891,14.938243,14.9109125,14.8874855,14.864059,14.836729,14.813302,14.774258,14.739119,14.700074,14.661031,14.625891,15.988527,17.351164,18.7138,20.076437,21.439074,20.537155,19.639143,18.737226,17.839214,16.937298,18.600573,20.263847,21.923218,23.586494,25.24977,25.335667,25.425468,25.511364,25.601166,25.687063,23.488884,21.2868,19.088623,16.88654,14.688361,1.2142692,1.2962615,1.3782539,1.4602464,1.542239,1.6242313,1.7608855,1.893635,2.0302892,2.1669433,2.2996929,2.3153105,2.330928,2.3465457,2.358259,2.3738766,2.366068,2.3543546,2.3465457,2.3348327,2.3231194,2.4675822,2.6081407,2.7526035,2.893162,3.0376248,2.900971,2.7643168,2.6237583,2.4871042,2.35045,4.493967,6.6335793,8.777096,10.920613,13.06413,10.760532,8.456935,6.153338,3.853645,1.5500476,1.4290112,1.3040704,1.183034,1.0580931,0.93705654,0.80040246,0.6637484,0.5231899,0.38653582,0.24988174,0.23816854,0.22645533,0.21083772,0.19912452,0.18741131,0.1717937,0.15227169,0.13665408,0.11713207,0.10151446,0.10151446,0.10541886,0.10932326,0.10932326,0.113227665,0.14055848,0.1678893,0.19522011,0.22255093,0.24988174,0.3318742,0.40996224,0.48805028,0.5700427,0.6481308,0.60908675,0.5700427,0.5309987,0.48805028,0.44900626,0.3709182,0.29673457,0.21864653,0.14055848,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.80040246,1.4485333,2.1005683,2.7486992,3.4007344,2.7213683,2.0380979,1.358732,0.679366,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.15617609,0.19131571,0.22255093,0.25378615,0.28892577,0.39044023,0.49195468,0.59346914,0.698888,0.80040246,0.698888,0.60127795,0.4997635,0.39824903,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.19131571,0.3318742,0.46852827,0.60908675,0.74964523,0.8433509,0.94096094,1.0346665,1.1283722,1.2259823,1.7218413,2.2137961,2.7096553,3.2055142,3.7013733,3.8106966,3.9239242,4.037152,4.1503797,4.263607,4.493967,4.728231,4.958591,5.192855,5.423215,4.9937305,4.560342,4.126953,3.6935644,3.2640803,3.1391394,3.0141985,2.8892577,2.7643168,2.639376,2.5651922,2.4910088,2.4207294,2.3465457,2.2762666,2.1591344,2.0380979,1.9209659,1.8038338,1.6867018,3.049338,4.40807,5.7668023,7.1294384,8.488171,8.4178915,8.347612,8.277332,8.207053,8.136774,7.746334,7.355894,6.969358,6.578918,6.1884775,6.297801,6.407124,6.5164475,6.6257706,6.7389984,6.7624245,6.785851,6.813182,6.8366084,6.8639393,6.387602,5.911265,5.4388323,4.9624953,4.4861584,4.9663997,5.446641,5.9268827,6.407124,6.8873653,7.098203,7.3129454,7.523783,7.7385254,7.9493628,6.473499,5.001539,3.5256753,2.0498111,0.57394713,1.4719596,2.3699722,3.2679846,4.165997,5.0640097,7.617489,10.170968,12.728352,15.281831,17.839214,20.849508,23.863707,26.874,29.888199,32.898495,28.74421,24.586021,20.427834,16.269644,12.111456,14.036326,15.961197,17.886066,19.810938,21.735807,22.99693,24.254147,25.511364,26.768581,28.025799,28.861341,29.696884,30.52852,31.364063,32.199604,34.097145,35.994686,37.892223,39.789764,41.6873,42.761013,43.838627,44.91234,45.98605,47.063663,47.864067,48.668373,49.468777,50.273083,51.073486,43.787872,36.498352,29.212738,21.923218,14.637604,13.196879,11.756155,10.319335,8.878611,7.437886,8.015738,8.597494,9.17925,9.757101,10.338858,10.967466,11.596075,12.228588,12.857197,13.4858055,13.204688,12.923572,12.63855,12.357433,12.076316,14.907008,17.741604,20.572296,23.40689,26.237583,23.71534,21.193096,18.67085,16.148607,13.626364,13.657599,13.688834,13.723974,13.755209,13.786445,14.243259,14.703979,15.160794,15.617609,16.074425,16.906061,17.733795,18.565434,19.393166,20.224804,20.5762,20.931501,21.282896,21.634293,21.98569,23.906654,25.823717,27.740778,29.657839,31.574902,31.71546,31.856018,31.996576,32.133232,32.27379,32.387016,32.500244,32.613472,32.7267,32.83602,37.251904,41.663876,46.07585,50.487827,54.8998,48.605904,42.312008,36.014206,29.72031,23.426414,19.557152,15.6917925,11.82253,7.9532676,4.087909,4.5993857,5.1108627,5.6262436,6.13772,6.649197,6.016684,5.380266,4.743849,4.1113358,3.474918,3.5178664,3.5608149,3.6037633,3.6467118,3.6857557,3.232845,2.77603,2.3231194,1.8663043,1.4133936,2.2372224,3.0610514,3.8887846,4.7126136,5.5364423,5.563773,5.5871997,5.610626,5.6379566,5.661383,5.3138914,4.9624953,4.6110992,4.263607,3.912211,3.8692627,3.8263142,3.7833657,3.7443218,3.7013733,3.4436827,3.1898966,2.9361105,2.67842,2.4246337,2.377781,2.330928,2.2840753,2.233318,2.1864653,2.15523,2.1239948,2.0888553,2.05762,2.0263848,2.3270237,2.631567,2.9322062,3.2367494,3.5373883,3.5608149,3.5842414,3.6037633,3.6271896,3.6506162,4.0801005,4.5095844,4.939069,5.368553,5.801942,5.8956475,5.989353,6.083059,6.180669,6.2743745,5.3334136,4.388548,3.4475873,2.5066261,1.5617609,1.7218413,1.8819219,2.0420024,2.2020829,2.3621633,2.3738766,2.3816853,2.3933985,2.4012074,2.4129205,2.463678,2.5183394,2.5690966,2.6237583,2.6745155,2.639376,2.6003318,2.5612879,2.5261483,2.4871042,3.2367494,3.9824903,4.728231,5.477876,6.223617,7.1841,8.144583,9.105066,10.065549,11.0260315,10.174872,9.323712,8.476458,7.6252975,6.774138,6.7780423,6.7819467,6.7819467,6.785851,6.785851,8.093826,9.397896,10.701966,12.006037,13.314012,13.930907,14.547803,15.164699,15.781594,16.398489,17.335546,18.268698,19.205755,20.138906,21.075964,19.229181,17.378494,15.531713,13.68493,11.838148,25.382519,38.92689,52.47126,66.01954,79.56391,65.38312,51.20233,37.02154,22.840754,8.663869,10.120211,11.576552,13.036799,14.493141,15.949483,15.051471,14.149553,13.251541,12.349625,11.4516115,9.628256,7.8088045,5.989353,4.169902,2.35045,1.8780174,1.4094892,0.94096094,0.46852827,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.11713207,0.14836729,0.1756981,0.20693332,0.23816854,0.23426414,0.22645533,0.22255093,0.21864653,0.21083772,0.1835069,0.15227169,0.12103647,0.093705654,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.08980125,0.11713207,0.14446288,0.1717937,0.19912452,0.3435874,0.48414588,0.62860876,0.76916724,0.9136301,0.76916724,0.62860876,0.48414588,0.3435874,0.19912452,0.1717937,0.14055848,0.10932326,0.078088045,0.05075723,0.92924774,1.8116426,2.690133,3.5686235,4.4510183,4.9156423,5.3841705,5.852699,6.321227,6.785851,6.7311897,6.676528,6.621866,6.5672045,6.5125427,6.3836975,6.2587566,6.1299114,6.001066,5.8761253,5.958118,6.044015,6.1299114,6.2158084,6.3017054,7.008402,7.715099,8.421796,9.128492,9.839094,9.475985,9.112875,8.749765,8.386656,8.023546,8.32809,8.636538,8.941081,9.245625,9.550168,9.284669,9.019169,8.75367,8.488171,8.226576,8.406178,8.589685,8.773191,8.956698,9.136301,9.397896,9.655587,9.917182,10.178777,10.436467,10.819098,11.20173,11.584361,11.966993,12.349625,12.24811,12.150499,12.0489855,11.951375,11.849861,11.970898,12.091934,12.209065,12.330102,12.4511385,12.950902,13.45457,13.958238,14.461906,14.96167,14.89139,14.821111,14.750832,14.6805525,14.614178,14.700074,14.785972,14.875772,14.96167,15.051471,16.421915,17.788456,19.158901,20.529346,21.899792,21.068155,20.236517,19.400974,18.569338,17.7377,18.84655,19.951496,21.060347,22.169195,23.274141,23.527927,23.781713,24.031595,24.285381,24.539167,22.7939,21.048632,19.303364,17.558098,15.812829,1.175225,1.2767396,1.3782539,1.4836729,1.5851873,1.6867018,1.8311646,1.9756275,2.1239948,2.2684577,2.4129205,2.3933985,2.3738766,2.3543546,2.330928,2.3114061,2.2918842,2.2723622,2.25284,2.233318,2.2137961,2.3738766,2.533957,2.6940374,2.854118,3.0141985,2.9361105,2.8619268,2.787743,2.7135596,2.639376,4.661856,6.6843367,8.706817,10.729298,12.751778,10.48332,8.214863,5.9464045,3.6818514,1.4133936,1.3040704,1.1986516,1.0893283,0.98390937,0.8745861,0.737932,0.60127795,0.46071947,0.3240654,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.1756981,0.1678893,0.15617609,0.14836729,0.13665408,0.14055848,0.14836729,0.15227169,0.15617609,0.1639849,0.1796025,0.19912452,0.21474212,0.23426414,0.24988174,0.3240654,0.39434463,0.46852827,0.5388075,0.61299115,0.5700427,0.5270943,0.48414588,0.44119745,0.39824903,0.3318742,0.26549935,0.19912452,0.12884527,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.60127795,1.0893283,1.5734742,2.0615244,2.5495746,2.0380979,1.5305257,1.0190489,0.5114767,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.30063897,0.3553006,0.40605783,0.46071947,0.5114767,0.5309987,0.5466163,0.5661383,0.58175594,0.60127795,0.5231899,0.44900626,0.37482262,0.30063897,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.23035973,0.359205,0.49195468,0.62079996,0.74964523,1.0034313,1.2533131,1.5070993,1.7608855,2.0107672,2.3543546,2.6940374,3.0337205,3.3734035,3.7130866,3.7989833,3.8887846,3.9746814,4.0605783,4.1503797,4.4041657,4.6540475,4.9078336,5.1616197,5.4115014,5.0483923,4.6813784,4.318269,3.951255,3.5881457,3.4866312,3.3890212,3.2875066,3.1859922,3.0883822,2.9907722,2.8970666,2.803361,2.7057507,2.612045,2.5261483,2.4441557,2.358259,2.2723622,2.1864653,3.4436827,4.7009,5.958118,7.2192397,8.476458,8.261715,8.043069,7.8283267,7.6135845,7.3988423,7.2582836,7.113821,6.9732623,6.8287997,6.688241,6.6687193,6.6531014,6.6335793,6.617962,6.5984397,6.473499,6.348558,6.223617,6.098676,5.9737353,5.700427,5.423215,5.1499066,4.8765984,4.5993857,5.0483923,5.493494,5.9425,6.3915067,6.8366084,6.8639393,6.8873653,6.910792,6.9381227,6.9615493,5.735567,4.513489,3.2875066,2.0615244,0.8394465,1.6827974,2.5261483,3.3734035,4.2167544,5.0640097,7.621393,10.182681,12.743969,15.3013525,17.86264,21.735807,25.612879,29.486046,33.363117,37.236286,32.109802,26.983324,21.85294,16.72646,11.599979,13.751305,15.8987255,18.05005,20.201378,22.348799,23.363943,24.379087,25.394232,26.409376,27.424522,28.3811,29.341583,30.29816,31.25474,32.21132,34.09324,35.979065,37.86099,39.742912,41.624832,42.0387,42.44866,42.86253,43.276394,43.686356,44.818634,45.947006,47.07928,48.207653,49.336025,42.800056,36.264088,29.724215,23.188246,16.64837,14.871868,13.091461,11.311053,9.530646,7.7502384,8.745861,9.745388,10.741011,11.740538,12.73616,12.67369,12.607315,12.54094,12.47847,12.412095,12.123169,11.834243,11.541413,11.252487,10.963562,13.040704,15.117846,17.194988,19.27213,21.349272,19.631334,17.909492,16.191557,14.469715,12.751778,12.70102,12.654168,12.607315,12.560462,12.513609,12.841579,13.165645,13.493614,13.821584,14.149553,14.9109125,15.668366,16.429726,17.191084,17.948538,18.104713,18.26089,18.41316,18.569338,18.725513,20.271656,21.821705,23.367847,24.91399,26.464039,26.61631,26.772486,26.928663,27.080935,27.23711,28.224924,29.212738,30.200552,31.188366,32.176178,36.061058,39.949844,43.838627,47.723507,51.612293,45.396484,39.18458,32.968773,26.752964,20.537155,17.112995,13.692739,10.268578,6.8483214,3.4241607,3.9239242,4.423688,4.9234514,5.423215,5.9268827,5.3177958,4.7087092,4.1035266,3.49444,2.8892577,2.998581,3.1079042,3.2172275,3.3265507,3.435874,3.0532427,2.6667068,2.2840753,1.8975395,1.5110037,2.0888553,2.6628022,3.2367494,3.8106966,4.388548,4.6735697,4.9624953,5.251421,5.5364423,5.825368,5.5989127,5.376362,5.1499066,4.9234514,4.7009,4.575959,4.454923,4.3338866,4.2089458,4.087909,3.8770714,3.6662338,3.4593005,3.2484627,3.0376248,2.893162,2.7486992,2.6042364,2.455869,2.3114061,2.436347,2.5573835,2.67842,2.803361,2.9243972,3.154757,3.3851168,3.6154766,3.8458362,4.0761957,4.169902,4.263607,4.3612175,4.454923,4.548629,4.8219366,5.095245,5.368553,5.6418614,5.911265,6.001066,6.0908675,6.180669,6.2743745,6.364176,5.5403466,4.716518,3.8965936,3.0727646,2.2489357,2.330928,2.416825,2.4988174,2.5808098,2.6628022,2.7213683,2.77603,2.8345962,2.893162,2.951728,3.1430438,3.3343596,3.5256753,3.7208953,3.912211,3.5764325,3.2367494,2.900971,2.5612879,2.2255092,3.2953155,4.365122,5.434928,6.504734,7.57454,8.144583,8.714626,9.284669,9.854712,10.424754,9.686822,8.94889,8.210958,7.47693,6.7389984,6.9537406,7.172387,7.3910336,7.605776,7.824422,9.698535,11.568744,13.442857,15.31697,17.18718,17.4722,17.757221,18.042242,18.327265,18.612286,19.506393,20.404406,21.298513,22.192623,23.086731,20.693333,18.296028,15.902631,13.509232,11.111929,23.664581,36.217236,48.76989,61.32254,73.8752,60.78764,47.703987,34.620335,21.536682,8.449126,11.904523,15.356014,18.807507,22.258997,25.714394,22.899319,20.08815,17.273075,14.461906,11.650736,9.671205,7.6955767,5.716045,3.7404175,1.7608855,1.4094892,1.0580931,0.7066968,0.3513962,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.16008049,0.20693332,0.25378615,0.30063897,0.3513962,0.339683,0.3318742,0.32016098,0.30844778,0.30063897,0.25378615,0.20693332,0.15617609,0.10932326,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.093705654,0.12103647,0.15227169,0.1835069,0.21083772,0.30844778,0.40605783,0.5036679,0.60127795,0.698888,0.58956474,0.48024148,0.3709182,0.26159495,0.14836729,0.12884527,0.10541886,0.08199245,0.058566034,0.039044023,0.698888,1.358732,2.018576,2.67842,3.338264,3.697469,4.056674,4.415879,4.7789884,5.138193,5.12648,5.1186714,5.1069584,5.099149,5.087436,5.009348,4.927356,4.8492675,4.7672753,4.689187,4.83365,4.9781127,5.1225758,5.267039,5.4115014,5.9151692,6.4188375,6.918601,7.422269,7.9259367,7.6643414,7.3988423,7.137247,6.8756523,6.6140575,6.9459314,7.28171,7.617489,7.9532676,8.289046,8.070399,7.8517528,7.633106,7.4183645,7.1997175,7.2543793,7.3051367,7.355894,7.4105554,7.461313,7.719003,7.9766936,8.234385,8.492075,8.749765,9.116779,9.479889,9.846903,10.2100115,10.573121,10.588739,10.600452,10.612165,10.6238785,10.6355915,10.815194,10.990892,11.170495,11.346193,11.525795,12.216875,12.911859,13.602938,14.294017,14.989,14.871868,14.75864,14.641508,14.528281,14.411149,14.625891,14.836729,15.051471,15.262308,15.473146,16.8514,18.229654,19.607908,20.986162,22.364416,21.599154,20.83389,20.068628,19.303364,18.538101,19.088623,19.643047,20.19357,20.747993,21.298513,21.716286,22.134056,22.551826,22.969599,23.38737,22.098917,20.80656,19.518106,18.22575,16.937298,1.1361811,1.261122,1.3821584,1.5031948,1.6281357,1.7491722,1.9053483,2.0615244,2.2137961,2.3699722,2.5261483,2.4714866,2.416825,2.358259,2.3035975,2.2489357,2.2216048,2.1903696,2.1591344,2.1318035,2.1005683,2.2762666,2.455869,2.631567,2.8111696,2.9868677,2.9751544,2.9634414,2.951728,2.9361105,2.9243972,4.825841,6.7311897,8.632633,10.534078,12.439425,10.206107,7.9727893,5.7394714,3.506153,1.2767396,1.183034,1.0893283,0.9956226,0.9058213,0.81211567,0.6754616,0.5388075,0.39824903,0.26159495,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.1835069,0.1835069,0.1796025,0.1756981,0.1756981,0.1835069,0.19131571,0.19912452,0.20693332,0.21083772,0.21864653,0.22645533,0.23426414,0.24207294,0.24988174,0.31625658,0.37872702,0.44510186,0.5114767,0.57394713,0.5309987,0.48414588,0.44119745,0.39434463,0.3513962,0.29283017,0.23426414,0.1756981,0.12103647,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.39824903,0.7262188,1.0502841,1.3743496,1.698415,1.358732,1.0190489,0.679366,0.339683,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.44900626,0.5192855,0.59346914,0.6637484,0.737932,0.6715572,0.60127795,0.5349031,0.46852827,0.39824903,0.3513962,0.30063897,0.24988174,0.19912452,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.26940376,0.39044023,0.5114767,0.62860876,0.74964523,1.1596074,1.5695697,1.979532,2.3894942,2.7994564,2.9868677,3.1703746,3.3538816,3.541293,3.7247996,3.78727,3.8497405,3.912211,3.9746814,4.037152,4.31046,4.5837684,4.853172,5.12648,5.3997884,5.1030536,4.806319,4.50568,4.2089458,3.912211,3.8380275,3.7638438,3.6857557,3.611572,3.5373883,3.4202564,3.3031244,3.1859922,3.06886,2.951728,2.8970666,2.8463092,2.7916477,2.7408905,2.6862288,3.8419318,4.997635,6.153338,7.309041,8.460839,8.101635,7.7424297,7.3832245,7.0240197,6.66091,6.7663293,6.871748,6.9771667,7.082586,7.1880045,7.043542,6.899079,6.7507114,6.606249,6.461786,6.1884775,5.911265,5.6379566,5.3607445,5.087436,5.0132523,4.939069,4.860981,4.786797,4.7126136,5.12648,5.5442514,5.958118,6.3719845,6.785851,6.6257706,6.461786,6.3017054,6.13772,5.9737353,5.001539,4.025439,3.049338,2.0732377,1.1010414,1.893635,2.6862288,3.4788225,4.271416,5.0640097,7.629202,10.19049,12.755682,15.320874,17.886066,22.62601,27.362051,32.101994,36.838036,41.574074,35.4793,29.380627,23.28195,17.183275,11.088503,13.462379,15.836256,18.214037,20.587914,22.96179,23.734861,24.507933,25.281004,26.054077,26.823244,27.904762,28.986282,30.063898,31.145416,32.226936,34.09324,35.959545,37.825848,39.696056,41.562363,41.31248,41.0626,40.812717,40.562836,40.312954,41.769295,43.225636,44.685883,46.142227,47.598568,41.812244,36.02592,30.235691,24.449368,18.663042,16.542952,14.422862,12.302772,10.182681,8.062591,9.475985,10.893282,12.306676,13.723974,15.137367,14.376009,13.618555,12.857197,12.095839,11.338385,11.04165,10.741011,10.444276,10.147541,9.850807,11.174399,12.494087,13.817679,15.141272,16.46096,15.543426,14.625891,13.708356,12.790822,11.873287,11.748346,11.619501,11.490656,11.365715,11.23687,11.435994,11.631214,11.8303385,12.025558,12.224684,12.915763,13.606842,14.294017,14.985096,15.676175,15.633226,15.590279,15.54733,15.504381,15.461433,16.640562,17.815788,18.994917,20.174046,21.349272,21.521065,21.688955,21.860748,22.028637,22.200432,24.062832,25.925232,27.78763,29.65003,31.51243,34.874123,38.235813,41.601406,44.963097,48.324787,42.19097,36.05325,29.919434,23.785618,17.651802,14.672744,11.693685,8.718531,5.7394714,2.7643168,3.2484627,3.736513,4.224563,4.7126136,5.2006636,4.618908,4.041056,3.4593005,2.8814487,2.2996929,2.4792955,2.6549935,2.8306916,3.0102942,3.1859922,2.87364,2.5573835,2.241127,1.9287747,1.6125181,1.9365835,2.260649,2.5886188,2.912684,3.2367494,3.78727,4.337791,4.8883114,5.4388323,5.989353,5.8878384,5.786324,5.688714,5.5871997,5.4856853,5.2865605,5.083532,4.8805027,4.677474,4.474445,4.31046,4.1464753,3.978586,3.814601,3.6506162,3.408543,3.1664703,2.9243972,2.67842,2.436347,2.7135596,2.9907722,3.2718892,3.5491016,3.8263142,3.9824903,4.138666,4.298747,4.454923,4.6110992,4.7789884,4.9468775,5.114767,5.282656,5.4505453,5.563773,5.6809053,5.794133,5.911265,6.0244927,6.1103897,6.196286,6.278279,6.364176,6.4500723,5.74728,5.044488,4.3416953,3.638903,2.9361105,2.9439192,2.9478238,2.951728,2.9556324,2.9634414,3.06886,3.174279,3.2757936,3.3812122,3.4866312,3.8185053,4.154284,4.4861584,4.8180323,5.1499066,4.513489,3.873167,3.2367494,2.6003318,1.9639144,3.3538816,4.747753,6.141625,7.531592,8.925464,9.105066,9.284669,9.464272,9.643873,9.823476,9.198771,8.574067,7.9493628,7.3246584,6.699954,7.1333427,7.5667315,7.996216,8.429605,8.862993,11.303245,13.743496,16.183748,18.623999,21.06425,21.013493,20.96664,20.919786,20.872934,20.826082,21.681147,22.53621,23.391273,24.246338,25.101402,22.157482,19.213564,16.273548,13.329629,10.38571,21.946646,33.50758,45.068516,56.62945,68.18648,56.19606,44.209545,32.21522,20.228708,8.238289,13.68493,19.13157,24.582117,30.028757,35.4754,30.751072,26.026745,21.298513,16.574188,11.849861,9.714153,7.578445,5.446641,3.310933,1.175225,0.94096094,0.7066968,0.46852827,0.23426414,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.13665408,0.20302892,0.26940376,0.3318742,0.39824903,0.46071947,0.44900626,0.43338865,0.41777104,0.40215343,0.38653582,0.3240654,0.25769055,0.19131571,0.12884527,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.093705654,0.12884527,0.16008049,0.19131571,0.22645533,0.27721256,0.3318742,0.38263142,0.43338865,0.48805028,0.40996224,0.3318742,0.25378615,0.1756981,0.10151446,0.08589685,0.07027924,0.05466163,0.039044023,0.023426414,0.46462387,0.9058213,1.3431144,1.7843118,2.2255092,2.4792955,2.7291772,2.9829633,3.2367494,3.4866312,3.521771,3.5569105,3.59205,3.6271896,3.6623292,3.631094,3.5959544,3.5647192,3.533484,3.4983444,3.7052777,3.9083066,4.11524,4.318269,4.5252023,4.8219366,5.1186714,5.4193106,5.716045,6.012779,5.8487945,5.688714,5.5247293,5.3607445,5.2006636,5.563773,5.930787,6.2938967,6.66091,7.0240197,6.8561306,6.6843367,6.5164475,6.3446536,6.1767645,6.098676,6.0205884,5.9425,5.8644123,5.786324,6.044015,6.297801,6.551587,6.8092775,7.0630636,7.4105554,7.758047,8.105539,8.453031,8.800523,8.925464,9.050405,9.175345,9.300286,9.425227,9.659492,9.893755,10.131924,10.366188,10.600452,11.482847,12.365242,13.247637,14.130032,15.012426,14.852346,14.6922655,14.532186,14.372105,14.212025,14.551707,14.8874855,15.223265,15.562947,15.8987255,17.284788,18.67085,20.056915,21.439074,22.825136,22.126247,21.431265,20.732376,20.033487,19.338505,19.3346,19.330696,19.330696,19.326792,19.326792,19.908546,20.490303,21.07206,21.653814,22.23557,21.403933,20.568392,19.73285,18.897306,18.061766,1.1010414,1.2415999,1.3860629,1.5266213,1.6710842,1.8116426,1.9756275,2.1435168,2.3075018,2.4714866,2.639376,2.5456703,2.455869,2.366068,2.2762666,2.1864653,2.1474214,2.1083772,2.069333,2.0263848,1.9873407,2.182561,2.377781,2.5730011,2.7682211,2.9634414,3.0141985,3.0610514,3.1118085,3.1625657,3.213323,4.9937305,6.7780423,8.55845,10.342762,12.123169,9.928895,7.7307167,5.532538,3.3343596,1.1361811,1.0580931,0.98390937,0.9058213,0.8277333,0.74964523,0.61299115,0.47633708,0.3357786,0.19912452,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.19131571,0.19912452,0.20302892,0.20693332,0.21083772,0.22255093,0.23426414,0.24207294,0.25378615,0.26159495,0.26159495,0.25769055,0.25378615,0.25378615,0.24988174,0.30844778,0.3631094,0.42167544,0.48024148,0.5388075,0.48805028,0.44119745,0.39434463,0.3474918,0.30063897,0.25378615,0.20693332,0.15617609,0.10932326,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.19912452,0.3631094,0.5231899,0.6871748,0.8511597,0.679366,0.5114767,0.339683,0.1717937,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.59346914,0.6832704,0.77697605,0.8706817,0.96438736,0.80821127,0.6559396,0.5036679,0.3513962,0.19912452,0.1756981,0.14836729,0.12494087,0.10151446,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.30844778,0.42167544,0.5309987,0.64032197,0.74964523,1.3157835,1.8858263,2.4519646,3.018103,3.5881457,3.619381,3.6467118,3.677947,3.7091823,3.736513,3.775557,3.8106966,3.8497405,3.8887846,3.9239242,4.2167544,4.5095844,4.802415,5.095245,5.388075,5.1577153,4.927356,4.6969957,4.466636,4.2362766,4.1894236,4.138666,4.087909,4.037152,3.9863946,3.8458362,3.7091823,3.5686235,3.4280653,3.2875066,3.2679846,3.2484627,3.2289407,3.2094188,3.1859922,4.240181,5.2943697,6.3446536,7.3988423,8.449126,7.9454584,7.4417906,6.9342184,6.4305506,5.9268827,6.278279,6.629675,6.9810715,7.336372,7.687768,7.4144597,7.141152,6.871748,6.5984397,6.3251314,5.899552,5.473972,5.0483923,4.6267166,4.2011366,4.3260775,4.4510183,4.575959,4.7009,4.825841,5.2084727,5.591104,5.9737353,6.356367,6.7389984,6.387602,6.036206,5.688714,5.337318,4.985922,4.263607,3.5373883,2.8111696,2.0888553,1.3626363,2.1005683,2.8424048,3.5842414,4.322173,5.0640097,7.633106,10.202203,12.771299,15.344301,17.913397,23.51231,29.111223,34.71404,40.312954,45.911865,38.8449,31.77793,24.710962,17.643993,10.573121,13.173453,15.773785,18.374117,20.97445,23.574781,24.10578,24.636778,25.163872,25.694872,26.22587,27.428427,28.630981,29.833538,31.036093,32.23865,34.089336,35.943928,37.794613,39.649204,41.499893,40.58626,39.676537,38.762905,37.849274,36.935646,38.72386,40.508175,42.292484,44.076797,45.86111,40.82443,35.78775,30.751072,25.71049,20.67381,18.214037,15.754263,13.29449,10.834716,8.374943,10.206107,12.041177,13.872341,15.7035055,17.538574,16.082233,14.625891,13.173453,11.717112,10.260769,9.956225,9.651682,9.347139,9.042596,8.738052,9.304191,9.874233,10.4403715,11.00651,11.576552,11.45942,11.346193,11.229061,11.115833,10.998701,10.791768,10.584834,10.377901,10.170968,9.964035,10.03041,10.096785,10.163159,10.2334385,10.299813,10.920613,11.541413,12.158309,12.779109,13.399908,13.16174,12.919667,12.681499,12.439425,12.201257,13.009468,13.813775,14.621986,15.430198,16.238409,16.421915,16.609327,16.792833,16.976341,17.163752,19.900738,22.637724,25.37471,28.111696,30.848682,33.687183,36.525684,39.364185,42.19878,45.03728,38.981552,32.925823,26.874,20.818274,14.762545,12.228588,9.698535,7.164578,4.630621,2.1005683,2.5769055,3.049338,3.5256753,3.998108,4.474445,3.9239242,3.3694992,2.8189783,2.2645533,1.7140326,1.9561055,2.2020829,2.4480603,2.6940374,2.9361105,2.6940374,2.4480603,2.2020829,1.9561055,1.7140326,1.7882162,1.8623998,1.9365835,2.0107672,2.0888553,2.900971,3.7130866,4.5252023,5.337318,6.1494336,6.1767645,6.2001905,6.223617,6.250948,6.2743745,5.9932575,5.708236,5.4271193,5.1460023,4.860981,4.743849,4.6228123,4.5017757,4.380739,4.263607,3.9239242,3.5842414,3.240654,2.900971,2.5612879,2.9946766,3.4280653,3.8614538,4.290938,4.7243266,4.8102236,4.8961205,4.9781127,5.0640097,5.1499066,5.388075,5.630148,5.8683167,6.1103897,6.348558,6.3056097,6.266566,6.223617,6.180669,6.13772,6.2158084,6.297801,6.375889,6.4578815,6.5359693,5.9542136,5.3724575,4.7907014,4.2089458,3.6232853,3.5530062,3.4788225,3.408543,3.3343596,3.2640803,3.416352,3.5686235,3.7208953,3.873167,4.025439,4.4978714,4.970304,5.4427366,5.9151692,6.387602,5.4505453,4.513489,3.5764325,2.639376,1.698415,3.416352,5.1303844,6.844417,8.55845,10.276386,10.065549,9.854712,9.643873,9.43694,9.226103,8.710721,8.1992445,7.687768,7.1762915,6.66091,7.309041,7.957172,8.605303,9.253433,9.901564,12.907954,15.914344,18.920732,21.931028,24.937418,24.558691,24.17606,23.79733,23.418604,23.035973,23.851994,24.668013,25.484034,26.296148,27.11217,23.621634,20.131098,16.640562,13.153932,9.663396,20.228708,30.797924,41.36714,51.932453,62.50167,51.604485,40.7112,29.814016,18.920732,8.023546,15.469242,22.911032,30.352823,37.794613,45.236404,38.59892,31.961437,25.323954,18.68647,12.0489855,9.757101,7.465217,5.173333,2.8814487,0.58566034,0.46852827,0.3513962,0.23426414,0.11713207,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.113227665,0.12494087,0.13665408,0.14836729,0.1639849,0.24597734,0.3279698,0.40996224,0.49195468,0.57394713,0.5544251,0.5349031,0.5153811,0.4958591,0.47633708,0.39434463,0.30844778,0.22645533,0.14446288,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.09761006,0.13274968,0.1678893,0.20302892,0.23816854,0.24597734,0.25378615,0.26159495,0.26940376,0.27330816,0.23035973,0.1835069,0.14055848,0.093705654,0.05075723,0.042948425,0.03513962,0.027330816,0.019522011,0.011713207,0.23426414,0.45291066,0.6715572,0.8941081,1.1127546,1.2572175,1.4016805,1.5461433,1.6906061,1.8389735,1.9170616,1.999054,2.077142,2.1591344,2.2372224,2.25284,2.2684577,2.2840753,2.2957885,2.3114061,2.5769055,2.8424048,3.1079042,3.3734035,3.638903,3.7287042,3.8224099,3.9161155,4.0059166,4.0996222,4.037152,3.9746814,3.912211,3.8497405,3.78727,4.181615,4.575959,4.9742084,5.368553,5.7628975,5.6418614,5.5169206,5.395884,5.270943,5.1499066,4.942973,4.73604,4.5291066,4.318269,4.1113358,4.365122,4.618908,4.8687897,5.1225758,5.376362,5.704332,6.036206,6.364176,6.6960497,7.0240197,7.262188,7.5003567,7.7385254,7.9766936,8.210958,8.503788,8.796618,9.089449,9.382278,9.675109,10.748819,11.818625,12.892336,13.966047,15.035853,14.832824,14.625891,14.422862,14.215929,14.012899,14.473619,14.938243,15.398962,15.863586,16.324306,17.718178,19.11205,20.502016,21.895887,23.285854,22.657246,22.028637,21.396124,20.767515,20.138906,19.580578,19.022247,18.463919,17.905588,17.351164,18.096905,18.84655,19.59229,20.338032,21.087677,20.70895,20.326319,19.947592,19.568865,19.186234,1.0619974,1.2259823,1.3860629,1.5500476,1.7140326,1.8741131,2.0498111,2.2255092,2.4012074,2.5769055,2.7486992,2.6237583,2.4988174,2.3738766,2.2489357,2.1239948,2.0732377,2.0263848,1.9756275,1.9248703,1.8741131,2.0888553,2.2996929,2.514435,2.7252727,2.9361105,3.049338,3.1625657,3.2757936,3.3890212,3.4983444,5.1616197,6.824895,8.488171,10.151445,11.810817,9.651682,7.4886436,5.3256044,3.1625657,0.999527,0.93705654,0.8745861,0.81211567,0.74964523,0.6871748,0.5505207,0.41386664,0.27330816,0.13665408,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,0.26159495,0.27330816,0.28892577,0.30063897,0.31235218,0.30063897,0.28892577,0.27330816,0.26159495,0.24988174,0.30063897,0.3513962,0.39824903,0.44900626,0.4997635,0.44900626,0.39824903,0.3513962,0.30063897,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,0.737932,0.8511597,0.96438736,1.0737107,1.1869383,0.94876975,0.7106012,0.47633708,0.23816854,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.3513962,0.44900626,0.5505207,0.6481308,0.74964523,1.475864,2.1981785,2.9243972,3.6506162,4.376835,4.251894,4.126953,3.998108,3.873167,3.7482262,3.7638438,3.775557,3.78727,3.7989833,3.8106966,4.123049,4.4393053,4.7516575,5.0640097,5.376362,5.212377,5.0483923,4.8883114,4.7243266,4.564246,4.5369153,4.513489,4.4861584,4.462732,4.4393053,4.2753205,4.1113358,3.951255,3.78727,3.6232853,3.638903,3.6506162,3.6623292,3.6740425,3.6857557,4.6384296,5.5871997,6.5359693,7.4886436,8.437413,7.7892823,7.137247,6.4891167,5.8370814,5.1889505,5.786324,6.387602,6.98888,7.5862536,8.187531,7.7892823,7.387129,6.98888,6.5867267,6.1884775,5.610626,5.036679,4.462732,3.8887846,3.310933,3.638903,3.9629683,4.2870336,4.6110992,4.939069,5.2865605,5.6379566,5.989353,6.336845,6.688241,6.1494336,5.610626,5.0757227,4.5369153,3.998108,3.5256753,3.049338,2.5769055,2.1005683,1.6242313,2.3114061,2.998581,3.6857557,4.376835,5.0640097,7.6370106,10.213917,12.786918,15.363823,17.936825,24.39861,30.860395,37.326084,43.787872,50.249657,42.214397,34.175232,26.136068,18.10081,10.061645,12.888432,15.711315,18.538101,21.360985,24.187773,24.476698,24.761719,25.050644,25.335667,25.624592,26.948185,28.27568,29.599274,30.926771,32.250362,34.089336,35.924404,37.76338,39.598446,41.43742,39.86395,38.286568,36.713093,35.135715,33.56224,35.674522,37.786804,39.899086,42.011368,44.12365,39.836617,35.549583,31.262548,26.975515,22.688482,19.889025,17.085665,14.286208,11.486752,8.687295,10.936231,13.189071,15.438006,17.686943,19.935879,17.788456,15.637131,13.4858055,11.338385,9.187058,8.874706,8.562354,8.250002,7.9376497,7.6252975,7.437886,7.250475,7.0630636,6.8756523,6.688241,7.375416,8.062591,8.749765,9.43694,10.124115,9.839094,9.550168,9.261242,8.976221,8.687295,8.624825,8.562354,8.499884,8.437413,8.374943,8.925464,9.475985,10.0265045,10.573121,11.123642,10.686349,10.249056,9.811763,9.37447,8.937177,9.37447,9.811763,10.249056,10.686349,11.123642,11.326671,11.525795,11.72492,11.924045,12.123169,15.738646,19.350218,22.96179,26.573362,30.188839,32.500244,34.81165,37.12696,39.438366,41.749775,35.77604,29.798397,23.824663,17.850927,11.873287,9.788337,7.699481,5.610626,3.5256753,1.43682,1.901444,2.3621633,2.8267872,3.2875066,3.7482262,3.2250361,2.7018464,2.174752,1.6515622,1.1244678,1.43682,1.7491722,2.0615244,2.3738766,2.6862288,2.514435,2.338737,2.1630387,1.9873407,1.8116426,1.6359446,1.4641509,1.2884527,1.1127546,0.93705654,2.0107672,3.0883822,4.1620927,5.2358036,6.3134184,6.461786,6.6140575,6.7624245,6.910792,7.0630636,6.699954,6.336845,5.9737353,5.610626,5.251421,5.173333,5.099149,5.024966,4.950782,4.8765984,4.4393053,3.998108,3.5608149,3.1235218,2.6862288,3.2757936,3.8614538,4.4510183,5.036679,5.6262436,5.6379566,5.64967,5.661383,5.6730967,5.688714,6.001066,6.3134184,6.6257706,6.9381227,7.250475,7.0513506,6.8483214,6.649197,6.4500723,6.250948,6.3251314,6.3993154,6.473499,6.551587,6.6257706,6.1611466,5.700427,5.2358036,4.775084,4.3143644,4.1620927,4.0137253,3.8614538,3.7130866,3.5608149,3.7638438,3.9629683,4.1620927,4.3612175,4.564246,5.173333,5.786324,6.3993154,7.012306,7.6252975,6.387602,5.1499066,3.912211,2.6745155,1.43682,3.474918,5.5130157,7.551114,9.589212,11.623405,11.0260315,10.424754,9.823476,9.226103,8.624825,8.226576,7.824422,7.426173,7.0240197,6.6257706,7.4886436,8.351517,9.21439,10.073358,10.936231,14.512663,18.089096,21.661623,25.238056,28.810585,28.099983,27.389381,26.674877,25.964275,25.24977,26.026745,26.799816,27.576794,28.349865,29.12684,25.085785,21.048632,17.01148,12.974329,8.937177,18.514675,28.08827,37.661865,47.239365,56.812958,47.01291,37.212856,27.412807,17.612759,7.812709,17.24965,26.68659,36.12353,45.564373,55.001316,46.450672,37.900032,29.349392,20.79875,12.24811,9.80005,7.3519893,4.900025,2.4480603,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.28892577,0.38653582,0.48805028,0.58566034,0.6871748,0.6637484,0.63641757,0.61299115,0.58566034,0.5622339,0.46071947,0.3631094,0.26159495,0.1639849,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.10151446,0.13665408,0.1756981,0.21083772,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.31235218,0.43729305,0.5622339,0.6871748,0.81211567,0.8745861,0.93705654,0.999527,1.0619974,1.1244678,1.4485333,1.7765031,2.1005683,2.4246337,2.7486992,2.639376,2.5261483,2.4129205,2.2996929,2.1864653,2.2255092,2.260649,2.2996929,2.338737,2.3738766,2.7994564,3.2250361,3.6506162,4.0761957,4.5017757,4.423688,4.349504,4.2753205,4.2011366,4.123049,3.78727,3.4514916,3.1118085,2.77603,2.436347,2.6862288,2.9361105,3.1859922,3.435874,3.6857557,3.998108,4.3143644,4.6267166,4.939069,5.251421,5.5989127,5.950309,6.3017054,6.649197,7.000593,7.348085,7.699481,8.050878,8.398369,8.749765,10.010887,11.275913,12.537036,13.798158,15.063184,14.813302,14.56342,14.313539,14.063657,13.813775,14.399435,14.989,15.57466,16.164225,16.749886,18.151566,19.549341,20.951023,22.348799,23.750479,23.188246,22.62601,22.063778,21.501543,20.93931,19.826555,18.7138,17.601046,16.48829,15.375536,16.289165,17.198893,18.112522,19.026152,19.935879,20.013966,20.08815,20.162333,20.236517,20.310701,1.0893283,1.2455044,1.4016805,1.5617609,1.717937,1.8741131,2.0380979,2.2059872,2.3699722,2.533957,2.7018464,2.5808098,2.463678,2.3465457,2.2294137,2.1122816,2.0810463,2.0459068,2.0146716,1.9834363,1.9482968,2.174752,2.4012074,2.6237583,2.8502135,3.076669,3.2094188,3.3460727,3.4788225,3.6154766,3.7482262,5.239708,6.7311897,8.218767,9.710248,11.20173,9.148014,7.094299,5.040583,2.9907722,0.93705654,0.8667773,0.79649806,0.7262188,0.6559396,0.58566034,0.47633708,0.3670138,0.25769055,0.14836729,0.039044023,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.1835069,0.20302892,0.22255093,0.24207294,0.26159495,0.26940376,0.27330816,0.27721256,0.28111696,0.28892577,0.27721256,0.26940376,0.25769055,0.24597734,0.23816854,0.28111696,0.3279698,0.3709182,0.41777104,0.46071947,0.42557985,0.38653582,0.3513962,0.31235218,0.27330816,0.24597734,0.21474212,0.1835069,0.15617609,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.11713207,0.21083772,0.30063897,0.39434463,0.48805028,0.59737355,0.7066968,0.8160201,0.92924774,1.038571,1.0502841,1.0619974,1.0737107,1.0893283,1.1010414,0.8941081,0.6910792,0.48414588,0.28111696,0.07418364,0.078088045,0.08589685,0.08980125,0.093705654,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.042948425,0.08589685,0.12884527,0.1717937,0.21083772,0.5114767,0.81211567,1.1127546,1.4133936,1.7140326,2.135708,2.5573835,2.979059,3.4007344,3.8263142,3.8614538,3.900498,3.9356375,3.9746814,4.0137253,4.1581883,4.3026514,4.447114,4.591577,4.73604,4.853172,4.9742084,5.0913405,5.2084727,5.3256044,5.196759,5.0718184,4.942973,4.814128,4.689187,4.747753,4.806319,4.8687897,4.927356,4.985922,4.8492675,4.7126136,4.575959,4.4393053,4.298747,4.2597027,4.220659,4.181615,4.138666,4.0996222,4.9156423,5.7316628,6.5437784,7.3597984,8.175818,7.8634663,7.5550184,7.2465706,6.9342184,6.6257706,7.1216297,7.6135845,8.109444,8.605303,9.101162,8.6131115,8.125061,7.6370106,7.1489606,6.66091,5.919074,5.173333,4.4275923,3.6818514,2.9361105,3.4788225,4.01763,4.5564375,5.099149,5.6379566,5.9620223,6.2860875,6.6140575,6.9381227,7.262188,7.012306,6.7624245,6.5125427,6.262661,6.012779,5.376362,4.73604,4.0996222,3.4632049,2.8267872,3.8497405,4.8765984,5.899552,6.9264097,7.9493628,10.877665,13.805966,16.734268,19.658665,22.586967,28.342056,34.097145,39.852234,45.607323,51.36241,43.420856,35.483208,27.541653,19.604004,11.66245,13.809871,15.957292,18.104713,20.252134,22.399555,23.153105,23.906654,24.6563,25.40985,26.163399,28.099983,30.036566,31.97315,33.91364,35.85022,36.849747,37.849274,38.8488,39.848328,40.85176,39.168964,37.49007,35.811176,34.12838,32.449486,33.839455,35.22942,36.61939,38.009357,39.399323,35.721375,32.04343,28.365482,24.69144,21.013493,19.326792,17.636185,15.949483,14.262781,12.576079,14.130032,15.683984,17.24184,18.795792,20.349745,18.206228,16.066616,13.923099,11.779582,9.636065,9.276859,8.913751,8.550641,8.187531,7.824422,7.387129,6.949836,6.5125427,6.0752497,5.6379566,6.3134184,6.98888,7.6643414,8.335898,9.01136,8.886419,8.761478,8.636538,8.511597,8.386656,8.550641,8.718531,8.882515,9.0465,9.21439,9.382278,9.554072,9.721962,9.893755,10.061645,9.698535,9.331521,8.968412,8.601398,8.238289,8.722435,9.20658,9.690726,10.178777,10.662923,12.373051,14.0831785,15.793307,17.503435,19.213564,22.286327,25.359093,28.431858,31.500717,34.573483,36.275803,37.974216,39.676537,41.37495,43.073364,36.455402,29.833538,23.215576,16.59371,9.975748,8.238289,6.504734,4.7711797,3.0337205,1.3001659,1.6437533,1.9912452,2.3348327,2.67842,3.0259118,2.6237583,2.2216048,1.815547,1.4133936,1.0112402,1.2767396,1.542239,1.8077383,2.0732377,2.338737,2.5300527,2.7213683,2.9165885,3.1079042,3.2992198,3.6857557,4.0761957,4.462732,4.8492675,5.2358036,6.0518236,6.8678436,7.6838636,8.495979,9.311999,8.987934,8.663869,8.335898,8.011833,7.687768,7.1880045,6.688241,6.1884775,5.688714,5.1889505,5.114767,5.040583,4.970304,4.8961205,4.825841,4.575959,4.3260775,4.0761957,3.8263142,3.5764325,3.8263142,4.0761957,4.3260775,4.575959,4.825841,5.12648,5.4310236,5.7316628,6.036206,6.336845,6.4578815,6.578918,6.6960497,6.817086,6.9381227,6.8483214,6.75852,6.6687193,6.578918,6.4891167,6.547683,6.606249,6.6687193,6.727285,6.785851,6.289992,5.794133,5.2943697,4.7985106,4.298747,4.271416,4.240181,4.2089458,4.181615,4.1503797,4.3612175,4.5681505,4.7789884,4.989826,5.2006636,5.7316628,6.2587566,6.7897553,7.320754,7.8517528,6.969358,6.0908675,5.2084727,4.3299823,3.4514916,5.0718184,6.688241,8.308568,9.928895,11.549222,10.889378,10.229534,9.56969,8.909846,8.250002,7.800996,7.355894,6.9068875,6.461786,6.012779,7.47693,8.937177,10.401327,11.861574,13.325725,16.519526,19.709423,22.903223,26.09312,29.28692,28.646599,28.006277,27.365955,26.725634,26.089216,26.987228,27.889145,28.787157,29.689075,30.587088,26.682686,22.778282,18.87388,14.965574,11.061172,19.014439,26.967707,34.920975,42.87424,50.823605,42.19097,33.55834,24.925705,16.29307,7.6643414,15.76988,23.871515,31.977055,40.082592,48.188133,40.523792,32.85945,25.191204,17.526861,9.86252,7.890797,5.9229784,3.951255,1.9834363,0.011713207,0.08589685,0.15617609,0.23035973,0.30063897,0.37482262,0.78868926,1.1986516,1.6125181,2.0263848,2.436347,1.9912452,1.542239,1.0932326,0.6481308,0.19912452,0.19912452,0.19912452,0.19912452,0.19912452,0.19912452,0.30063897,0.39824903,0.4997635,0.60127795,0.698888,0.6559396,0.60908675,0.5661383,0.5192855,0.47633708,0.39434463,0.31625658,0.23426414,0.15617609,0.07418364,0.078088045,0.078088045,0.08199245,0.08589685,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.21083772,0.19912452,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12103647,0.10541886,0.08980125,0.07418364,0.07418364,0.07027924,0.06637484,0.06637484,0.062470436,0.05466163,0.046852827,0.039044023,0.031235218,0.023426414,0.05075723,0.078088045,0.10932326,0.13665408,0.1639849,0.26159495,0.3631094,0.46071947,0.5622339,0.6637484,0.7106012,0.75745404,0.80430686,0.8511597,0.9019169,1.1674163,1.43682,1.7023194,1.9717231,2.2372224,2.1513257,2.069333,1.9834363,1.8975395,1.8116426,1.8428779,1.8741131,1.901444,1.9326792,1.9639144,2.3035975,2.6432803,2.9829633,3.3226464,3.6623292,3.6154766,3.5686235,3.521771,3.4710135,3.4241607,3.174279,2.9243972,2.6745155,2.4246337,2.174752,2.416825,2.6588979,2.900971,3.1430438,3.3890212,3.6740425,3.959064,4.2440853,4.5291066,4.814128,5.3217,5.8292727,6.336845,6.844417,7.348085,7.4886436,7.629202,7.7697606,7.910319,8.050878,9.093353,10.139732,11.186112,12.228588,13.274967,13.1266,12.974329,12.825961,12.67369,12.525322,13.173453,13.821584,14.465811,15.113941,15.762072,17.226223,18.694279,20.158428,21.62258,23.086731,22.629915,22.1731,21.716286,21.25947,20.79875,19.889025,18.9793,18.069574,17.159847,16.250122,16.91387,17.573715,18.237463,18.90121,19.561056,19.73285,19.900738,20.072533,20.244326,20.412214,1.1127546,1.2650263,1.4172981,1.5695697,1.7218413,1.8741131,2.0302892,2.1864653,2.338737,2.494913,2.6510892,2.541766,2.4285383,2.3192148,2.2098918,2.1005683,2.084951,2.069333,2.0537157,2.0380979,2.0263848,2.260649,2.4988174,2.736986,2.9751544,3.213323,3.3694992,3.5256753,3.6857557,3.8419318,3.998108,5.3177958,6.6335793,7.9532676,9.269051,10.588739,8.644346,6.703859,4.759466,2.8189783,0.8745861,0.79649806,0.71841,0.6442264,0.5661383,0.48805028,0.40605783,0.3240654,0.23816854,0.15617609,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.13665408,0.1639849,0.19131571,0.21864653,0.24597734,0.27330816,0.27330816,0.26940376,0.26940376,0.26549935,0.26159495,0.25378615,0.24597734,0.23816854,0.23426414,0.22645533,0.26549935,0.30454338,0.3435874,0.38653582,0.42557985,0.39824903,0.37482262,0.3513962,0.3240654,0.30063897,0.27721256,0.25378615,0.23426414,0.21083772,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.23426414,0.42167544,0.60518235,0.78868926,0.97610056,1.0698062,1.1635119,1.261122,1.3548276,1.4485333,1.3626363,1.2767396,1.1869383,1.1010414,1.0112402,0.8394465,0.6676528,0.4958591,0.3240654,0.14836729,0.16008049,0.1717937,0.1796025,0.19131571,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.6754616,1.175225,1.6749885,2.174752,2.6745155,2.795552,2.9165885,3.0337205,3.154757,3.2757936,3.474918,3.6740425,3.873167,4.0761957,4.2753205,4.552533,4.829746,5.1069584,5.3841705,5.661383,5.5832953,5.5091114,5.4310236,5.3529353,5.2748475,5.181142,5.0913405,4.997635,4.903929,4.814128,4.958591,5.1030536,5.2475166,5.3919797,5.5364423,5.423215,5.3138914,5.2006636,5.087436,4.9742084,4.884407,4.7907014,4.6969957,4.60329,4.513489,5.192855,5.872221,6.551587,7.230953,7.914223,7.941554,7.9727893,8.0040245,8.031356,8.062591,8.453031,8.843472,9.2339115,9.6243515,10.010887,9.43694,8.862993,8.289046,7.7111945,7.137247,6.223617,5.3060827,4.3924527,3.4788225,2.5612879,3.3187418,4.0722914,4.825841,5.5832953,6.336845,6.6374836,6.9381227,7.238762,7.5394006,7.8361354,7.8751793,7.914223,7.9493628,7.988407,8.023546,7.223144,6.426646,5.6262436,4.825841,4.025439,5.388075,6.7507114,8.113348,9.475985,10.838621,14.118319,17.398016,20.677715,23.957413,27.23711,32.285503,37.333893,42.378384,47.426773,52.475166,44.63122,36.791183,28.947239,21.103294,13.263254,14.73131,16.20327,17.671324,19.143284,20.61134,21.829514,23.047686,24.26586,25.484034,26.698303,29.251781,31.801357,34.35093,36.900505,39.45008,39.614067,39.774147,39.93813,40.09821,40.262196,38.477882,36.693573,34.90926,33.121044,31.336733,32.004387,32.67204,33.33969,34.007343,34.674995,31.606136,28.54118,25.47232,22.40346,19.338505,18.760653,18.186707,17.612759,17.03881,16.46096,17.323833,18.182802,19.041769,19.900738,20.76361,18.627903,16.492195,14.356487,12.220779,10.088976,9.675109,9.261242,8.85128,8.437413,8.023546,7.336372,6.649197,5.9620223,5.2748475,4.5876727,5.251421,5.911265,6.575013,7.238762,7.898606,7.9376497,7.9766936,8.011833,8.050878,8.086017,8.480362,8.870802,9.265146,9.655587,10.049932,9.839094,9.628256,9.421323,9.2104845,8.999647,8.706817,8.413987,8.121157,7.8283267,7.5394006,8.070399,8.601398,9.136301,9.6673,10.198298,13.419431,16.640562,19.861694,23.078922,26.300053,28.834011,31.364063,33.89802,36.431976,38.96203,40.051357,41.136784,42.22611,43.311535,44.400864,37.13477,29.868677,22.60649,15.340397,8.074304,6.6921453,5.309987,3.9278288,2.5456703,1.1635119,1.3899672,1.6164225,1.8467822,2.0732377,2.2996929,2.018576,1.7413634,1.4602464,1.1791295,0.9019169,1.116659,1.3353056,1.5539521,1.7686942,1.9873407,2.5456703,3.1079042,3.6662338,4.2284675,4.786797,5.7394714,6.688241,7.6370106,8.58578,9.538455,10.09288,10.647305,11.20173,11.756155,12.31058,11.514082,10.71368,9.913278,9.112875,8.312472,7.676055,7.0357327,6.3993154,5.7628975,5.12648,5.056201,4.985922,4.9156423,4.845363,4.775084,4.7126136,4.650143,4.5876727,4.5252023,4.462732,4.376835,4.2870336,4.2011366,4.1113358,4.025439,4.618908,5.2084727,5.801942,6.395411,6.98888,6.914696,6.844417,6.7702336,6.6960497,6.6257706,6.6452928,6.6648145,6.6843367,6.703859,6.7233806,6.7702336,6.813182,6.860035,6.9068875,6.949836,6.4188375,5.883934,5.3529353,4.8219366,4.2870336,4.376835,4.466636,4.5564375,4.646239,4.73604,4.958591,5.1772375,5.395884,5.618435,5.8370814,6.2860875,6.7311897,7.180196,7.629202,8.074304,7.551114,7.0318284,6.5086384,5.985449,5.462259,6.6648145,7.8673706,9.069926,10.272482,11.475039,10.756628,10.034314,9.315904,8.59359,7.8751793,7.37932,6.883461,6.3915067,5.8956475,5.3997884,7.461313,9.526741,11.588266,13.64979,15.711315,18.522484,21.333654,24.140919,26.95209,29.763258,29.193216,28.627077,28.06094,27.490896,26.924759,27.951616,28.97457,30.001427,31.02438,32.05124,28.27568,24.504028,20.732376,16.960724,13.189071,19.518106,25.847143,32.176178,38.50912,44.838154,37.37294,29.90772,22.442505,14.977287,7.5120697,14.286208,21.056442,27.83058,34.60081,41.37495,34.593002,27.814962,21.033014,14.254972,7.47693,5.985449,4.493967,3.0063896,1.5149081,0.023426414,0.1717937,0.31625658,0.46071947,0.60518235,0.74964523,1.5500476,2.35045,3.1508527,3.951255,4.7516575,3.853645,2.959537,2.0654287,1.1713207,0.27330816,0.26159495,0.24988174,0.23816854,0.22645533,0.21083772,0.31235218,0.41386664,0.5114767,0.61299115,0.7106012,0.6481308,0.58175594,0.5192855,0.45291066,0.38653582,0.3279698,0.26940376,0.20693332,0.14836729,0.08589685,0.093705654,0.09761006,0.10151446,0.10932326,0.113227665,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.21864653,0.20302892,0.1835069,0.1678893,0.14836729,0.14446288,0.14055848,0.13665408,0.12884527,0.12494087,0.10932326,0.093705654,0.078088045,0.06637484,0.05075723,0.06637484,0.08589685,0.10151446,0.12103647,0.13665408,0.21083772,0.28892577,0.3631094,0.43729305,0.5114767,0.5466163,0.57785153,0.60908675,0.6442264,0.6754616,0.8862993,1.0932326,1.3040704,1.5149081,1.7257458,1.6671798,1.6086137,1.5539521,1.4953861,1.43682,1.4602464,1.4836729,1.5031948,1.5266213,1.5500476,1.8038338,2.0615244,2.3153105,2.5690966,2.8267872,2.803361,2.7838387,2.7643168,2.7447948,2.7252727,2.5612879,2.4012074,2.2372224,2.0732377,1.9131571,2.1474214,2.3816853,2.6159496,2.854118,3.0883822,3.3460727,3.6037633,3.8614538,4.1191444,4.376835,5.040583,5.704332,6.36808,7.0357327,7.699481,7.629202,7.558923,7.4886436,7.4183645,7.348085,8.175818,9.0035515,9.8312845,10.6590185,11.486752,11.435994,11.389141,11.338385,11.287627,11.23687,11.943566,12.654168,13.360865,14.067561,14.774258,16.304783,17.83531,19.365835,20.89636,22.426888,22.071587,21.72019,21.368793,21.013493,20.662096,19.9554,19.248703,18.538101,17.831406,17.124708,17.538574,17.948538,18.362404,18.77627,19.186234,19.451733,19.717232,19.98273,20.24823,20.51373,1.1361811,1.2845483,1.4329157,1.5812829,1.7257458,1.8741131,2.018576,2.1669433,2.3114061,2.455869,2.6003318,2.4988174,2.3933985,2.2918842,2.1903696,2.0888553,2.0888553,2.0927596,2.096664,2.096664,2.1005683,2.35045,2.6003318,2.8502135,3.1000953,3.349977,3.5295796,3.7091823,3.8887846,4.068387,4.251894,5.395884,6.5398736,7.6838636,8.831758,9.975748,8.140678,6.309514,4.478349,2.6432803,0.81211567,0.7262188,0.6442264,0.5583295,0.47243267,0.38653582,0.3318742,0.27721256,0.22255093,0.1678893,0.113227665,0.113227665,0.113227665,0.113227665,0.113227665,0.113227665,0.14836729,0.1835069,0.21864653,0.25378615,0.28892577,0.27721256,0.26940376,0.25769055,0.24597734,0.23816854,0.23426414,0.22645533,0.22255093,0.21864653,0.21083772,0.24597734,0.28111696,0.31625658,0.3513962,0.38653582,0.37482262,0.3631094,0.3513962,0.3357786,0.3240654,0.30844778,0.29673457,0.28111696,0.26549935,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.3513962,0.62860876,0.9058213,1.1869383,1.4641509,1.542239,1.6242313,1.7023194,1.7843118,1.8623998,1.6749885,1.4875772,1.3001659,1.1127546,0.92534333,0.78478485,0.6442264,0.5036679,0.3631094,0.22645533,0.23816854,0.25378615,0.26940376,0.28502136,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.8355421,1.5383345,2.2372224,2.9361105,3.638903,3.455396,3.2718892,3.0883822,2.9087796,2.7252727,3.0883822,3.4514916,3.8106966,4.173806,4.5369153,4.9468775,5.35684,5.7668023,6.1767645,6.5867267,6.3134184,6.044015,5.7707067,5.4973984,5.22409,5.169429,5.1108627,5.0522966,4.9937305,4.939069,5.169429,5.395884,5.6262436,5.8566036,6.086963,6.001066,5.911265,5.825368,5.735567,5.64967,5.505207,5.3607445,5.2162814,5.0718184,4.9234514,5.4700675,6.016684,6.559396,7.1060123,7.648724,8.019642,8.39056,8.761478,9.128492,9.499411,9.784432,10.069453,10.354475,10.639496,10.924518,10.260769,9.600925,8.937177,8.273428,7.6135845,6.5281606,5.4427366,4.357313,3.2718892,2.1864653,3.1586614,4.126953,5.099149,6.067441,7.0357327,7.3129454,7.5862536,7.8634663,8.136774,8.413987,8.738052,9.062118,9.386183,9.714153,10.0382185,9.073831,8.113348,7.1489606,6.1884775,5.22409,6.9264097,8.624825,10.323239,12.025558,13.723974,17.358973,20.990067,24.62116,28.256159,31.887253,36.228947,40.56674,44.908436,49.246227,53.58792,45.841587,38.099155,30.352823,22.60649,14.864059,15.656653,16.449247,17.24184,18.034433,18.823124,20.50592,22.188719,23.871515,25.554314,27.23711,30.399675,33.56224,36.724808,39.887375,43.04994,42.374477,41.699017,41.023556,40.34809,39.676537,37.786804,35.89317,34.00344,32.11371,30.223978,30.169315,30.114655,30.059994,30.005331,29.95067,27.490896,25.035027,22.579159,20.119385,17.663515,18.19842,18.737226,19.276033,19.810938,20.349745,20.51373,20.68162,20.845604,21.009588,21.173573,19.045673,16.921679,14.79378,12.665881,10.537982,10.073358,9.612638,9.151918,8.687295,8.226576,7.2856145,6.348558,5.4115014,4.474445,3.5373883,4.1894236,4.8375545,5.4856853,6.13772,6.785851,6.98888,7.1880045,7.387129,7.5862536,7.7892823,8.406178,9.026978,9.647778,10.268578,10.889378,10.295909,9.706344,9.116779,8.527214,7.9376497,7.719003,7.4964523,7.277806,7.0591593,6.8366084,7.4183645,7.996216,8.577971,9.155824,9.737579,14.469715,19.197947,23.926178,28.658312,33.386543,35.381695,37.37294,39.364185,41.359333,43.35058,43.826916,44.299347,44.775684,45.24812,45.724453,37.814137,29.903816,21.993498,14.0831785,6.1767645,5.1460023,4.11524,3.084478,2.0537157,1.0268579,1.1361811,1.2455044,1.3548276,1.4641509,1.5734742,1.4172981,1.261122,1.1010414,0.94486535,0.78868926,0.95657855,1.1283722,1.2962615,1.4680552,1.6359446,2.5651922,3.4905357,4.4197836,5.349031,6.2743745,7.7892823,9.300286,10.81129,12.326198,13.837202,14.133936,14.426766,14.723501,15.016331,15.313066,14.036326,12.763491,11.486752,10.213917,8.937177,8.164105,7.387129,6.6140575,5.8370814,5.0640097,4.9937305,4.927356,4.860981,4.7907014,4.7243266,4.8492675,4.9742084,5.099149,5.22409,5.349031,4.9234514,4.5017757,4.0761957,3.6506162,3.2250361,4.1074314,4.989826,5.872221,6.754616,7.6370106,7.3715115,7.1060123,6.844417,6.578918,6.3134184,6.4422636,6.571109,6.703859,6.832704,6.9615493,6.9927845,7.0240197,7.0513506,7.082586,7.113821,6.5437784,5.9776397,5.4115014,4.841459,4.2753205,4.4861584,4.6930914,4.903929,5.114767,5.3256044,5.5559645,5.786324,6.016684,6.2431393,6.473499,6.8405128,7.2036223,7.570636,7.9337454,8.300759,8.136774,7.968885,7.8049,7.6409154,7.47693,8.261715,9.0465,9.8312845,10.61607,11.400854,10.619974,9.839094,9.058213,8.281238,7.5003567,6.957645,6.4149327,5.872221,5.3295093,4.786797,7.4495993,10.112402,12.775204,15.438006,18.10081,20.529346,22.953981,25.382519,27.811058,30.235691,29.743736,29.247877,28.752018,28.256159,27.764204,28.912098,30.063898,31.211792,32.36359,33.511486,29.872581,26.233679,22.590872,18.95197,15.313066,20.021774,24.72658,29.43529,34.143997,38.8488,32.551003,26.2532,19.9554,13.661504,7.363703,12.802535,18.241367,23.684105,29.122936,34.561768,28.66612,22.774378,16.87873,10.983084,5.087436,4.0761957,3.06886,2.05762,1.0463798,0.039044023,0.25378615,0.47243267,0.6910792,0.9058213,1.1244678,2.3114061,3.4983444,4.689187,5.8761253,7.0630636,5.7199492,4.376835,3.0337205,1.6906061,0.3513962,0.3240654,0.30063897,0.27330816,0.24988174,0.22645533,0.3240654,0.42557985,0.5231899,0.62470436,0.7262188,0.64032197,0.5544251,0.46852827,0.38653582,0.30063897,0.26159495,0.21864653,0.1796025,0.14055848,0.10151446,0.10932326,0.113227665,0.12103647,0.12884527,0.13665408,0.13665408,0.13665408,0.13665408,0.13665408,0.13665408,0.1756981,0.21083772,0.24988174,0.28892577,0.3240654,0.30454338,0.28502136,0.26549935,0.24597734,0.22645533,0.21864653,0.21083772,0.20302892,0.19522011,0.18741131,0.1639849,0.14055848,0.12103647,0.09761006,0.07418364,0.08199245,0.08980125,0.09761006,0.10541886,0.113227665,0.1639849,0.21083772,0.26159495,0.31235218,0.3631094,0.37872702,0.39824903,0.41386664,0.43338865,0.44900626,0.60127795,0.75354964,0.9058213,1.0580931,1.2142692,1.183034,1.1517987,1.1205635,1.0932326,1.0619974,1.077615,1.0932326,1.1088502,1.1205635,1.1361811,1.3079748,1.475864,1.6476578,1.815547,1.9873407,1.9951496,2.0029583,2.0107672,2.018576,2.0263848,1.9482968,1.8741131,1.7999294,1.7257458,1.6515622,1.8780174,2.1044729,2.330928,2.5612879,2.787743,3.018103,3.2484627,3.4788225,3.7091823,3.9356375,4.759466,5.5832953,6.4032197,7.2270484,8.050878,7.7697606,7.4886436,7.211431,6.930314,6.649197,7.2582836,7.871275,8.480362,9.089449,9.698535,9.749292,9.80005,9.850807,9.901564,9.948417,10.717585,11.486752,12.252014,13.021181,13.786445,15.383345,16.976341,18.573242,20.166237,21.763138,21.513256,21.267279,21.021301,20.77142,20.525442,20.021774,19.514202,19.010534,18.506866,17.999294,18.163279,18.32336,18.487345,18.651329,18.81141,19.170614,19.533724,19.89293,20.252134,20.61134,1.1635119,1.3040704,1.4485333,1.5890918,1.7335546,1.8741131,2.0107672,2.1435168,2.280171,2.416825,2.5495746,2.455869,2.358259,2.2645533,2.1708477,2.0732377,2.096664,2.1161861,2.135708,2.15523,2.174752,2.436347,2.7018464,2.9634414,3.2250361,3.4866312,3.68966,3.892689,4.095718,4.298747,4.5017757,5.473972,6.446168,7.4183645,8.39056,9.362757,7.6409154,5.919074,4.193328,2.4714866,0.74964523,0.6559396,0.5661383,0.47243267,0.37872702,0.28892577,0.26159495,0.23426414,0.20693332,0.1756981,0.14836729,0.13665408,0.12494087,0.113227665,0.10151446,0.08589685,0.12884527,0.1717937,0.21474212,0.25769055,0.30063897,0.28111696,0.26549935,0.24597734,0.23035973,0.21083772,0.21083772,0.20693332,0.20693332,0.20302892,0.19912452,0.23035973,0.26159495,0.28892577,0.32016098,0.3513962,0.3513962,0.3513962,0.3513962,0.3513962,0.3513962,0.3435874,0.3357786,0.3279698,0.32016098,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.46852827,0.8394465,1.2103647,1.5812829,1.9482968,2.0146716,2.0810463,2.1435168,2.2098918,2.2762666,1.9873407,1.698415,1.4133936,1.1244678,0.8394465,0.7301232,0.62079996,0.5153811,0.40605783,0.30063897,0.32016098,0.339683,0.359205,0.37872702,0.39824903,0.32016098,0.23816854,0.16008049,0.078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.999527,1.901444,2.7994564,3.7013733,4.5993857,4.11524,3.631094,3.1430438,2.6588979,2.174752,2.7018464,3.2250361,3.7482262,4.2753205,4.7985106,5.3412223,5.883934,6.426646,6.969358,7.5120697,7.043542,6.578918,6.1103897,5.6418614,5.173333,5.153811,5.1303844,5.1069584,5.083532,5.0640097,5.376362,5.6926184,6.008875,6.321227,6.6374836,6.575013,6.5125427,6.4500723,6.387602,6.3251314,6.126007,5.930787,5.7316628,5.5364423,5.337318,5.74728,6.1572423,6.5672045,6.9771667,7.387129,8.097731,8.8083315,9.518932,10.22563,10.936231,11.115833,11.29934,11.478943,11.6585455,11.838148,11.088503,10.338858,9.589212,8.835662,8.086017,6.832704,5.579391,4.322173,3.06886,1.8116426,2.998581,4.181615,5.368553,6.551587,7.7385254,7.988407,8.238289,8.488171,8.738052,8.987934,9.600925,10.213917,10.826907,11.435994,12.0489855,10.924518,9.80005,8.675582,7.551114,6.426646,8.460839,10.498938,12.537036,14.575133,16.613232,20.595722,24.582117,28.568512,32.551003,36.537395,40.16849,43.80349,47.43458,51.065678,54.700676,47.051952,39.40713,31.758408,24.109684,16.46096,16.578093,16.69132,16.808453,16.921679,17.03881,19.186234,21.333654,23.481075,25.628496,27.775917,31.551476,35.323128,39.098682,42.87424,46.6498,45.138794,43.623886,42.112885,40.60188,39.08697,37.09182,35.096672,33.10152,31.106373,29.111223,28.334248,27.557272,26.780294,26.003319,25.226343,23.375656,21.528873,19.682093,17.83531,15.988527,17.636185,19.287746,20.93931,22.586967,24.23853,23.707531,23.176533,22.645533,22.118439,21.58744,19.46735,17.34726,15.227169,13.107079,10.986988,10.475512,9.964035,9.448653,8.937177,8.4257,7.238762,6.0518236,4.860981,3.6740425,2.4871042,3.1235218,3.7638438,4.4002614,5.036679,5.6730967,6.036206,6.3993154,6.7624245,7.125534,7.4886436,8.335898,9.183154,10.03041,10.877665,11.72492,10.756628,9.784432,8.81614,7.843944,6.8756523,6.727285,6.578918,6.4305506,6.2860875,6.13772,6.7663293,7.3910336,8.019642,8.648251,9.276859,15.516094,21.75533,27.994564,34.2338,40.473034,41.929375,43.381813,44.83425,46.28669,47.73913,47.598568,47.461914,47.32526,47.188606,47.048046,38.493504,29.938957,21.38441,12.829865,4.2753205,3.5959544,2.920493,2.241127,1.5656652,0.8862993,0.8784905,0.8706817,0.8667773,0.8589685,0.8511597,0.8160201,0.78088045,0.74574083,0.7106012,0.6754616,0.79649806,0.92143893,1.0424755,1.1635119,1.2884527,2.5808098,3.8770714,5.173333,6.46569,7.7619514,9.839094,11.912332,13.989473,16.062712,18.135948,18.171087,18.206228,18.241367,18.276506,18.311647,16.562475,14.813302,13.06413,11.311053,9.561881,8.648251,7.7385254,6.824895,5.911265,5.001539,4.9351645,4.8687897,4.806319,4.7399445,4.6735697,4.985922,5.298274,5.610626,5.9268827,6.239235,5.473972,4.7126136,3.951255,3.1859922,2.4246337,3.5959544,4.7711797,5.9425,7.113821,8.289046,7.8283267,7.3715115,6.914696,6.4578815,6.001066,6.239235,6.481308,6.719476,6.9615493,7.1997175,7.2153354,7.230953,7.2465706,7.2582836,7.2739015,6.6726236,6.0713453,5.466163,4.8648853,4.263607,4.591577,4.9234514,5.251421,5.5832953,5.911265,6.153338,6.3915067,6.6335793,6.871748,7.113821,7.394938,7.676055,7.9610763,8.242193,8.52331,8.718531,8.909846,9.101162,9.296382,9.487698,9.854712,10.221725,10.588739,10.955752,11.326671,10.48332,9.643873,8.804427,7.9649806,7.125534,6.5359693,5.9464045,5.35684,4.7633705,4.173806,7.437886,10.698062,13.962143,17.226223,20.486399,22.532305,24.578213,26.624119,28.66612,30.712029,30.290352,29.868677,29.443098,29.021421,28.599747,29.876486,31.14932,32.42606,33.698895,34.975636,31.465578,27.959425,24.453272,20.943214,17.437061,20.521538,23.606016,26.694399,29.778875,32.863354,27.73297,22.602585,17.4722,12.341816,7.211431,11.318862,15.426293,19.533724,23.641155,27.748587,22.739239,17.72989,12.720543,7.7111945,2.7018464,2.1708477,1.639849,1.1088502,0.58175594,0.05075723,0.339683,0.62860876,0.92143893,1.2103647,1.4992905,3.076669,4.650143,6.223617,7.800996,9.37447,7.5862536,5.794133,4.0059166,2.2137961,0.42557985,0.38653582,0.3513962,0.31235218,0.27330816,0.23816854,0.3357786,0.43729305,0.5388075,0.63641757,0.737932,0.63251317,0.5270943,0.42167544,0.31625658,0.21083772,0.19131571,0.1717937,0.15227169,0.13274968,0.113227665,0.12103647,0.13274968,0.14055848,0.15227169,0.1639849,0.14836729,0.13665408,0.12494087,0.113227665,0.10151446,0.1639849,0.22645533,0.28892577,0.3513962,0.41386664,0.39044023,0.3670138,0.3435874,0.3240654,0.30063897,0.28892577,0.28111696,0.26940376,0.26159495,0.24988174,0.21864653,0.19131571,0.16008049,0.12884527,0.10151446,0.09761006,0.093705654,0.093705654,0.08980125,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.21083772,0.21474212,0.21864653,0.21864653,0.22255093,0.22645533,0.32016098,0.41386664,0.5114767,0.60518235,0.698888,0.698888,0.6949836,0.6910792,0.6910792,0.6871748,0.6949836,0.7027924,0.7106012,0.71841,0.7262188,0.80821127,0.8941081,0.98000497,1.0659018,1.1517987,1.1869383,1.2181735,1.2533131,1.2884527,1.3235924,1.33921,1.3509232,1.3626363,1.3743496,1.3860629,1.6086137,1.8272603,2.0459068,2.2684577,2.4871042,2.690133,2.893162,3.096191,3.2992198,3.4983444,4.478349,5.4583545,6.4383593,7.4183645,8.398369,7.910319,7.4183645,6.930314,6.4383593,5.950309,6.3407493,6.735094,7.1294384,7.519879,7.914223,8.062591,8.210958,8.36323,8.511597,8.663869,9.491602,10.319335,11.143164,11.970898,12.798631,14.461906,16.121277,17.780647,19.44002,21.09939,20.958832,20.81437,20.67381,20.529346,20.388788,20.084246,19.783606,19.479063,19.178425,18.87388,18.787983,18.698183,18.612286,18.526388,18.436588,18.893402,19.346313,19.803127,20.256039,20.712854,1.1869383,1.3235924,1.4641509,1.6008049,1.737459,1.8741131,1.999054,2.1239948,2.2489357,2.3738766,2.4988174,2.4129205,2.3231194,2.2372224,2.1513257,2.0615244,2.1005683,2.135708,2.174752,2.2137961,2.2489357,2.5261483,2.7994564,3.076669,3.349977,3.6232853,3.8497405,4.0761957,4.298747,4.5252023,4.7516575,5.548156,6.348558,7.1489606,7.9493628,8.749765,7.137247,5.5247293,3.912211,2.2996929,0.6871748,0.58566034,0.48805028,0.38653582,0.28892577,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.113227665,0.1639849,0.21083772,0.26159495,0.31235218,0.28892577,0.26159495,0.23816854,0.21083772,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.21083772,0.23816854,0.26159495,0.28892577,0.31235218,0.3240654,0.3357786,0.3513962,0.3631094,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.58566034,1.0502841,1.5110037,1.9756275,2.436347,2.4871042,2.5378613,2.5886188,2.639376,2.6862288,2.2996929,1.9131571,1.5266213,1.1361811,0.74964523,0.6754616,0.60127795,0.5231899,0.44900626,0.37482262,0.39824903,0.42557985,0.44900626,0.47633708,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,1.1635119,2.260649,3.3616903,4.462732,5.563773,4.775084,3.9863946,3.2016098,2.4129205,1.6242313,2.3114061,2.998581,3.6857557,4.376835,5.0640097,5.735567,6.4110284,7.08649,7.7619514,8.437413,7.773665,7.113821,6.4500723,5.786324,5.12648,5.138193,5.1499066,5.1616197,5.173333,5.1889505,5.5871997,5.989353,6.387602,6.785851,7.1880045,7.1489606,7.113821,7.0747766,7.0357327,7.000593,6.7507114,6.5008297,6.250948,6.001066,5.7511845,6.0244927,6.3017054,6.575013,6.8483214,7.125534,8.175818,9.226103,10.276386,11.326671,12.373051,12.4511385,12.525322,12.599506,12.67369,12.751778,11.912332,11.076789,10.237343,9.4018,8.562354,7.137247,5.7121406,4.2870336,2.8619268,1.43682,2.8385005,4.2362766,5.6379566,7.0357327,8.437413,8.663869,8.886419,9.112875,9.339331,9.561881,10.4637985,11.361811,12.263727,13.16174,14.063657,12.775204,11.486752,10.198298,8.913751,7.6252975,9.999174,12.373051,14.750832,17.124708,19.498585,23.836376,28.174168,32.51196,36.849747,41.18754,44.11194,47.036335,49.96073,52.889034,55.81343,48.262318,40.7112,33.163994,25.612879,18.061766,17.49953,16.937298,16.375063,15.812829,15.250595,17.86264,20.474686,23.086731,25.698776,28.310822,32.699368,37.087917,41.476463,45.86111,50.249657,47.899208,45.548756,43.198307,40.85176,38.501312,36.40074,34.300175,32.199604,30.099037,27.998468,26.499178,24.999887,23.500597,22.001307,20.498112,19.26432,18.026625,16.788929,15.551234,14.313539,17.073952,19.838268,22.59868,25.362997,28.12341,26.90133,25.67535,24.449368,23.223385,22.001307,19.889025,17.776743,15.660558,13.548276,11.435994,10.87376,10.311526,9.749292,9.187058,8.624825,7.1880045,5.7511845,4.3143644,2.87364,1.43682,2.0615244,2.6862288,3.310933,3.9356375,4.564246,5.087436,5.610626,6.13772,6.66091,7.1880045,8.261715,9.339331,10.413041,11.486752,12.564366,11.213444,9.86252,8.511597,7.1606736,5.813655,5.735567,5.661383,5.5871997,5.5130157,5.4388323,6.114294,6.785851,7.461313,8.136774,8.812236,16.562475,24.312714,32.06295,39.81319,47.563427,48.473152,49.386784,50.300415,51.214043,52.12377,51.374126,50.62448,49.874836,49.12519,48.375546,39.172867,29.974096,20.775324,11.576552,2.3738766,2.0498111,1.7257458,1.4016805,1.0737107,0.74964523,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.21083772,0.30063897,0.38653582,0.47633708,0.5622339,0.63641757,0.7106012,0.78868926,0.8628729,0.93705654,2.6003318,4.263607,5.9268827,7.5862536,9.249529,11.888905,14.524376,17.163752,19.799223,22.4386,22.212145,21.98569,21.763138,21.536682,21.314133,19.088623,16.863113,14.637604,12.412095,10.186585,9.136301,8.086017,7.0357327,5.989353,4.939069,4.8765984,4.814128,4.7516575,4.689187,4.6267166,5.12648,5.6262436,6.126007,6.6257706,7.125534,6.0244927,4.9234514,3.8263142,2.7252727,1.6242313,3.0883822,4.548629,6.012779,7.47693,8.937177,8.289046,7.6370106,6.98888,6.336845,5.688714,6.036206,6.387602,6.7389984,7.08649,7.437886,7.437886,7.437886,7.437886,7.437886,7.437886,6.801469,6.1611466,5.5247293,4.8883114,4.251894,4.7009,5.1499066,5.5989127,6.0518236,6.5008297,6.7507114,7.000593,7.250475,7.5003567,7.7502384,7.9493628,8.148487,8.351517,8.550641,8.749765,9.300286,9.850807,10.401327,10.951848,11.498465,11.4516115,11.400854,11.350098,11.29934,11.248583,10.350571,9.448653,8.550641,7.648724,6.7507114,6.114294,5.473972,4.8375545,4.2011366,3.5608149,7.426173,11.287627,15.14908,19.014439,22.875893,24.539167,26.19854,27.861814,29.52509,31.188366,30.83697,30.485573,30.13808,29.786684,29.439194,30.83697,32.23865,33.636425,35.038105,36.435883,33.062477,29.689075,26.311768,22.938364,19.561056,21.025206,22.489357,23.949604,25.413754,26.874,22.911032,18.95197,14.989,11.0260315,7.0630636,9.839094,12.611219,15.387249,18.163279,20.93931,16.812357,12.689307,8.562354,4.4393053,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.42557985,0.78868926,1.1517987,1.5110037,1.8741131,3.8380275,5.7980375,7.7619514,9.725866,11.685876,9.448653,7.211431,4.9742084,2.736986,0.4997635,0.44900626,0.39824903,0.3513962,0.30063897,0.24988174,0.3513962,0.44900626,0.5505207,0.6481308,0.74964523,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.14836729,0.23816854,0.3240654,0.41386664,0.4997635,0.47633708,0.44900626,0.42557985,0.39824903,0.37482262,0.3631094,0.3513962,0.3357786,0.3240654,0.31235218,0.27330816,0.23816854,0.19912452,0.1639849,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.21083772,0.23816854,0.26159495,0.28892577,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.37482262,0.43729305,0.4997635,0.5622339,0.62470436,0.7262188,0.8238289,0.92534333,1.0268579,1.1244678,1.33921,1.5500476,1.7608855,1.9756275,2.1864653,2.3621633,2.5378613,2.7135596,2.8892577,3.0610514,4.2011366,5.337318,6.473499,7.6135845,8.749765,8.050878,7.348085,6.649197,5.950309,5.251421,5.423215,5.5989127,5.774611,5.950309,6.126007,6.375889,6.6257706,6.8756523,7.125534,7.375416,8.261715,9.151918,10.0382185,10.924518,11.810817,13.536563,15.262308,16.988054,18.7138,20.435642,20.400501,20.361458,20.326319,20.287273,20.24823,20.15062,20.049105,19.951496,19.849981,19.748466,19.412687,19.07691,18.737226,18.401447,18.061766,18.612286,19.162806,19.713327,20.263847,20.81437,1.2142692,1.3431144,1.475864,1.6086137,1.7413634,1.8741131,1.9834363,2.096664,2.2059872,2.3153105,2.4246337,2.3621633,2.2996929,2.2372224,2.174752,2.1122816,2.1513257,2.1864653,2.2255092,2.260649,2.2996929,2.5495746,2.7994564,3.049338,3.2992198,3.5491016,3.8770714,4.2050414,4.533011,4.860981,5.1889505,5.8370814,6.4891167,7.137247,7.7892823,8.437413,6.8951745,5.3529353,3.8106966,2.2684577,0.7262188,0.61689556,0.5114767,0.40215343,0.29673457,0.18741131,0.21083772,0.23426414,0.25378615,0.27721256,0.30063897,0.25769055,0.21474212,0.1717937,0.12884527,0.08589685,0.12103647,0.15227169,0.1835069,0.21864653,0.24988174,0.23426414,0.21474212,0.19912452,0.1796025,0.1639849,0.1639849,0.1678893,0.1717937,0.1717937,0.1756981,0.19131571,0.20693332,0.21864653,0.23426414,0.24988174,0.27721256,0.30454338,0.3318742,0.359205,0.38653582,0.38653582,0.38263142,0.37872702,0.37872702,0.37482262,0.30844778,0.23816854,0.1717937,0.10541886,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.5349031,0.92143893,1.3040704,1.6906061,2.0732377,2.1278992,2.1786566,2.233318,2.2840753,2.338737,2.0888553,1.8389735,1.5890918,1.33921,1.0893283,1.2923572,1.4992905,1.7023194,1.9092526,2.1122816,1.8819219,1.6476578,1.4133936,1.183034,0.94876975,0.76135844,0.5700427,0.37872702,0.19131571,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,1.0541886,2.0537157,3.057147,4.0605783,5.0640097,4.3729305,3.6818514,2.9907722,2.3035975,1.6125181,2.358259,3.1039999,3.8458362,4.591577,5.337318,5.7824197,6.2275214,6.6726236,7.1177254,7.562827,7.1333427,6.703859,6.2743745,5.840986,5.4115014,5.3841705,5.35684,5.3295093,5.3021784,5.2748475,5.5871997,5.899552,6.211904,6.524256,6.8366084,6.813182,6.79366,6.7702336,6.746807,6.7233806,6.5984397,6.473499,6.348558,6.223617,6.098676,6.3836975,6.6687193,6.9537406,7.238762,7.523783,8.433509,9.339331,10.249056,11.154878,12.0606985,12.056794,12.0489855,12.041177,12.033368,12.025558,11.170495,10.315431,9.460366,8.605303,7.7502384,6.504734,5.2592297,4.0137253,2.7682211,1.5266213,2.8892577,4.2557983,5.618435,6.984976,8.351517,8.683391,9.0152645,9.347139,9.679013,10.010887,11.506273,12.997755,14.489237,15.980719,17.476105,16.65618,15.836256,15.016331,14.196406,13.376482,15.313066,17.24965,19.186234,21.12672,23.063305,26.90133,30.735455,34.573483,38.41151,42.24954,44.763973,47.2745,49.788937,52.29947,54.813904,47.07928,39.34466,31.606136,23.871515,16.136894,15.793307,15.453624,15.110037,14.766449,14.426766,17.811884,21.200905,24.586021,27.975042,31.364063,34.26113,37.1621,40.063072,42.964043,45.86111,47.001194,48.137375,49.273556,50.413643,51.549824,46.08366,40.621403,35.15524,29.689075,24.226816,23.488884,22.750952,22.01302,21.275087,20.537155,21.661623,22.78609,23.914463,25.03893,26.163399,26.534317,26.90914,27.280058,27.650976,28.025799,26.526508,25.023314,23.524023,22.024733,20.525442,18.7138,16.898252,15.086611,13.274967,11.4633255,10.912805,10.362284,9.811763,9.261242,8.710721,7.348085,5.9815445,4.618908,3.252367,1.8858263,2.416825,2.9478238,3.4788225,4.0059166,4.5369153,5.153811,5.7707067,6.3915067,7.008402,7.6252975,8.480362,9.335425,10.19049,11.045554,11.900618,10.682445,9.464272,8.246098,7.0318284,5.813655,6.860035,7.9064145,8.956698,10.003078,11.0494585,11.615597,12.181735,12.743969,13.310107,13.8762455,21.868557,29.864773,37.86099,45.853302,53.849518,54.16187,54.470314,54.778763,55.091114,55.399563,52.237,49.074432,45.911865,42.749302,39.586735,32.22303,24.85933,17.491722,10.128019,2.7643168,2.377781,1.9912452,1.6086137,1.2220778,0.8394465,0.6910792,0.5466163,0.40215343,0.25769055,0.113227665,0.25378615,0.39824903,0.5388075,0.6832704,0.8238289,0.8667773,0.9058213,0.94486535,0.98390937,1.0268579,2.9361105,4.8492675,6.7624245,8.675582,10.588739,13.118792,15.652749,18.186707,20.716759,23.250715,22.62601,22.001307,21.376602,20.751898,20.12329,17.839214,15.555139,13.271063,10.983084,8.699008,7.8634663,7.0240197,6.1884775,5.349031,4.513489,4.60329,4.6930914,4.7828927,4.872694,4.9624953,5.2592297,5.55206,5.8487945,6.141625,6.4383593,5.840986,5.2475166,4.6540475,4.056674,3.4632049,4.5993857,5.735567,6.8756523,8.011833,9.151918,8.476458,7.8049,7.1333427,6.461786,5.786324,6.04011,6.2938967,6.5437784,6.7975645,7.0513506,6.949836,6.8483214,6.7507114,6.649197,6.551587,6.036206,5.520825,5.0054436,4.4900627,3.9746814,4.4002614,4.825841,5.251421,5.6730967,6.098676,6.3993154,6.6960497,6.9927845,7.289519,7.5862536,7.8400397,8.093826,8.343708,8.597494,8.85128,9.327617,9.803954,10.284196,10.760532,11.23687,11.154878,11.072885,10.990892,10.9089,10.826907,9.889851,8.956698,8.019642,7.08649,6.1494336,6.094772,6.04011,5.985449,5.930787,5.8761253,8.652155,11.428185,14.208119,16.98415,19.764084,21.02911,22.294136,23.559164,24.82419,26.089216,25.784672,25.484034,25.179491,24.87885,24.574308,25.901804,27.229301,28.556799,29.884295,31.211792,28.107792,25.003792,21.895887,18.791887,15.687888,17.202797,18.717705,20.232613,21.74752,23.262428,19.740658,16.222792,12.70102,9.183154,5.661383,7.882988,10.100689,12.322293,14.543899,16.761599,13.466284,10.167064,6.871748,3.5725281,0.27330816,0.23035973,0.1835069,0.14055848,0.093705654,0.05075723,0.39824903,0.74964523,1.1010414,1.4485333,1.7999294,3.3538816,4.903929,6.4578815,8.011833,9.561881,8.043069,6.5281606,5.009348,3.4905357,1.9756275,1.9717231,1.9639144,1.9600099,1.9561055,1.9482968,2.2957885,2.639376,2.9868677,3.330455,3.6740425,3.6506162,3.6232853,3.5998588,3.5764325,3.5491016,3.4436827,3.338264,3.2367494,3.1313305,3.0259118,2.4831998,1.9443923,1.4055848,0.8667773,0.3240654,0.27330816,0.21864653,0.1678893,0.113227665,0.062470436,0.13665408,0.20693332,0.28111696,0.3513962,0.42557985,0.44119745,0.46071947,0.47633708,0.4958591,0.5114767,0.4958591,0.47633708,0.46071947,0.44119745,0.42557985,0.37482262,0.3240654,0.27330816,0.22645533,0.1756981,0.1835069,0.19131571,0.19912452,0.20693332,0.21083772,0.23426414,0.25769055,0.28111696,0.30063897,0.3240654,0.3435874,0.3631094,0.38653582,0.40605783,0.42557985,0.42948425,0.43338865,0.44119745,0.44510186,0.44900626,0.46852827,0.48805028,0.5114767,0.5309987,0.5505207,0.5153811,0.48024148,0.44510186,0.40996224,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.40996224,0.44510186,0.48024148,0.5153811,0.5505207,0.62079996,0.6949836,0.76916724,0.8394465,0.9136301,1.0893283,1.2689307,1.4446288,1.6242313,1.7999294,1.9482968,2.096664,2.241127,2.3894942,2.5378613,3.4905357,4.4432096,5.395884,6.348558,7.3012323,6.9732623,6.6452928,6.3173227,5.989353,5.661383,6.001066,6.336845,6.676528,7.012306,7.348085,7.5862536,7.824422,8.062591,8.300759,8.538928,9.042596,9.546264,10.053836,10.557504,11.061172,12.579984,14.098797,15.613705,17.132517,18.651329,18.791887,18.928543,19.069101,19.20966,19.350218,19.20185,19.049578,18.90121,18.74894,18.600573,18.420969,18.241367,18.061766,17.878258,17.698656,18.471727,19.244799,20.01787,20.790941,21.564014,1.2376955,1.3665408,1.4914817,1.620327,1.7491722,1.8741131,1.9717231,2.0654287,2.1591344,2.2567444,2.35045,2.3114061,2.2762666,2.2372224,2.1981785,2.1630387,2.1981785,2.2372224,2.2762666,2.3114061,2.35045,2.5769055,2.7994564,3.0259118,3.2484627,3.474918,3.9044023,4.3338866,4.7633705,5.196759,5.6262436,6.126007,6.6257706,7.125534,7.6252975,8.125061,6.6531014,5.181142,3.7091823,2.233318,0.76135844,0.6481308,0.5309987,0.41777104,0.30063897,0.18741131,0.23426414,0.27721256,0.3240654,0.3670138,0.41386664,0.3513962,0.29283017,0.23426414,0.1717937,0.113227665,0.12884527,0.14055848,0.15617609,0.1717937,0.18741131,0.1756981,0.1678893,0.15617609,0.14836729,0.13665408,0.14055848,0.14836729,0.15227169,0.15617609,0.1639849,0.1678893,0.1717937,0.1756981,0.1835069,0.18741131,0.23035973,0.27330816,0.31625658,0.359205,0.39824903,0.39434463,0.39044023,0.38653582,0.37872702,0.37482262,0.31625658,0.25378615,0.19522011,0.13665408,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.48414588,0.78868926,1.097137,1.4055848,1.7140326,1.7686942,1.8233559,1.8780174,1.9326792,1.9873407,1.8741131,1.7608855,1.6515622,1.5383345,1.4251068,1.9092526,2.3933985,2.8814487,3.3655949,3.8497405,3.3616903,2.8697357,2.3816853,1.8897307,1.4016805,1.1205635,0.8394465,0.5583295,0.28111696,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.94096094,1.8467822,2.7526035,3.6584249,4.564246,3.970777,3.377308,2.7838387,2.194274,1.6008049,2.4012074,3.2055142,4.0059166,4.8102236,5.610626,5.8292727,6.044015,6.2587566,6.473499,6.688241,6.4891167,6.2938967,6.094772,5.8956475,5.700427,5.6340523,5.563773,5.4973984,5.4310236,5.3607445,5.5871997,5.813655,6.036206,6.262661,6.4891167,6.481308,6.473499,6.46569,6.4578815,6.4500723,6.4500723,6.4500723,6.4500723,6.4500723,6.4500723,6.746807,7.039637,7.336372,7.629202,7.9259367,8.691199,9.456462,10.221725,10.983084,11.748346,11.6585455,11.568744,11.478943,11.389141,11.29934,10.4286585,9.554072,8.683391,7.8088045,6.9381227,5.872221,4.806319,3.7443218,2.67842,1.6125181,2.9439192,4.271416,5.602817,6.9342184,8.261715,8.702912,9.14411,9.581403,10.0226,10.4637985,12.548749,14.633699,16.71865,18.8036,20.888552,20.53325,20.181856,19.83046,19.479063,19.123762,20.626957,22.126247,23.625538,25.124828,26.624119,29.962383,33.300648,36.638912,39.97327,43.311535,45.4121,47.512672,49.61324,51.713806,53.814377,45.892345,37.974216,30.052185,22.134056,14.212025,14.090988,13.966047,13.845011,13.723974,13.599033,17.761126,21.923218,26.089216,30.251308,34.413403,35.826794,37.236286,38.649677,40.063072,41.476463,46.099277,50.725994,55.34881,59.975525,64.598335,55.77048,46.938725,38.11087,29.279112,20.45126,20.474686,20.498112,20.525442,20.548868,20.5762,24.062832,27.549461,31.036093,34.52663,38.01326,35.994686,33.97611,31.961437,29.942862,27.924286,26.151686,24.375183,22.59868,20.826082,19.049578,17.538574,16.023666,14.512663,13.001659,11.486752,10.951848,10.413041,9.874233,9.339331,8.800523,7.5081654,6.2158084,4.9234514,3.631094,2.338737,2.7721257,3.2094188,3.6428072,4.0761957,4.513489,5.22409,5.930787,6.6413884,7.3519893,8.062591,8.699008,9.331521,9.967939,10.604357,11.23687,10.151445,9.066022,7.9805984,6.899079,5.813655,7.984503,10.151445,12.322293,14.493141,16.663988,17.1169,17.573715,18.026625,18.48344,18.936352,27.178545,35.416832,43.659027,51.897316,60.135605,59.84668,59.55385,59.261017,58.968185,58.675358,53.09987,47.524384,41.9489,36.373413,30.80183,25.26929,19.740658,14.208119,8.679486,3.1508527,2.7057507,2.260649,1.815547,1.3704453,0.92534333,0.76135844,0.59346914,0.42948425,0.26549935,0.10151446,0.29673457,0.4958591,0.6910792,0.8902037,1.0893283,1.0932326,1.097137,1.1010414,1.1088502,1.1127546,3.2757936,5.4388323,7.601871,9.761005,11.924045,14.352583,16.78112,19.205755,21.634293,24.062832,23.035973,22.01302,20.986162,19.96321,18.936352,16.59371,14.247164,11.900618,9.557977,7.211431,6.5867267,5.9620223,5.337318,4.7126136,4.087909,4.3299823,4.572055,4.814128,5.056201,5.298274,5.388075,5.481781,5.571582,5.661383,5.7511845,5.661383,5.571582,5.481781,5.388075,5.298274,6.114294,6.9264097,7.7385254,8.550641,9.362757,8.667773,7.9727893,7.277806,6.5828223,5.8878384,6.044015,6.196286,6.3524623,6.5086384,6.66091,6.461786,6.262661,6.0635366,5.8644123,5.661383,5.270943,4.8765984,4.4861584,4.0918136,3.7013733,4.0996222,4.5017757,4.900025,5.298274,5.700427,6.044015,6.3915067,6.735094,7.0786815,7.426173,7.7307167,8.03526,8.339804,8.644346,8.94889,9.354948,9.761005,10.163159,10.569217,10.975275,10.858143,10.744915,10.631687,10.514555,10.401327,9.4291315,8.460839,7.4886436,6.520352,5.548156,6.0791545,6.606249,7.1333427,7.660437,8.187531,9.882042,11.572648,13.263254,14.957765,16.64837,17.519053,18.38583,19.252607,20.119385,20.986162,20.732376,20.47859,20.2209,19.967113,19.713327,20.96664,22.223858,23.47717,24.734388,25.987701,23.153105,20.31851,17.483913,14.649317,11.810817,13.380386,14.946052,16.515621,18.081287,19.650856,16.574188,13.493614,10.416945,7.3402762,4.263607,5.9268827,7.5940623,9.257338,10.920613,12.587793,10.116306,7.648724,5.1772375,2.7057507,0.23816854,0.19912452,0.15617609,0.11713207,0.078088045,0.039044023,0.37482262,0.7106012,1.0502841,1.3860629,1.7257458,2.8658314,4.009821,5.153811,6.2938967,7.437886,6.6413884,5.840986,5.044488,4.2479897,3.4514916,3.4905357,3.5295796,3.5686235,3.611572,3.6506162,4.240181,4.829746,5.4193106,6.008875,6.5984397,6.676528,6.7507114,6.824895,6.899079,6.9732623,6.7663293,6.5554914,6.3446536,6.133816,5.9268827,4.83365,3.7404175,2.6471848,1.5539521,0.46071947,0.38263142,0.30063897,0.22255093,0.14055848,0.062470436,0.12103647,0.1756981,0.23426414,0.29283017,0.3513962,0.40996224,0.46852827,0.5309987,0.58956474,0.6481308,0.62860876,0.60518235,0.58175594,0.5583295,0.5388075,0.47633708,0.41386664,0.3513962,0.28892577,0.22645533,0.25378615,0.28111696,0.30844778,0.3357786,0.3631094,0.40605783,0.45291066,0.4958591,0.5427119,0.58566034,0.64032197,0.6910792,0.74574083,0.79649806,0.8511597,0.8238289,0.79649806,0.76916724,0.7418364,0.7106012,0.7262188,0.7418364,0.75745404,0.77307165,0.78868926,0.71841,0.6481308,0.57785153,0.5075723,0.43729305,0.43729305,0.43729305,0.43729305,0.43729305,0.43729305,0.44510186,0.45291066,0.46071947,0.46852827,0.47633708,0.5192855,0.5661383,0.60908675,0.6559396,0.698888,0.8433509,0.98390937,1.1283722,1.2689307,1.4133936,1.53443,1.6515622,1.7725986,1.893635,2.0107672,2.7799344,3.5491016,4.3143644,5.083532,5.8487945,5.8956475,5.938596,5.985449,6.028397,6.0752497,6.575013,7.0747766,7.57454,8.074304,8.574067,8.800523,9.026978,9.249529,9.475985,9.698535,9.823476,9.944512,10.069453,10.19049,10.311526,11.623405,12.93138,14.243259,15.551234,16.863113,17.17937,17.495626,17.815788,18.132044,18.448301,18.249176,18.05005,17.850927,17.651802,17.448774,17.429253,17.405825,17.382399,17.358973,17.33945,18.33117,19.326792,20.322414,21.318037,22.31366,1.261122,1.3860629,1.5070993,1.6281357,1.7530766,1.8741131,1.9561055,2.0341935,2.1161861,2.194274,2.2762666,2.260649,2.2489357,2.2372224,2.2255092,2.2137961,2.2489357,2.2879796,2.3231194,2.3621633,2.4012074,2.6003318,2.7994564,2.998581,3.2016098,3.4007344,3.9317331,4.466636,4.997635,5.5286336,6.0635366,6.4110284,6.7624245,7.113821,7.461313,7.812709,6.4110284,5.009348,3.6037633,2.2020829,0.80040246,0.679366,0.5544251,0.43338865,0.30844778,0.18741131,0.25378615,0.3240654,0.39044023,0.45681506,0.5231899,0.44900626,0.3709182,0.29283017,0.21474212,0.13665408,0.13665408,0.13274968,0.12884527,0.12884527,0.12494087,0.12103647,0.12103647,0.11713207,0.113227665,0.113227665,0.12103647,0.12884527,0.13665408,0.14055848,0.14836729,0.14446288,0.14055848,0.13665408,0.12884527,0.12494087,0.1835069,0.23816854,0.29673457,0.3553006,0.41386664,0.40605783,0.39824903,0.39044023,0.38263142,0.37482262,0.3240654,0.26940376,0.21864653,0.1639849,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.42948425,0.659844,0.8902037,1.1205635,1.3509232,1.4055848,1.4641509,1.5227169,1.5812829,1.6359446,1.6632754,1.6867018,1.7140326,1.737459,1.7608855,2.5261483,3.2914112,4.056674,4.8219366,5.5871997,4.841459,4.0918136,3.3460727,2.5964274,1.8506867,1.4797685,1.1088502,0.7418364,0.3709182,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.8316377,1.639849,2.4480603,3.2562714,4.0605783,3.5686235,3.0727646,2.5769055,2.0810463,1.5890918,2.4480603,3.3070288,4.165997,5.02887,5.8878384,5.872221,5.8566036,5.840986,5.8292727,5.813655,5.8487945,5.883934,5.919074,5.9542136,5.989353,5.8800297,5.7707067,5.6652875,5.5559645,5.4505453,5.5871997,5.7238536,5.8644123,6.001066,6.13772,6.1455293,6.153338,6.1611466,6.168956,6.1767645,6.3017054,6.426646,6.551587,6.676528,6.801469,7.1060123,7.4105554,7.715099,8.019642,8.324185,8.94889,9.56969,10.194394,10.815194,11.435994,11.2642,11.092407,10.920613,10.748819,10.573121,9.686822,8.796618,7.9064145,7.016211,6.126007,5.239708,4.3534083,3.4710135,2.5847144,1.698415,2.9946766,4.290938,5.5832953,6.8795567,8.175818,8.722435,9.269051,9.815667,10.366188,10.912805,13.591225,16.26574,18.94416,21.62258,24.300999,24.414227,24.531359,24.644587,24.761719,24.874947,25.936945,26.998941,28.06094,29.12684,30.188839,33.023434,35.861935,38.700436,41.538937,44.37353,46.064137,47.75084,49.437542,51.124245,52.810944,44.70931,36.60377,28.498232,20.392693,12.287154,12.384764,12.482374,12.579984,12.677594,12.775204,17.714273,22.649437,27.588507,32.52367,37.462738,37.388557,37.314373,37.236286,37.1621,37.087917,45.201263,53.310707,61.424057,69.53741,77.65075,65.4534,53.259953,41.0665,28.86915,16.675701,17.464392,18.249176,19.037865,19.826555,20.61134,26.464039,32.31283,38.16163,44.014328,49.86312,45.45505,41.04698,36.638912,32.23084,27.826675,25.776863,23.723148,21.673336,19.623526,17.573715,16.36335,15.14908,13.938716,12.724447,11.514082,10.986988,10.4637985,9.936704,9.413514,8.886419,7.6682463,6.446168,5.2279944,4.0059166,2.787743,3.1274261,3.4671092,3.8067923,4.1464753,4.4861584,5.290465,6.0908675,6.8951745,7.6955767,8.499884,8.913751,9.331521,9.745388,10.159255,10.573121,9.6243515,8.671678,7.719003,6.7663293,5.813655,9.105066,12.396477,15.6917925,18.983204,22.274614,22.618202,22.965694,23.309282,23.656773,24.00036,32.484627,40.96889,49.45706,57.94133,66.4256,65.53149,64.63348,63.73937,62.84526,61.95115,53.96274,45.974335,37.98593,30.001427,22.01302,18.315552,14.621986,10.928422,7.230953,3.5373883,3.0337205,2.5261483,2.0224805,1.5188124,1.0112402,0.8277333,0.6442264,0.45681506,0.27330816,0.08589685,0.339683,0.59346914,0.8433509,1.097137,1.3509232,1.319688,1.2884527,1.261122,1.2298868,1.1986516,3.611572,6.0244927,8.437413,10.850334,13.263254,15.586374,17.905588,20.228708,22.551826,24.874947,23.44984,22.024733,20.599627,19.174519,17.749413,15.344301,12.939189,10.534078,8.128965,5.7238536,5.3138914,4.900025,4.4861584,4.0761957,3.6623292,4.056674,4.4510183,4.8492675,5.2436123,5.6379566,5.520825,5.407597,5.2943697,5.1772375,5.0640097,5.477876,5.891743,6.3056097,6.7233806,7.137247,7.6252975,8.113348,8.601398,9.089449,9.573594,8.859089,8.140678,7.422269,6.703859,5.989353,6.044015,6.1025805,6.1611466,6.2158084,6.2743745,5.9737353,5.6730967,5.376362,5.0757227,4.775084,4.50568,4.2362766,3.9668727,3.6935644,3.4241607,3.7989833,4.173806,4.548629,4.9234514,5.298274,5.6926184,6.083059,6.477403,6.871748,7.262188,7.621393,7.9766936,8.335898,8.691199,9.050405,9.382278,9.714153,10.046027,10.381805,10.71368,10.565312,10.416945,10.268578,10.124115,9.975748,8.968412,7.9649806,6.9615493,5.9542136,4.950782,6.0596323,7.168483,8.281238,9.390087,10.498938,11.108025,11.713207,12.322293,12.93138,13.536563,14.008995,14.477524,14.946052,15.418485,15.8870125,15.680079,15.473146,15.266212,15.059279,14.848442,16.031475,17.21451,18.397543,19.580578,20.76361,18.19842,15.633226,13.068034,10.502842,7.9376497,9.557977,11.178304,12.798631,14.418958,16.039284,13.403813,10.768341,8.13287,5.4973984,2.8619268,3.970777,5.083532,6.192382,7.3012323,8.413987,6.7702336,5.12648,3.4866312,1.8428779,0.19912452,0.1639849,0.12884527,0.093705654,0.058566034,0.023426414,0.3513962,0.6754616,0.999527,1.3235924,1.6515622,2.3816853,3.1157131,3.8458362,4.579864,5.3138914,5.2358036,5.1577153,5.0796275,5.001539,4.9234514,5.009348,5.095245,5.181142,5.263134,5.349031,6.184573,7.0201154,7.8556576,8.691199,9.526741,9.698535,9.874233,10.049932,10.22563,10.401327,10.085071,9.768814,9.456462,9.140205,8.823949,7.180196,5.5364423,3.8887846,2.2450314,0.60127795,0.49195468,0.38653582,0.27721256,0.1717937,0.062470436,0.10541886,0.14836729,0.19131571,0.23426414,0.27330816,0.37872702,0.48024148,0.58175594,0.6832704,0.78868926,0.76135844,0.7340276,0.7066968,0.679366,0.6481308,0.57394713,0.4997635,0.42557985,0.3513962,0.27330816,0.3240654,0.3709182,0.41777104,0.46462387,0.5114767,0.58175594,0.6481308,0.7145056,0.78088045,0.8511597,0.93315214,1.0190489,1.1049459,1.1908426,1.2767396,1.2142692,1.1557031,1.0932326,1.0346665,0.97610056,0.98390937,0.9956226,1.0034313,1.0151446,1.0268579,0.92143893,0.8160201,0.7106012,0.60518235,0.4997635,0.4997635,0.4997635,0.4997635,0.4997635,0.4997635,0.48024148,0.46071947,0.44119745,0.42167544,0.39824903,0.41777104,0.43338865,0.45291066,0.46852827,0.48805028,0.59346914,0.7027924,0.80821127,0.91753453,1.0268579,1.116659,1.2103647,1.3040704,1.3938715,1.4875772,2.069333,2.6510892,3.2367494,3.8185053,4.4002614,4.8180323,5.2358036,5.6535745,6.0713453,6.4891167,7.1489606,7.812709,8.476458,9.136301,9.80005,10.010887,10.22563,10.436467,10.651209,10.862047,10.604357,10.342762,10.081166,9.823476,9.561881,10.666827,11.767868,12.86891,13.973856,15.074897,15.570756,16.066616,16.55857,17.054428,17.550287,17.300406,17.050524,16.800642,16.55076,16.300879,16.43363,16.570284,16.706938,16.839687,16.976341,18.194515,19.408783,20.626957,21.84513,23.063305,1.2884527,1.4055848,1.5227169,1.639849,1.756981,1.8741131,1.9404879,2.0068626,2.069333,2.135708,2.1981785,2.2137961,2.2255092,2.2372224,2.2489357,2.260649,2.2996929,2.338737,2.3738766,2.4129205,2.4480603,2.6237583,2.7994564,2.9751544,3.1508527,3.3265507,3.959064,4.5954814,5.2318993,5.8644123,6.5008297,6.699954,6.899079,7.098203,7.3012323,7.5003567,6.168956,4.83365,3.5022488,2.1708477,0.8394465,0.7066968,0.57785153,0.44900626,0.31625658,0.18741131,0.27721256,0.3670138,0.45681506,0.5466163,0.63641757,0.5427119,0.44900626,0.3513962,0.25769055,0.1639849,0.14055848,0.12103647,0.10151446,0.08199245,0.062470436,0.06637484,0.07418364,0.078088045,0.08199245,0.08589685,0.09761006,0.10932326,0.11713207,0.12884527,0.13665408,0.12103647,0.10932326,0.093705654,0.078088045,0.062470436,0.13665408,0.20693332,0.28111696,0.3513962,0.42557985,0.41386664,0.40605783,0.39434463,0.38653582,0.37482262,0.3318742,0.28502136,0.23816854,0.19522011,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.046852827,0.08980125,0.13665408,0.1796025,0.22645533,0.37872702,0.5309987,0.6832704,0.8355421,0.9878138,1.0463798,1.1088502,1.1674163,1.2259823,1.2884527,1.4485333,1.6125181,1.7765031,1.9365835,2.1005683,3.1430438,4.1894236,5.2358036,6.278279,7.3246584,6.321227,5.3138914,4.31046,3.3031244,2.2996929,1.8389735,1.3782539,0.92143893,0.46071947,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.7223144,1.4329157,2.1435168,2.854118,3.5608149,3.1664703,2.7682211,2.3699722,1.9717231,1.5734742,2.4910088,3.408543,4.3260775,5.2436123,6.1611466,5.919074,5.6730967,5.4271193,5.181142,4.939069,5.2045684,5.473972,5.7394714,6.008875,6.2743745,6.126007,5.9815445,5.833177,5.6848097,5.5364423,5.5871997,5.6379566,5.688714,5.735567,5.786324,5.8097506,5.833177,5.8566036,5.8761253,5.899552,6.1494336,6.3993154,6.649197,6.899079,7.1489606,7.465217,7.7814736,8.093826,8.410083,8.726339,9.20658,9.686822,10.163159,10.6434,11.123642,10.869856,10.61607,10.358379,10.104593,9.850807,8.941081,8.03526,7.125534,6.2197127,5.3138914,4.607195,3.9044023,3.1977055,2.4910088,1.7882162,3.049338,4.3065557,5.5676775,6.8287997,8.086017,8.741957,9.397896,10.053836,10.705871,11.361811,14.633699,17.901684,21.173573,24.441559,27.713448,28.295202,28.876959,29.458715,30.044374,30.626131,31.250835,31.87554,32.500244,33.12495,33.749653,36.08839,38.42322,40.76196,43.100697,45.439434,46.71227,47.98901,49.261845,50.53858,51.811417,43.522373,35.233326,26.940376,18.651329,10.362284,10.67854,10.998701,11.314958,11.631214,11.951375,17.663515,23.375656,29.087797,34.79994,40.512077,38.950317,37.388557,35.826794,34.26113,32.699368,44.299347,55.899326,67.499306,79.09929,90.699265,75.14022,59.581177,44.01823,28.459188,12.900145,14.450192,16.00024,17.550287,19.100336,20.650383,28.861341,37.076202,45.287163,53.502026,61.712982,54.915417,48.117855,41.32029,34.522724,27.72516,25.398136,23.075018,20.747993,18.424873,16.101755,15.188125,14.274494,13.360865,12.4511385,11.537509,11.0260315,10.510651,9.999174,9.487698,8.976221,7.8283267,6.6804323,5.532538,4.3846436,3.2367494,3.4827268,3.7287042,3.970777,4.2167544,4.462732,5.35684,6.250948,7.1489606,8.043069,8.937177,9.132397,9.327617,9.522837,9.718058,9.913278,9.093353,8.273428,7.453504,6.6335793,5.813655,10.229534,14.641508,19.057388,23.473267,27.889145,28.12341,28.357674,28.591938,28.826202,29.064371,37.794613,46.520954,55.251198,63.98144,72.711685,71.21629,69.71701,68.22162,66.72233,65.226944,54.825615,44.42429,34.02296,23.625538,13.224211,11.365715,9.503315,7.6448197,5.786324,3.9239242,3.3616903,2.795552,2.2294137,1.6632754,1.1010414,0.8941081,0.6910792,0.48414588,0.28111696,0.07418364,0.38263142,0.6910792,0.9956226,1.3040704,1.6125181,1.5461433,1.4836729,1.4172981,1.3509232,1.2884527,3.951255,6.6140575,9.276859,11.935758,14.59856,16.816261,19.03396,21.251661,23.469362,25.687063,23.863707,22.036446,20.21309,18.38583,16.562475,14.098797,11.631214,9.167537,6.703859,4.2362766,4.037152,3.8380275,3.638903,3.435874,3.2367494,3.7833657,4.3338866,4.8805027,5.4271193,5.9737353,5.6535745,5.3334136,5.0132523,4.6930914,4.376835,5.2943697,6.2158084,7.1333427,8.054782,8.976221,9.136301,9.300286,9.464272,9.6243515,9.788337,9.0465,8.308568,7.5667315,6.8287997,6.086963,6.0479193,6.008875,5.9659266,5.9268827,5.8878384,5.4856853,5.087436,4.689187,4.2870336,3.8887846,3.7404175,3.59205,3.4436827,3.2992198,3.1508527,3.4983444,3.8497405,4.2011366,4.548629,4.900025,5.3412223,5.7785153,6.2197127,6.66091,7.098203,7.5081654,7.918128,8.32809,8.741957,9.151918,9.40961,9.671205,9.928895,10.19049,10.44818,10.268578,10.088976,9.909373,9.729771,9.550168,8.511597,7.4691215,6.4305506,5.388075,4.349504,6.044015,7.734621,9.4291315,11.119738,12.814248,12.334006,11.85767,11.381332,10.901091,10.424754,10.498938,10.569217,10.6434,10.71368,10.787864,10.627783,10.467703,10.307622,10.147541,9.987461,11.096312,12.209065,13.317916,14.426766,15.535617,13.243732,10.947944,8.652155,6.356367,4.0605783,5.735567,7.406651,9.081639,10.752724,12.423808,10.2334385,8.039165,5.8487945,3.6545205,1.4641509,2.018576,2.5730011,3.1274261,3.6818514,4.2362766,3.4241607,2.6081407,1.7921207,0.97610056,0.1639849,0.13274968,0.10151446,0.07418364,0.042948425,0.011713207,0.3240654,0.63641757,0.94876975,1.261122,1.5734742,1.8975395,2.2216048,2.541766,2.8658314,3.1859922,3.8302186,4.4705405,5.114767,5.758993,6.3993154,6.5281606,6.66091,6.7897553,6.918601,7.0513506,8.128965,9.2104845,10.2881,11.369619,12.4511385,12.724447,13.001659,13.274967,13.548276,13.825488,13.403813,12.986042,12.564366,12.146595,11.72492,9.526741,7.328563,5.134289,2.9361105,0.737932,0.60127795,0.46852827,0.3318742,0.19912452,0.062470436,0.08980125,0.11713207,0.14446288,0.1717937,0.19912452,0.3435874,0.48805028,0.63641757,0.78088045,0.92534333,0.8941081,0.8589685,0.8277333,0.79649806,0.76135844,0.6754616,0.58566034,0.4997635,0.41386664,0.3240654,0.39434463,0.46071947,0.5270943,0.59346914,0.6637484,0.75354964,0.8433509,0.93315214,1.0229534,1.1127546,1.2298868,1.3470187,1.4641509,1.5812829,1.698415,1.6086137,1.5149081,1.4212024,1.3314011,1.2376955,1.2415999,1.2494087,1.2533131,1.2572175,1.261122,1.1205635,0.98390937,0.8433509,0.7027924,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.5153811,0.46852827,0.42167544,0.3709182,0.3240654,0.31625658,0.30454338,0.29673457,0.28502136,0.27330816,0.3474918,0.42167544,0.49195468,0.5661383,0.63641757,0.7027924,0.76916724,0.8316377,0.8980125,0.96438736,1.358732,1.756981,2.15523,2.5534792,2.951728,3.7404175,4.5291066,5.3217,6.1103897,6.899079,7.726812,8.550641,9.37447,10.198298,11.0260315,11.225157,11.424281,11.623405,11.826434,12.025558,11.381332,10.741011,10.096785,9.456462,8.812236,9.706344,10.604357,11.498465,12.392572,13.286681,13.958238,14.633699,15.305257,15.976814,16.64837,16.351637,16.050997,15.750359,15.449719,15.14908,15.441911,15.734741,16.02757,16.320402,16.613232,18.053955,19.490776,20.931501,22.372225,23.81295,1.3118792,1.4251068,1.5383345,1.6515622,1.7608855,1.8741131,1.9248703,1.9756275,2.0263848,2.0732377,2.1239948,2.1630387,2.1981785,2.2372224,2.2762666,2.3114061,2.35045,2.3855898,2.4246337,2.463678,2.4988174,2.6510892,2.7994564,2.951728,3.1000953,3.2484627,3.9863946,4.7243266,5.462259,6.2001905,6.9381227,6.98888,7.0357327,7.08649,7.137247,7.1880045,5.9268827,4.661856,3.4007344,2.135708,0.8745861,0.737932,0.60127795,0.46071947,0.3240654,0.18741131,0.30063897,0.41386664,0.5231899,0.63641757,0.74964523,0.63641757,0.5231899,0.41386664,0.30063897,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.42557985,0.41386664,0.39824903,0.38653582,0.37482262,0.3357786,0.30063897,0.26159495,0.22645533,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.3240654,0.39824903,0.47633708,0.5505207,0.62470436,0.6871748,0.74964523,0.81211567,0.8745861,0.93705654,1.2376955,1.5383345,1.8389735,2.135708,2.436347,3.7638438,5.087436,6.4110284,7.7385254,9.062118,7.800996,6.5359693,5.2748475,4.0137253,2.7486992,2.1981785,1.6515622,1.1010414,0.5505207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.61299115,1.2259823,1.8389735,2.4480603,3.0610514,2.7643168,2.463678,2.1630387,1.8623998,1.5617609,2.5378613,3.513962,4.4861584,5.462259,6.4383593,5.9620223,5.4856853,5.0132523,4.5369153,4.0605783,4.564246,5.0640097,5.563773,6.0635366,6.5633,6.375889,6.1884775,6.001066,5.813655,5.6262436,5.5871997,5.548156,5.5130157,5.473972,5.4388323,5.473972,5.5130157,5.548156,5.5871997,5.6262436,6.001066,6.375889,6.7507114,7.125534,7.5003567,7.824422,8.148487,8.476458,8.800523,9.124588,9.464272,9.80005,10.135828,10.475512,10.81129,10.475512,10.135828,9.80005,9.464272,9.124588,8.1992445,7.2739015,6.348558,5.423215,4.5017757,3.9746814,3.4514916,2.9243972,2.4012074,1.8741131,3.1000953,4.3260775,5.548156,6.774138,8.00012,8.761478,9.526741,10.2881,11.0494585,11.810817,15.676175,19.537628,23.399082,27.26444,31.125895,32.176178,33.226463,34.27675,35.323128,36.373413,36.56082,36.748234,36.935646,37.12306,37.314373,39.14944,40.988415,42.823483,44.662457,46.50143,47.364304,48.22327,49.086143,49.949017,50.81189,42.339336,33.86288,25.386423,16.91387,8.437413,8.976221,9.511124,10.049932,10.588739,11.123642,17.612759,24.097971,30.587088,37.076202,43.561417,40.512077,37.462738,34.413403,31.364063,28.310822,43.401337,58.487946,73.574554,88.66116,103.75168,84.82704,65.902405,46.97386,28.049225,9.124588,11.435994,13.751305,16.062712,18.374117,20.689428,31.262548,41.83567,52.412697,62.985817,73.56284,64.375786,55.188725,46.001667,36.810703,27.623646,25.023314,22.426888,19.826555,17.226223,14.625891,14.012899,13.399908,12.786918,12.173926,11.560935,11.061172,10.561408,10.061645,9.561881,9.062118,7.988407,6.910792,5.8370814,4.7633705,3.6857557,3.8380275,3.9863946,4.138666,4.2870336,4.4393053,5.423215,6.4110284,7.3988423,8.386656,9.37447,9.351044,9.323712,9.300286,9.276859,9.249529,8.562354,7.8751793,7.1880045,6.5008297,5.813655,11.350098,16.88654,22.426888,27.96333,33.49977,33.624714,33.749653,33.874596,33.999535,34.124477,43.100697,52.073013,61.049232,70.02545,79.00168,76.90111,74.80054,72.69997,70.5994,68.49883,55.688488,42.87424,30.063898,17.24965,4.4393053,4.4119744,4.388548,4.3612175,4.337791,4.3143644,3.6857557,3.0610514,2.436347,1.8116426,1.1869383,0.96438736,0.737932,0.5114767,0.28892577,0.062470436,0.42557985,0.78868926,1.1517987,1.5110037,1.8741131,1.7765031,1.6749885,1.5734742,1.475864,1.3743496,4.2870336,7.1997175,10.112402,13.025085,15.93777,18.05005,20.162333,22.274614,24.386896,26.499178,24.273668,22.048159,19.826555,17.601046,15.375536,12.849388,10.323239,7.800996,5.2748475,2.7486992,2.7643168,2.77603,2.787743,2.7994564,2.8111696,3.513962,4.21285,4.911738,5.610626,6.3134184,5.786324,5.263134,4.73604,4.21285,3.6857557,5.1108627,6.5359693,7.9610763,9.386183,10.81129,10.651209,10.487225,10.323239,10.163159,9.999174,9.237816,8.476458,7.7111945,6.949836,6.1884775,6.0518236,5.911265,5.774611,5.6379566,5.5013027,5.001539,4.5017757,3.998108,3.4983444,2.998581,2.9751544,2.951728,2.9243972,2.900971,2.87364,3.2016098,3.5256753,3.8497405,4.173806,4.5017757,4.985922,5.473972,5.9620223,6.4500723,6.9381227,7.3988423,7.8634663,8.324185,8.78881,9.249529,9.43694,9.6243515,9.811763,9.999174,10.186585,9.975748,9.761005,9.550168,9.339331,9.124588,8.050878,6.9732623,5.899552,4.825841,3.7482262,6.0244927,8.300759,10.573121,12.849388,15.125654,13.563893,11.998228,10.436467,8.874706,7.3129454,6.98888,6.66091,6.336845,6.012779,5.688714,5.575486,5.462259,5.349031,5.2358036,5.12648,6.1611466,7.1997175,8.238289,9.276859,10.311526,8.289046,6.262661,4.2362766,2.2137961,0.18741131,1.9131571,3.638903,5.3607445,7.08649,8.812236,7.0630636,5.3138914,3.5608149,1.8116426,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.30063897,0.60127795,0.9019169,1.1986516,1.4992905,1.4133936,1.3235924,1.2376955,1.1517987,1.0619974,2.4246337,3.78727,5.1499066,6.5125427,7.8751793,8.050878,8.226576,8.398369,8.574067,8.749765,10.073358,11.400854,12.724447,14.051944,15.375536,15.750359,16.125181,16.500004,16.874826,17.24965,16.72646,16.199366,15.676175,15.14908,14.625891,11.873287,9.124588,6.375889,3.6232853,0.8745861,0.7106012,0.5505207,0.38653582,0.22645533,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.31235218,0.4997635,0.6871748,0.8745861,1.0619974,1.0268579,0.9878138,0.94876975,0.9136301,0.8745861,0.77307165,0.6754616,0.57394713,0.47633708,0.37482262,0.46071947,0.5505207,0.63641757,0.7262188,0.81211567,0.92534333,1.038571,1.1517987,1.261122,1.3743496,1.5266213,1.6749885,1.8233559,1.9756275,2.1239948,1.999054,1.8741131,1.7491722,1.6242313,1.4992905,1.4992905,1.4992905,1.4992905,1.4992905,1.4992905,1.3235924,1.1517987,0.97610056,0.80040246,0.62470436,0.62470436,0.62470436,0.62470436,0.62470436,0.62470436,0.5505207,0.47633708,0.39824903,0.3240654,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,0.10151446,0.13665408,0.1756981,0.21083772,0.24988174,0.28892577,0.3240654,0.3631094,0.39824903,0.43729305,0.6481308,0.8628729,1.0737107,1.2884527,1.4992905,2.6628022,3.8263142,4.985922,6.1494336,7.3129454,8.300759,9.288573,10.276386,11.2642,12.24811,12.439425,12.626837,12.814248,13.001659,13.189071,12.162213,11.139259,10.112402,9.089449,8.062591,8.749765,9.43694,10.124115,10.81129,11.498465,12.349625,13.200784,14.051944,14.899199,15.750359,15.398962,15.051471,14.700074,14.348679,14.001186,14.450192,14.899199,15.348206,15.801116,16.250122,17.913397,19.576674,21.236044,22.899319,24.562595,1.3509232,1.456342,1.5656652,1.6710842,1.7804074,1.8858263,1.9365835,1.9834363,2.0302892,2.077142,2.1239948,2.1708477,2.2216048,2.2684577,2.3153105,2.3621633,2.397303,2.4324427,2.4675822,2.5027218,2.5378613,2.67842,2.822883,2.9634414,3.1079042,3.2484627,3.951255,4.650143,5.349031,6.0518236,6.7507114,6.7663293,6.785851,6.801469,6.8209906,6.8366084,5.704332,4.572055,3.4397783,2.3075018,1.175225,1.0346665,0.8941081,0.75354964,0.61689556,0.47633708,0.5114767,0.5466163,0.58175594,0.61689556,0.6481308,0.5544251,0.45681506,0.359205,0.26159495,0.1639849,0.12884527,0.09761006,0.06637484,0.031235218,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.058566034,0.07027924,0.078088045,0.08980125,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.07027924,0.14055848,0.21083772,0.28111696,0.3513962,0.3435874,0.3357786,0.3279698,0.32016098,0.31235218,0.28111696,0.24597734,0.21474212,0.1835069,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.60127795,0.8941081,1.183034,1.4719596,1.7608855,1.7921207,1.8233559,1.8506867,1.8819219,1.9131571,2.0263848,2.135708,2.2489357,2.3621633,2.475391,3.6232853,4.7711797,5.919074,7.0630636,8.210958,7.2426662,6.2743745,5.3021784,4.3338866,3.3616903,2.7838387,2.2059872,1.6281357,1.0541886,0.47633708,0.46071947,0.44510186,0.42948425,0.41386664,0.39824903,0.48414588,0.5700427,0.6559396,0.7418364,0.8238289,1.1517987,1.475864,1.7999294,2.1239948,2.4480603,2.358259,2.2684577,2.1786566,2.0888553,1.999054,2.854118,3.7052777,4.5564375,5.4115014,6.262661,5.891743,5.5169206,5.1460023,4.7711797,4.4002614,4.8375545,5.2748475,5.7121406,6.1494336,6.5867267,6.473499,6.356367,6.2431393,6.126007,6.012779,5.852699,5.6926184,5.532538,5.3724575,5.212377,5.196759,5.181142,5.169429,5.153811,5.138193,5.5676775,5.997162,6.426646,6.8561306,7.2856145,7.629202,7.968885,8.308568,8.648251,8.987934,9.323712,9.663396,9.999174,10.338858,10.674636,10.350571,10.0265045,9.698535,9.37447,9.050405,8.378847,7.703386,7.0318284,6.3602715,5.688714,5.1772375,4.6657605,4.1581883,3.6467118,3.1391394,4.1113358,5.083532,6.055728,7.027924,8.00012,8.695104,9.390087,10.085071,10.780055,11.475039,15.453624,19.428307,23.40689,27.385477,31.364063,33.620808,35.877552,38.134296,40.39104,42.65169,42.382286,42.116787,41.84738,41.581882,41.31248,41.913757,42.51113,43.11241,43.713688,44.31106,45.166126,46.017284,46.868446,47.723507,48.57467,40.590164,32.605663,24.62116,16.636658,8.648251,9.042596,9.43694,9.82738,10.221725,10.612165,16.995863,23.375656,29.759354,36.14305,42.52675,39.75072,36.978592,34.206467,31.434343,28.662216,41.289055,53.911987,66.538826,79.16176,91.78859,75.3003,58.81201,42.32372,25.83543,9.351044,11.908427,14.465811,17.023193,19.580578,22.13796,30.950197,39.762432,48.57467,57.386906,66.19914,58.183403,50.17157,42.15583,34.140095,26.124355,25.378614,24.636778,23.891037,23.145296,22.399555,20.51373,18.631807,16.745981,14.860155,12.974329,13.083652,13.189071,13.298394,13.403813,13.513136,11.553126,9.597021,7.6409154,5.6809053,3.7247996,3.8341231,3.9434462,4.056674,4.165997,4.2753205,5.153811,6.028397,6.9068875,7.785378,8.663869,8.546737,8.433509,8.316377,8.203149,8.086017,7.9337454,7.7775693,7.621393,7.4691215,7.3129454,11.221252,15.133463,19.041769,22.953981,26.862288,28.525562,30.188839,31.84821,33.511486,35.17476,41.851288,48.52391,55.20044,61.87697,68.54959,66.20695,63.864307,61.521667,59.179024,56.836384,46.720078,36.607674,26.49137,16.378967,6.262661,5.716045,5.169429,4.618908,4.0722914,3.5256753,3.3187418,3.1118085,2.900971,2.6940374,2.4871042,2.018576,1.5461433,1.077615,0.60908675,0.13665408,0.7418364,1.3470187,1.9522011,2.5573835,3.1625657,3.0610514,2.9556324,2.854118,2.7526035,2.6510892,5.337318,8.023546,10.71368,13.399908,16.086138,17.26917,18.448301,19.62743,20.80656,21.98569,20.076437,18.167183,16.25793,14.348679,12.439425,10.545791,8.652155,6.75852,4.8687897,2.9751544,2.8306916,2.6862288,2.541766,2.3933985,2.2489357,3.1039999,3.9551594,4.806319,5.661383,6.5125427,5.9425,5.3724575,4.802415,4.2323723,3.6623292,5.6262436,7.5940623,9.557977,11.521891,13.4858055,12.790822,12.091934,11.393045,10.698062,9.999174,9.218294,8.441318,7.660437,6.8795567,6.098676,5.8761253,5.64967,5.423215,5.2006636,4.9742084,4.552533,4.1308575,3.7091823,3.2836022,2.8619268,2.920493,2.979059,3.0337205,3.0922866,3.1508527,3.4827268,3.814601,4.1464753,4.478349,4.814128,5.2201858,5.6262436,6.036206,6.4422636,6.8483214,7.211431,7.57454,7.9376497,8.300759,8.663869,9.261242,9.858616,10.455989,11.053363,11.650736,11.100216,10.549695,9.999174,9.448653,8.898132,7.918128,6.9381227,5.958118,4.9781127,3.998108,5.677001,7.355894,9.030883,10.709775,12.388668,11.350098,10.311526,9.276859,8.238289,7.1997175,7.0240197,6.844417,6.6687193,6.4891167,6.3134184,6.001066,5.688714,5.376362,5.0640097,4.7516575,5.4505453,6.1494336,6.8483214,7.551114,8.250002,6.6843367,5.114767,3.5491016,1.979532,0.41386664,2.1122816,3.8106966,5.5130157,7.211431,8.913751,7.223144,5.5364423,3.8497405,2.1630387,0.47633708,0.39044023,0.30454338,0.21864653,0.13665408,0.05075723,0.06637484,0.078088045,0.093705654,0.10932326,0.12494087,0.10932326,0.08980125,0.07418364,0.05466163,0.039044023,0.28892577,0.5388075,0.78868926,1.038571,1.2884527,1.5461433,1.8077383,2.069333,2.3270237,2.5886188,3.8302186,5.0718184,6.3134184,7.558923,8.800523,8.956698,9.116779,9.272955,9.4291315,9.589212,10.561408,11.537509,12.513609,13.4858055,14.461906,14.836729,15.207646,15.578565,15.953387,16.324306,15.543426,14.75864,13.97776,13.196879,12.412095,10.155351,7.898606,5.6418614,3.3812122,1.1244678,0.96438736,0.80430686,0.6442264,0.48414588,0.3240654,0.3240654,0.3240654,0.3240654,0.3240654,0.3240654,0.45291066,0.58175594,0.7066968,0.8355421,0.96438736,0.92534333,0.8862993,0.8511597,0.81211567,0.77307165,0.7340276,0.6910792,0.6481308,0.60518235,0.5622339,0.679366,0.79649806,0.9136301,1.0307622,1.1517987,1.2220778,1.2962615,1.3665408,1.4407244,1.5110037,1.6008049,1.6867018,1.7765031,1.8623998,1.9482968,1.8116426,1.6710842,1.5305257,1.3899672,1.2494087,1.2455044,1.2415999,1.2337911,1.2298868,1.2259823,1.0893283,0.94876975,0.81211567,0.6754616,0.5388075,0.5388075,0.5388075,0.5388075,0.5388075,0.5388075,0.47633708,0.41777104,0.359205,0.29673457,0.23816854,0.20693332,0.1717937,0.14055848,0.10932326,0.07418364,0.10151446,0.12884527,0.15617609,0.1835069,0.21083772,0.23816854,0.26940376,0.29673457,0.3240654,0.3513962,0.5192855,0.6910792,0.8589685,1.0307622,1.1986516,2.1318035,3.0649557,3.998108,4.93126,5.8644123,6.6648145,7.4691215,8.269524,9.073831,9.874233,10.124115,10.370092,10.61607,10.865952,11.111929,10.725393,10.338858,9.948417,9.561881,9.175345,9.839094,10.506746,11.170495,11.834243,12.501896,13.286681,14.07537,14.864059,15.648844,16.437534,15.808925,15.176412,14.547803,13.919194,13.286681,13.532659,13.778636,14.020708,14.2666855,14.512663,16.019762,17.526861,19.03396,20.54106,22.048159,1.3860629,1.4914817,1.5929961,1.6945106,1.796025,1.901444,1.9443923,1.9912452,2.0341935,2.0810463,2.1239948,2.182561,2.241127,2.2957885,2.3543546,2.4129205,2.4441557,2.4792955,2.5105307,2.541766,2.5769055,2.7096553,2.8463092,2.979059,3.1157131,3.2484627,3.912211,4.575959,5.2358036,5.899552,6.5633,6.547683,6.532065,6.5164475,6.5008297,6.4891167,5.4856853,4.482254,3.4788225,2.4792955,1.475864,1.3314011,1.1908426,1.0463798,0.9058213,0.76135844,0.71841,0.679366,0.63641757,0.59346914,0.5505207,0.46852827,0.38653582,0.30063897,0.21864653,0.13665408,0.10932326,0.08199245,0.05466163,0.027330816,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.046852827,0.05075723,0.058566034,0.06637484,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.05075723,0.10541886,0.15617609,0.21083772,0.26159495,0.26159495,0.25769055,0.25378615,0.25378615,0.24988174,0.22255093,0.19522011,0.1678893,0.14055848,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.8784905,1.3860629,1.8897307,2.3933985,2.900971,2.8970666,2.893162,2.893162,2.8892577,2.8892577,2.8111696,2.736986,2.6628022,2.5886188,2.514435,3.4827268,4.4510183,5.423215,6.3915067,7.363703,6.6843367,6.008875,5.3295093,4.6540475,3.9746814,3.3694992,2.7643168,2.1591344,1.5539521,0.94876975,0.92143893,0.8902037,0.8589685,0.8316377,0.80040246,0.96829176,1.1400855,1.3118792,1.4797685,1.6515622,1.6867018,1.7257458,1.7608855,1.7999294,1.8389735,1.9561055,2.077142,2.1981785,2.3192148,2.436347,3.1664703,3.8965936,4.6267166,5.35684,6.086963,5.8175592,5.548156,5.278752,5.009348,4.73604,5.1108627,5.4856853,5.8644123,6.239235,6.6140575,6.571109,6.5281606,6.4852123,6.4422636,6.3993154,6.1181984,5.833177,5.55206,5.270943,4.985922,4.919547,4.853172,4.786797,4.716518,4.650143,5.134289,5.618435,6.1064854,6.590631,7.0747766,7.4300776,7.785378,8.140678,8.495979,8.85128,9.187058,9.526741,9.86252,10.198298,10.537982,10.22563,9.913278,9.600925,9.288573,8.976221,8.554545,8.136774,7.715099,7.2934237,6.8756523,6.379793,5.883934,5.388075,4.8961205,4.4002614,5.1186714,5.840986,6.559396,7.28171,8.00012,8.628729,9.253433,9.882042,10.510651,11.139259,15.231073,19.322887,23.4147,27.506514,31.598328,35.065437,38.52864,41.99575,45.458954,48.926064,48.20375,47.481438,46.75912,46.036808,45.31059,44.67417,44.037754,43.401337,42.761013,42.124596,42.967945,43.8113,44.650745,45.494095,46.337444,38.840992,31.348446,23.851994,16.355541,8.862993,9.108971,9.358852,9.60483,9.850807,10.100689,16.378967,22.653341,28.931622,35.2099,41.48818,38.993267,36.498352,34.00344,31.508526,29.013613,39.176773,49.336025,59.499187,69.662346,79.8255,65.77356,51.72552,37.673576,23.625538,9.573594,12.376955,15.180316,17.983677,20.783133,23.586494,30.637844,37.689194,44.73664,51.78799,58.83934,51.994926,45.15441,38.309994,31.465578,24.625065,25.733915,26.84667,27.95552,29.064371,30.173222,27.018463,23.859802,20.701141,17.546383,14.387722,15.102228,15.816733,16.531239,17.245745,17.964155,15.12175,12.28325,9.440845,6.602344,3.7638438,3.8341231,3.9044023,3.970777,4.041056,4.1113358,4.8805027,5.645766,6.4149327,7.1841,7.9493628,7.746334,7.5394006,7.336372,7.1294384,6.9264097,7.3012323,7.6799593,8.058686,8.433509,8.812236,11.096312,13.376482,15.660558,17.94073,20.224804,23.426414,26.624119,29.82573,33.023434,36.225044,40.60188,44.974808,49.351646,53.724575,58.10141,55.516697,52.928078,50.34336,47.758648,45.173935,37.75557,30.34111,22.922745,15.504381,8.086017,7.016211,5.9464045,4.8765984,3.8067923,2.736986,2.9478238,3.1586614,3.3655949,3.5764325,3.78727,3.0727646,2.358259,1.6437533,0.92924774,0.21083772,1.0619974,1.9092526,2.7565079,3.6037633,4.4510183,4.3455997,4.240181,4.134762,4.029343,3.9239242,6.387602,8.85128,11.311053,13.774731,16.238409,16.484386,16.734268,16.980246,17.226223,17.476105,15.879204,14.286208,12.689307,11.096312,9.499411,8.238289,6.9810715,5.7199492,4.4588275,3.2016098,2.8970666,2.5964274,2.2918842,1.9912452,1.6867018,2.6940374,3.697469,4.7009,5.708236,6.7116675,6.098676,5.481781,4.8687897,4.251894,3.638903,6.141625,8.648251,11.150972,13.657599,16.164225,14.930434,13.696643,12.466757,11.232965,9.999174,9.202676,8.406178,7.605776,6.8092775,6.012779,5.700427,5.388075,5.0757227,4.7633705,4.4510183,4.1035266,3.7599394,3.416352,3.06886,2.7252727,2.8658314,3.0063896,3.1469483,3.2836022,3.4241607,3.7638438,4.1035266,4.4432096,4.786797,5.12648,5.45445,5.7785153,6.1064854,6.434455,6.7624245,7.0240197,7.2856145,7.551114,7.812709,8.074304,9.081639,10.088976,11.096312,12.103647,13.110983,12.224684,11.338385,10.44818,9.561881,8.675582,7.7892823,6.9068875,6.0205884,5.134289,4.251894,5.3295093,6.4110284,7.4886436,8.570163,9.651682,9.136301,8.624825,8.113348,7.601871,7.08649,7.0591593,7.027924,6.996689,6.969358,6.9381227,6.426646,5.911265,5.3997884,4.8883114,4.376835,4.73604,5.099149,5.462259,5.825368,6.1884775,5.0757227,3.9668727,2.8580225,1.7491722,0.63641757,2.3114061,3.9863946,5.661383,7.336372,9.01136,7.387129,5.7628975,4.138666,2.5105307,0.8862993,0.71841,0.5466163,0.37872702,0.20693332,0.039044023,0.05466163,0.07418364,0.08980125,0.10932326,0.12494087,0.113227665,0.10541886,0.093705654,0.08589685,0.07418364,0.27330816,0.47633708,0.6754616,0.8745861,1.0737107,1.6827974,2.2918842,2.8970666,3.506153,4.1113358,5.2358036,6.356367,7.480835,8.601398,9.725866,9.866425,10.003078,10.143637,10.284196,10.424754,11.0494585,11.674163,12.298867,12.923572,13.548276,13.919194,14.2901125,14.661031,15.031949,15.398962,14.360392,13.32182,12.2793455,11.240774,10.198298,8.433509,6.6687193,4.903929,3.1391394,1.3743496,1.2181735,1.0580931,0.9019169,0.74574083,0.58566034,0.57394713,0.5622339,0.5505207,0.5388075,0.5231899,0.59346914,0.659844,0.7262188,0.79649806,0.8628729,0.8238289,0.78868926,0.74964523,0.7106012,0.6754616,0.6910792,0.7066968,0.71841,0.7340276,0.74964523,0.8980125,1.0463798,1.1908426,1.33921,1.4875772,1.5188124,1.5539521,1.5851873,1.6164225,1.6515622,1.6749885,1.698415,1.7257458,1.7491722,1.7765031,1.620327,1.4641509,1.3118792,1.1557031,0.999527,0.9917182,0.98000497,0.96829176,0.96048295,0.94876975,0.8511597,0.74964523,0.6481308,0.5505207,0.44900626,0.44900626,0.44900626,0.44900626,0.44900626,0.44900626,0.40605783,0.359205,0.31625658,0.26940376,0.22645533,0.19912452,0.1717937,0.14055848,0.113227665,0.08589685,0.10541886,0.12103647,0.14055848,0.15617609,0.1756981,0.19131571,0.21083772,0.22645533,0.24597734,0.26159495,0.39044023,0.5192855,0.6442264,0.77307165,0.9019169,1.6008049,2.3035975,3.0063896,3.7091823,4.4119744,5.02887,5.645766,6.266566,6.883461,7.5003567,7.8088045,8.113348,8.421796,8.730244,9.0386915,9.288573,9.538455,9.788337,10.0382185,10.2881,10.928422,11.572648,12.216875,12.857197,13.501423,14.223738,14.949956,15.676175,16.398489,17.124708,16.214983,15.305257,14.395531,13.4858055,12.576079,12.615124,12.654168,12.693212,12.73616,12.775204,14.126127,15.480955,16.831879,18.186707,19.537628,1.4251068,1.5227169,1.620327,1.717937,1.815547,1.9131571,1.9561055,1.999054,2.0380979,2.0810463,2.1239948,2.194274,2.260649,2.3270237,2.3933985,2.463678,2.4910088,2.522244,2.5534792,2.5808098,2.612045,2.7408905,2.8658314,2.9946766,3.1235218,3.2484627,3.873167,4.5017757,5.12648,5.7511845,6.375889,6.329036,6.278279,6.2314262,6.184573,6.13772,5.263134,4.3924527,3.521771,2.6471848,1.7765031,1.6281357,1.4836729,1.33921,1.1947471,1.0502841,0.92924774,0.80821127,0.6910792,0.5700427,0.44900626,0.38263142,0.31625658,0.24597734,0.1796025,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.031235218,0.03513962,0.039044023,0.046852827,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.1756981,0.1796025,0.1835069,0.1835069,0.18741131,0.1639849,0.14055848,0.12103647,0.09761006,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,1.1557031,1.8780174,2.5964274,3.3187418,4.037152,4.0020123,3.9668727,3.9317331,3.8965936,3.8614538,3.5998588,3.338264,3.076669,2.8111696,2.5495746,3.3421683,4.134762,4.927356,5.7199492,6.5125427,6.126007,5.743376,5.35684,4.9742084,4.5876727,3.9551594,3.3226464,2.690133,2.05762,1.4251068,1.3782539,1.3353056,1.2884527,1.2455044,1.1986516,1.456342,1.7101282,1.9639144,2.2216048,2.475391,2.2255092,1.9756275,1.7257458,1.475864,1.2259823,1.5539521,1.8858263,2.2137961,2.5456703,2.87364,3.4827268,4.0918136,4.6969957,5.3060827,5.911265,5.743376,5.579391,5.4115014,5.2436123,5.0757227,5.388075,5.700427,6.012779,6.3251314,6.6374836,6.6687193,6.6960497,6.727285,6.75852,6.785851,6.3836975,5.9776397,5.571582,5.169429,4.7633705,4.6423345,4.521298,4.4041657,4.283129,4.1620927,4.7009,5.2436123,5.7824197,6.321227,6.8639393,7.230953,7.601871,7.9727893,8.343708,8.710721,9.050405,9.386183,9.725866,10.061645,10.401327,10.100689,9.80005,9.499411,9.198771,8.898132,8.734148,8.566258,8.398369,8.23048,8.062591,7.5823493,7.1021075,6.621866,6.141625,5.661383,6.1299114,6.5984397,7.066968,7.531592,8.00012,8.55845,9.120684,9.679013,10.241247,10.799577,15.008522,19.213564,23.422508,27.631454,31.836496,36.510067,41.183636,45.853302,50.52687,55.20044,54.02131,52.846085,51.666954,50.49173,49.3126,47.438488,45.564373,43.686356,41.812244,39.93813,40.769768,41.601406,42.436947,43.268585,44.100224,37.095726,30.091228,23.086731,16.07833,9.073831,9.17925,9.280765,9.382278,9.483793,9.589212,15.758167,21.931028,28.103888,34.27675,40.449608,38.231907,36.014206,33.796505,31.578806,29.361105,37.060585,44.763973,52.46345,60.162933,67.86242,56.250725,44.63903,33.023434,21.411741,9.80005,12.849388,15.894821,18.94416,21.989594,25.03893,30.325493,35.612053,40.898613,46.18908,51.47564,45.806446,40.13335,34.464157,28.794966,23.125774,26.089216,29.056562,32.020004,34.983444,37.95079,33.519295,29.091702,24.660204,20.228708,15.801116,17.120804,18.444397,19.767988,21.091581,22.411268,18.690374,14.969479,11.2446785,7.523783,3.7989833,3.8302186,3.8614538,3.8887846,3.9200199,3.951255,4.607195,5.263134,5.9229784,6.578918,7.238762,6.942027,6.649197,6.3524623,6.055728,5.7628975,6.6726236,7.5823493,8.492075,9.4018,10.311526,10.967466,11.623405,12.2793455,12.93138,13.58732,18.32336,23.063305,27.799343,32.539288,37.27533,39.348564,41.42571,43.498947,45.576088,47.649326,44.822536,41.99575,39.168964,36.338272,33.511486,28.791061,24.07064,19.354122,14.633699,9.913278,8.320281,6.727285,5.134289,3.541293,1.9482968,2.5769055,3.2055142,3.8341231,4.4588275,5.087436,4.126953,3.1664703,2.2059872,1.2494087,0.28892577,1.3782539,2.4675822,3.5569105,4.646239,5.735567,5.630148,5.520825,5.4154058,5.3060827,5.2006636,7.437886,9.675109,11.912332,14.149553,16.386776,15.7035055,15.016331,14.33306,13.645885,12.962616,11.681972,10.401327,9.120684,7.843944,6.5633,5.9346914,5.3060827,4.6813784,4.0527697,3.4241607,2.9634414,2.5066261,2.0459068,1.5851873,1.1244678,2.2840753,3.4397783,4.5993857,5.755089,6.910792,6.250948,5.591104,4.93126,4.271416,3.611572,6.657006,9.702439,12.747873,15.793307,18.838741,17.070047,15.3013525,13.536563,11.767868,9.999174,9.183154,8.371038,7.5550184,6.7389984,5.9268827,5.5247293,5.12648,4.7243266,4.3260775,3.9239242,3.6584249,3.3890212,3.1235218,2.854118,2.5886188,2.8111696,3.0337205,3.2562714,3.4788225,3.7013733,4.0488653,4.396357,4.743849,5.0913405,5.4388323,5.6848097,5.930787,6.180669,6.426646,6.676528,6.8366084,7.000593,7.1606736,7.3246584,7.4886436,8.905942,10.323239,11.740538,13.157836,14.575133,13.349152,12.123169,10.901091,9.675109,8.449126,7.660437,6.871748,6.0791545,5.290465,4.5017757,4.9820175,5.466163,5.9464045,6.4305506,6.910792,6.9264097,6.9381227,6.949836,6.9615493,6.9732623,7.094299,7.211431,7.328563,7.445695,7.562827,6.8483214,6.13772,5.423215,4.7126136,3.998108,4.025439,4.0488653,4.0761957,4.0996222,4.123049,3.4710135,2.8189783,2.1669433,1.5149081,0.8628729,2.514435,4.1620927,5.813655,7.461313,9.112875,7.551114,5.989353,4.423688,2.8619268,1.3001659,1.0463798,0.78868926,0.5349031,0.28111696,0.023426414,0.046852827,0.06637484,0.08589685,0.10541886,0.12494087,0.12103647,0.12103647,0.11713207,0.113227665,0.113227665,0.26159495,0.41386664,0.5622339,0.7106012,0.8628729,1.8194515,2.7721257,3.7287042,4.6813784,5.6379566,6.6413884,7.6409154,8.644346,9.647778,10.651209,10.772245,10.893282,11.018223,11.139259,11.2642,11.537509,11.810817,12.08803,12.361338,12.63855,13.005564,13.372578,13.739592,14.106606,14.473619,13.177358,11.881096,10.58093,9.284669,7.988407,6.715572,5.4427366,4.169902,2.8970666,1.6242313,1.4680552,1.3157835,1.1596074,1.0034313,0.8511597,0.8238289,0.80040246,0.77307165,0.74964523,0.7262188,0.7340276,0.7418364,0.74574083,0.75354964,0.76135844,0.7262188,0.6871748,0.6481308,0.61299115,0.57394713,0.6481308,0.71841,0.79259366,0.8667773,0.93705654,1.116659,1.2923572,1.4719596,1.6476578,1.8233559,1.8194515,1.8116426,1.8038338,1.796025,1.7882162,1.7491722,1.7140326,1.6749885,1.6359446,1.6008049,1.4290112,1.261122,1.0893283,0.92143893,0.74964523,0.7340276,0.71841,0.7066968,0.6910792,0.6754616,0.61299115,0.5505207,0.48805028,0.42557985,0.3631094,0.3631094,0.3631094,0.3631094,0.3631094,0.3631094,0.3318742,0.30063897,0.27330816,0.24207294,0.21083772,0.19131571,0.1678893,0.14446288,0.12103647,0.10151446,0.10932326,0.113227665,0.12103647,0.12884527,0.13665408,0.14446288,0.15227169,0.16008049,0.1678893,0.1756981,0.26159495,0.3435874,0.42948425,0.5153811,0.60127795,1.0737107,1.5461433,2.018576,2.4910088,2.9634414,3.39683,3.8263142,4.2597027,4.6930914,5.12648,5.493494,5.860508,6.2275214,6.5945354,6.9615493,7.8517528,8.738052,9.6243515,10.510651,11.400854,12.021654,12.63855,13.25935,13.88015,14.50095,15.160794,15.824542,16.48829,17.148134,17.811884,16.62104,15.434102,14.243259,13.052417,11.861574,11.697589,11.533605,11.365715,11.20173,11.037745,12.236397,13.431144,14.629795,15.828446,17.023193,1.4641509,1.5539521,1.6476578,1.7413634,1.8311646,1.9248703,1.9639144,2.0068626,2.0459068,2.084951,2.1239948,2.2020829,2.280171,2.358259,2.436347,2.514435,2.541766,2.5690966,2.5964274,2.6237583,2.6510892,2.7682211,2.8892577,3.0102942,3.1313305,3.2484627,3.8380275,4.423688,5.0132523,5.5989127,6.1884775,6.1064854,6.028397,5.9464045,5.8683167,5.786324,5.044488,4.3026514,3.5608149,2.8189783,2.0732377,1.9287747,1.7804074,1.6320401,1.4836729,1.33921,1.1400855,0.94096094,0.74574083,0.5466163,0.3513962,0.29673457,0.24597734,0.19131571,0.14055848,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.015617609,0.015617609,0.019522011,0.023426414,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.093705654,0.10151446,0.10932326,0.11713207,0.12494087,0.10932326,0.08980125,0.07418364,0.05466163,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,1.43682,2.3699722,3.3031244,4.240181,5.173333,5.1069584,5.040583,4.9742084,4.903929,4.8375545,4.388548,3.9356375,3.4866312,3.0376248,2.5886188,3.2016098,3.8185053,4.4314966,5.0483923,5.661383,5.571582,5.477876,5.3841705,5.2943697,5.2006636,4.5408196,3.8809757,3.2211318,2.5612879,1.901444,1.8389735,1.7804074,1.7218413,1.6593709,1.6008049,1.9404879,2.280171,2.619854,2.959537,3.2992198,2.7643168,2.2255092,1.6867018,1.1517987,0.61299115,1.1517987,1.6906061,2.233318,2.7721257,3.310933,3.7989833,4.283129,4.7672753,5.251421,5.735567,5.6730967,5.606722,5.5442514,5.477876,5.4115014,5.661383,5.911265,6.1611466,6.4110284,6.66091,6.7663293,6.8678436,6.969358,7.0708723,7.1762915,6.649197,6.1181984,5.591104,5.0640097,4.5369153,4.365122,4.193328,4.0215344,3.8458362,3.6740425,4.271416,4.8648853,5.4583545,6.055728,6.649197,7.0357327,7.4183645,7.8049,8.191436,8.574067,8.913751,9.249529,9.589212,9.924991,10.260769,9.975748,9.686822,9.4018,9.112875,8.823949,8.909846,8.995743,9.081639,9.163632,9.249529,8.784905,8.320281,7.8556576,7.3910336,6.9264097,7.141152,7.355894,7.570636,7.785378,8.00012,8.492075,8.98403,9.475985,9.971844,10.4637985,14.785972,19.108145,23.430319,27.752491,32.074665,37.954693,43.834724,49.714752,55.594784,61.474815,59.842773,58.21073,56.578693,54.94665,53.310707,50.1989,47.08709,43.97528,40.863476,37.751667,38.57159,39.39542,40.219246,41.039173,41.863003,35.346554,28.834011,22.317564,15.801116,9.288573,9.245625,9.202676,9.159728,9.116779,9.073831,15.141272,21.208714,27.276154,33.343594,39.411037,37.474453,35.533966,33.593475,31.652988,29.712502,34.948303,40.18801,45.423817,50.663525,55.899326,46.72398,37.548637,28.373291,19.197947,10.0265045,13.317916,16.609327,19.900738,23.196054,26.487465,30.01314,33.538815,37.06449,40.58626,44.11194,39.614067,35.116196,30.618322,26.124355,21.626484,26.444517,31.266453,36.084484,40.90642,45.724453,40.02403,34.319695,28.615364,22.914936,17.210606,19.143284,21.07206,23.000834,24.933514,26.862288,22.258997,17.651802,13.048512,8.441318,3.8380275,3.8263142,3.8185053,3.8067923,3.7989833,3.78727,4.3338866,4.884407,5.4310236,5.9776397,6.524256,6.141625,5.755089,5.368553,4.985922,4.5993857,6.044015,7.4847393,8.929368,10.370092,11.810817,10.838621,9.866425,8.894228,7.9220324,6.949836,13.224211,19.498585,25.776863,32.05124,38.32561,38.099155,37.876606,37.65015,37.423695,37.201145,34.12838,31.05952,27.99066,24.921799,21.849035,19.826555,17.804073,15.781594,13.759113,11.736633,9.620447,7.5081654,5.3919797,3.2757936,1.1635119,2.2059872,3.252367,4.298747,5.3412223,6.387602,5.181142,3.978586,2.7721257,1.5656652,0.3631094,1.6945106,3.0259118,4.3612175,5.6926184,7.0240197,6.914696,6.805373,6.6960497,6.5867267,6.473499,8.488171,10.498938,12.513609,14.524376,16.539047,14.918721,13.302299,11.685876,10.065549,8.449126,7.4847393,6.520352,5.5559645,4.591577,3.6232853,3.631094,3.6349986,3.638903,3.6467118,3.6506162,3.0337205,2.416825,1.796025,1.1791295,0.5622339,1.8741131,3.182088,4.493967,5.801942,7.113821,6.407124,5.704332,4.997635,4.290938,3.5881457,7.172387,10.756628,14.34087,17.929016,21.513256,19.20966,16.906061,14.606369,12.302772,9.999174,9.167537,8.335898,7.504261,6.6687193,5.8370814,5.349031,4.860981,4.376835,3.8887846,3.4007344,3.2094188,3.018103,2.8306916,2.639376,2.4480603,2.7565079,3.0610514,3.3655949,3.6701381,3.9746814,4.3299823,4.6852827,5.040583,5.395884,5.7511845,5.919074,6.083059,6.250948,6.4188375,6.5867267,6.649197,6.7116675,6.774138,6.8366084,6.899079,8.726339,10.553599,12.380859,14.208119,16.039284,14.473619,12.911859,11.350098,9.788337,8.226576,7.531592,6.8366084,6.141625,5.446641,4.7516575,4.6345253,4.521298,4.4041657,4.290938,4.173806,4.7126136,5.251421,5.786324,6.3251314,6.8639393,7.1294384,7.3910336,7.656533,7.9220324,8.187531,7.2739015,6.364176,5.4505453,4.5369153,3.6232853,3.310933,2.998581,2.6862288,2.3738766,2.0615244,1.8663043,1.6710842,1.475864,1.2806439,1.0893283,2.7135596,4.337791,5.9620223,7.5862536,9.21439,7.7111945,6.211904,4.7126136,3.213323,1.7140326,1.3743496,1.0307622,0.6910792,0.3513962,0.011713207,0.03513962,0.058566034,0.078088045,0.10151446,0.12494087,0.12884527,0.13665408,0.14055848,0.14446288,0.14836729,0.24988174,0.3513962,0.44900626,0.5505207,0.6481308,1.9522011,3.2562714,4.5564375,5.860508,7.1606736,8.046973,8.929368,9.811763,10.694158,11.576552,11.678067,11.783486,11.888905,11.994324,12.099743,12.025558,11.951375,11.873287,11.799104,11.72492,12.091934,12.455043,12.818152,13.185166,13.548276,11.994324,10.4403715,8.886419,7.328563,5.774611,4.9937305,4.2167544,3.435874,2.6549935,1.8741131,1.7218413,1.5695697,1.4172981,1.2650263,1.1127546,1.0737107,1.038571,0.999527,0.96438736,0.92534333,0.8706817,0.8199245,0.76916724,0.7145056,0.6637484,0.62470436,0.58566034,0.5505207,0.5114767,0.47633708,0.60518235,0.7340276,0.8667773,0.9956226,1.1244678,1.3314011,1.5383345,1.7491722,1.9561055,2.1630387,2.1161861,2.069333,2.018576,1.9717231,1.9248703,1.8233559,1.7257458,1.6242313,1.5266213,1.4251068,1.2415999,1.0541886,0.8706817,0.6832704,0.4997635,0.48024148,0.46071947,0.44119745,0.42167544,0.39824903,0.37482262,0.3513962,0.3240654,0.30063897,0.27330816,0.27330816,0.27330816,0.27330816,0.27330816,0.27330816,0.26159495,0.24597734,0.23035973,0.21474212,0.19912452,0.1835069,0.1639849,0.14836729,0.12884527,0.113227665,0.10932326,0.10932326,0.10541886,0.10151446,0.10151446,0.09761006,0.093705654,0.093705654,0.08980125,0.08589685,0.12884527,0.1717937,0.21474212,0.25769055,0.30063897,0.5427119,0.78478485,1.0268579,1.2689307,1.5110037,1.7608855,2.0068626,2.2567444,2.5027218,2.7486992,3.1781836,3.6037633,4.0332475,4.4588275,4.8883114,6.4110284,7.9376497,9.464272,10.986988,12.513609,13.110983,13.708356,14.30573,14.903104,15.500477,16.101755,16.69913,17.300406,17.901684,18.499058,17.031002,15.559043,14.090988,12.619028,11.150972,10.780055,10.409137,10.0382185,9.671205,9.300286,10.342762,11.385237,12.427712,13.470188,14.512663,1.4992905,1.5890918,1.6749885,1.7608855,1.8506867,1.9365835,1.9756275,2.0107672,2.0498111,2.0888553,2.1239948,2.2137961,2.2996929,2.3855898,2.475391,2.5612879,2.5886188,2.612045,2.639376,2.6628022,2.6862288,2.7994564,2.912684,3.0259118,3.1391394,3.2484627,3.7989833,4.349504,4.900025,5.4505453,6.001066,5.8878384,5.774611,5.661383,5.548156,5.4388323,4.825841,4.21285,3.5998588,2.9868677,2.3738766,2.2255092,2.0732377,1.9248703,1.7765031,1.6242313,1.3509232,1.0737107,0.80040246,0.5231899,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.113227665,0.22645533,0.3357786,0.44900626,0.5622339,1.7140326,2.8619268,4.0137253,5.1616197,6.3134184,6.211904,6.114294,6.012779,5.911265,5.813655,5.173333,4.5369153,3.900498,3.2640803,2.6237583,3.0610514,3.4983444,3.9356375,4.376835,4.814128,5.0132523,5.212377,5.4115014,5.610626,5.813655,5.12648,4.4393053,3.7482262,3.0610514,2.3738766,2.2996929,2.2255092,2.1513257,2.0732377,1.999054,2.4246337,2.8502135,3.2757936,3.7013733,4.123049,3.2992198,2.475391,1.6515622,0.8238289,0.0,0.74964523,1.4992905,2.2489357,2.998581,3.7482262,4.1113358,4.474445,4.8375545,5.2006636,5.563773,5.5989127,5.6379566,5.6730967,5.7121406,5.7511845,5.938596,6.126007,6.3134184,6.5008297,6.688241,6.8639393,7.0357327,7.211431,7.387129,7.562827,6.910792,6.262661,5.610626,4.9624953,4.3143644,4.087909,3.8614538,3.638903,3.4124475,3.1859922,3.8380275,4.4861584,5.138193,5.786324,6.4383593,6.8366084,7.238762,7.6370106,8.039165,8.437413,8.773191,9.112875,9.448653,9.788337,10.124115,9.850807,9.573594,9.300286,9.023073,8.749765,9.085544,9.425227,9.761005,10.100689,10.436467,9.987461,9.538455,9.085544,8.636538,8.187531,8.148487,8.113348,8.074304,8.039165,8.00012,8.4257,8.85128,9.276859,9.698535,10.124115,14.56342,18.998821,23.438128,27.873528,32.31283,39.399323,46.485813,53.576206,60.662697,67.74919,65.66424,63.575382,61.486526,59.401577,57.31272,52.963215,48.613712,44.26421,39.9108,35.561295,36.373413,37.185528,38.00155,38.813663,39.62578,33.601284,27.576794,21.548395,15.523903,9.499411,9.311999,9.124588,8.937177,8.749765,8.562354,14.524376,20.486399,26.448421,32.41435,38.37637,36.713093,35.04982,33.386543,31.723269,30.063898,32.83602,35.612053,38.388084,41.164112,43.936237,37.201145,30.462147,23.723148,16.988054,10.249056,13.786445,17.323833,20.861221,24.39861,27.935999,29.700788,31.461674,33.226463,34.98735,36.748234,33.425587,30.099037,26.77639,23.44984,20.12329,26.799816,33.476345,40.148968,46.825497,53.49812,46.524857,39.551594,32.57443,25.601166,18.623999,21.16186,23.699722,26.237583,28.775444,31.313307,25.823717,20.338032,14.848442,9.362757,3.873167,3.8263142,3.775557,3.7247996,3.6740425,3.6232853,4.0605783,4.5017757,4.939069,5.376362,5.813655,5.337318,4.860981,4.388548,3.912211,3.435874,5.4115014,7.387129,9.362757,11.338385,13.314012,10.71368,8.113348,5.5130157,2.912684,0.31235218,8.125061,15.93777,23.750479,31.563189,39.375896,36.849747,34.3236,31.801357,29.275208,26.74906,23.438128,20.12329,16.812357,13.501423,10.186585,10.862047,11.537509,12.212971,12.888432,13.563893,10.924518,8.289046,5.64967,3.0141985,0.37482262,1.8389735,3.2992198,4.7633705,6.223617,7.687768,6.239235,4.786797,3.338264,1.8858263,0.43729305,2.0107672,3.5881457,5.1616197,6.7389984,8.312472,8.1992445,8.086017,7.9766936,7.8634663,7.7502384,9.538455,11.326671,13.110983,14.899199,16.687416,14.13784,11.588266,9.0386915,6.4891167,3.9356375,3.2875066,2.639376,1.9873407,1.33921,0.6871748,1.3235924,1.9639144,2.6003318,3.2367494,3.873167,3.1000953,2.3231194,1.5500476,0.77307165,0.0,1.4641509,2.9243972,4.388548,5.8487945,7.3129454,6.5633,5.813655,5.0640097,4.3143644,3.5608149,7.687768,11.810817,15.93777,20.06082,24.187773,21.349272,18.51077,15.676175,12.837675,9.999174,9.148014,8.300759,7.4495993,6.5984397,5.7511845,5.173333,4.5993857,4.025439,3.4514916,2.87364,2.7643168,2.6510892,2.5378613,2.4246337,2.3114061,2.7018464,3.0883822,3.474918,3.8614538,4.251894,4.6110992,4.9742084,5.337318,5.700427,6.0635366,6.1494336,6.239235,6.3251314,6.4110284,6.5008297,6.461786,6.426646,6.387602,6.348558,6.3134184,8.550641,10.787864,13.025085,15.262308,17.49953,15.598087,13.700547,11.799104,9.901564,8.00012,7.3988423,6.801469,6.2001905,5.5989127,5.001539,4.2870336,3.5764325,2.8619268,2.1513257,1.43682,2.4988174,3.5608149,4.6267166,5.688714,6.7507114,7.1606736,7.57454,7.988407,8.398369,8.812236,7.699481,6.5867267,5.473972,4.3612175,3.2484627,2.6003318,1.9482968,1.3001659,0.6481308,0.0,0.26159495,0.5231899,0.78868926,1.0502841,1.3118792,2.912684,4.513489,6.114294,7.7111945,9.311999,7.8751793,6.4383593,5.001539,3.5608149,2.1239948,1.698415,1.2767396,0.8511597,0.42557985,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.23816854,0.28892577,0.3357786,0.38653582,0.43729305,2.0888553,3.736513,5.388075,7.0357327,8.687295,9.448653,10.213917,10.975275,11.736633,12.501896,12.587793,12.67369,12.763491,12.849388,12.939189,12.513609,12.08803,11.66245,11.23687,10.81129,11.174399,11.537509,11.900618,12.263727,12.626837,10.81129,8.999647,7.1880045,5.376362,3.5608149,3.2757936,2.9868677,2.7018464,2.4129205,2.1239948,1.9756275,1.8233559,1.6749885,1.5266213,1.3743496,1.3235924,1.2767396,1.2259823,1.175225,1.1244678,1.0112402,0.9019169,0.78868926,0.6754616,0.5622339,0.5231899,0.48805028,0.44900626,0.41386664,0.37482262,0.5622339,0.74964523,0.93705654,1.1244678,1.3118792,1.5500476,1.7882162,2.0263848,2.260649,2.4988174,2.4129205,2.3231194,2.2372224,2.1513257,2.0615244,1.901444,1.737459,1.5734742,1.4133936,1.2494087,1.0502841,0.8511597,0.6481308,0.44900626,0.24988174,0.22645533,0.19912452,0.1756981,0.14836729,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.37482262,0.8628729,1.3509232,1.8389735,2.3231194,2.8111696,4.9742084,7.137247,9.300286,11.4633255,13.626364,14.200311,14.774258,15.348206,15.926057,16.500004,17.03881,17.573715,18.112522,18.651329,19.186234,17.437061,15.687888,13.938716,12.189544,10.436467,9.86252,9.288573,8.710721,8.136774,7.562827,8.449126,9.339331,10.22563,11.111929,11.998228,1.5110037,1.5969005,1.678893,1.7608855,1.8428779,1.9248703,1.9639144,1.999054,2.0380979,2.0732377,2.1122816,2.1981785,2.2840753,2.366068,2.4519646,2.5378613,2.5769055,2.6159496,2.6588979,2.697942,2.736986,2.87364,3.0141985,3.1508527,3.2875066,3.4241607,3.9083066,4.388548,4.872694,5.35684,5.8370814,5.9815445,6.1221027,6.266566,6.407124,6.551587,5.6535745,4.755562,3.8575494,2.959537,2.0615244,1.9131571,1.7608855,1.6125181,1.4641509,1.3118792,1.1010414,0.8862993,0.6754616,0.46071947,0.24988174,0.21474212,0.1796025,0.14446288,0.10932326,0.07418364,0.07027924,0.06637484,0.058566034,0.05466163,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.046852827,0.039044023,0.03513962,0.031235218,0.023426414,0.023426414,0.019522011,0.015617609,0.015617609,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.12884527,0.11713207,0.10932326,0.09761006,0.08589685,0.12494087,0.1639849,0.19912452,0.23816854,0.27330816,0.6481308,1.0268579,1.4016805,1.7765031,2.1513257,3.0883822,4.025439,4.9624953,5.899552,6.8366084,6.6335793,6.434455,6.2314262,6.028397,5.825368,5.270943,4.716518,4.1581883,3.6037633,3.049338,3.3031244,3.5569105,3.8067923,4.0605783,4.3143644,4.7399445,5.169429,5.5950084,6.0205884,6.4500723,5.8683167,5.2865605,4.7009,4.1191444,3.5373883,3.4788225,3.4241607,3.3655949,3.3070288,3.2484627,3.3421683,3.435874,3.5256753,3.619381,3.7130866,2.97125,2.2294137,1.4836729,0.7418364,0.0,0.60518235,1.2103647,1.815547,2.4207294,3.0259118,3.59205,4.1581883,4.728231,5.2943697,5.8644123,5.813655,5.7628975,5.7121406,5.661383,5.610626,5.7668023,5.9229784,6.0791545,6.2314262,6.387602,6.5984397,6.8092775,7.016211,7.2270484,7.437886,6.8483214,6.2587566,5.6691923,5.0757227,4.4861584,4.447114,4.40807,4.369026,4.3260775,4.2870336,4.7516575,5.212377,5.6730967,6.13772,6.5984397,7.0474463,7.4964523,7.941554,8.39056,8.835662,9.124588,9.413514,9.698535,9.987461,10.276386,10.073358,9.870329,9.6673,9.464272,9.261242,9.534551,9.807858,10.081166,10.350571,10.6238785,10.4286585,10.229534,10.034314,9.835189,9.636065,9.651682,9.6673,9.682918,9.698535,9.714153,9.983557,10.256865,10.530173,10.803481,11.076789,15.285735,19.49468,23.703627,27.916475,32.125423,40.01622,47.91092,55.801716,63.69642,71.58721,70.02155,68.45589,66.89413,65.32846,63.762794,58.808105,53.85342,48.898735,43.944046,38.98936,38.32171,37.654057,36.986404,36.31875,35.651096,30.204456,24.761719,19.315079,13.868437,8.4257,8.359325,8.296855,8.23048,8.164105,8.101635,13.224211,18.346786,23.469362,28.591938,33.71061,33.253796,32.793076,32.332355,31.871635,31.410915,33.253796,35.096672,36.93955,38.78243,40.625305,34.725754,28.830107,22.930555,17.034906,11.139259,14.309634,17.483913,20.654287,23.828568,26.998941,28.357674,29.716406,31.071234,32.429966,33.788696,31.086851,28.388908,25.687063,22.98912,20.287273,26.61631,32.94925,39.278286,45.607323,51.93636,45.138794,38.34123,31.543665,24.746101,17.948538,20.423927,22.895414,25.366901,27.838388,30.31378,25.14435,19.978827,14.809398,9.643873,4.474445,4.853172,5.2358036,5.6145306,5.9932575,6.375889,6.832704,7.289519,7.746334,8.203149,8.663869,7.8205175,6.9810715,6.141625,5.3021784,4.462732,5.801942,7.141152,8.484266,9.823476,11.162686,9.245625,7.3324676,5.4193106,3.5022488,1.5890918,8.382751,15.176412,21.973976,28.767635,35.561295,33.171803,30.782307,28.392813,26.003319,23.613825,21.22433,18.838741,16.449247,14.063657,11.674163,11.650736,11.623405,11.599979,11.576552,11.549222,9.300286,7.0513506,4.7985106,2.5495746,0.30063897,2.0146716,3.7287042,5.446641,7.1606736,8.874706,8.449126,8.023546,7.601871,7.1762915,6.7507114,8.078208,9.405705,10.733202,12.0606985,13.388195,13.16174,12.93138,12.704925,12.47847,12.24811,12.86891,13.4858055,14.102701,14.719597,15.336493,12.900145,10.4637985,8.023546,5.5871997,3.1508527,3.3812122,3.6154766,3.8458362,4.0801005,4.3143644,5.1225758,5.930787,6.7429028,7.551114,8.36323,7.785378,7.2075267,6.629675,6.0518236,5.473972,5.688714,5.899552,6.114294,6.3251314,6.5359693,5.919074,5.298274,4.677474,4.056674,3.435874,7.6838636,11.927949,16.172033,20.416119,24.664108,21.439074,18.217941,14.996809,11.771772,8.550641,8.011833,7.4691215,6.930314,6.3915067,5.8487945,5.185046,4.521298,3.853645,3.1898966,2.5261483,2.6042364,2.67842,2.7565079,2.8345962,2.912684,3.3187418,3.7208953,4.126953,4.533011,4.939069,5.270943,5.602817,5.9346914,6.266566,6.5984397,6.524256,6.446168,6.36808,6.289992,6.211904,6.2938967,6.3719845,6.453977,6.532065,6.6140575,8.98403,11.354002,13.723974,16.093946,18.463919,16.570284,14.676648,12.783013,10.893282,8.999647,8.214863,7.4300776,6.6452928,5.860508,5.0757227,4.5564375,4.0332475,3.513962,2.9946766,2.475391,3.2718892,4.0644827,4.860981,5.6535745,6.4500723,6.6960497,6.9459314,7.191909,7.4417906,7.687768,6.8209906,5.9542136,5.083532,4.2167544,3.349977,2.6940374,2.0341935,1.3782539,0.71841,0.062470436,0.41386664,0.76916724,1.1205635,1.4719596,1.8233559,3.2640803,4.7009,6.13772,7.57454,9.01136,7.6838636,6.356367,5.02887,3.7013733,2.3738766,1.901444,1.4251068,0.94876975,0.47633708,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.14836729,0.19522011,0.24207294,0.28892577,0.3357786,0.63251317,0.92924774,1.2220778,1.5188124,1.8116426,2.8892577,3.9668727,5.044488,6.1221027,7.1997175,8.117252,9.034787,9.952321,10.869856,11.787391,11.533605,11.275913,11.022127,10.768341,10.510651,10.178777,9.8429985,9.507219,9.171441,8.835662,9.136301,9.43694,9.737579,10.0382185,10.338858,8.85128,7.363703,5.8761253,4.388548,2.900971,2.6628022,2.4246337,2.1864653,1.9482968,1.7140326,1.5929961,1.4719596,1.3509232,1.2337911,1.1127546,1.1010414,1.0932326,1.0815194,1.0737107,1.0619974,0.96048295,0.8589685,0.75354964,0.6520352,0.5505207,0.5388075,0.5231899,0.5114767,0.4997635,0.48805028,0.62860876,0.77307165,0.9136301,1.0580931,1.1986516,1.3743496,1.5500476,1.7257458,1.901444,2.0732377,1.9951496,1.9131571,1.8350691,1.7530766,1.6749885,1.5461433,1.4212024,1.2923572,1.1635119,1.038571,0.8823949,0.7262188,0.57394713,0.41777104,0.26159495,0.24597734,0.22645533,0.21083772,0.19131571,0.1756981,0.1835069,0.19522011,0.20693332,0.21474212,0.22645533,0.21864653,0.21083772,0.20302892,0.19522011,0.18741131,0.19912452,0.20693332,0.21864653,0.22645533,0.23816854,0.24988174,0.26159495,0.27330816,0.28892577,0.30063897,0.3357786,0.37482262,0.41386664,0.44900626,0.48805028,0.5114767,0.5388075,0.5622339,0.58566034,0.61299115,0.5583295,0.5075723,0.45681506,0.40215343,0.3513962,0.30454338,0.26159495,0.21474212,0.1717937,0.12494087,0.1678893,0.21083772,0.25378615,0.29673457,0.3357786,0.7340276,1.1322767,1.5305257,1.9287747,2.3231194,4.084005,5.840986,7.5979667,9.354948,11.111929,11.795199,12.47847,13.16174,13.841106,14.524376,15.270117,16.015858,16.761599,17.503435,18.249176,16.644466,15.039758,13.435048,11.8303385,10.22563,9.761005,9.296382,8.831758,8.36323,7.898606,8.745861,9.597021,10.444276,11.291532,12.138786,1.5266213,1.6008049,1.678893,1.756981,1.8350691,1.9131571,1.9482968,1.9873407,2.0263848,2.0615244,2.1005683,2.182561,2.2645533,2.3465457,2.4285383,2.514435,2.5690966,2.6237583,2.67842,2.7330816,2.787743,2.951728,3.1118085,3.2757936,3.435874,3.5998588,4.0137253,4.4314966,4.845363,5.2592297,5.6730967,6.0713453,6.4695945,6.8678436,7.266093,7.6643414,6.481308,5.298274,4.11524,2.9322062,1.7491722,1.6008049,1.4485333,1.3001659,1.1517987,0.999527,0.8511597,0.698888,0.5505207,0.39824903,0.24988174,0.21864653,0.1835069,0.15227169,0.12103647,0.08589685,0.08980125,0.093705654,0.093705654,0.09761006,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.046852827,0.039044023,0.03513962,0.031235218,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.042948425,0.08589685,0.12884527,0.1717937,0.21083772,0.20693332,0.19912452,0.19131571,0.1835069,0.1756981,0.24988174,0.3240654,0.39824903,0.47633708,0.5505207,1.1869383,1.8233559,2.463678,3.1000953,3.736513,4.462732,5.1889505,5.911265,6.6374836,7.363703,7.0591593,6.7507114,6.446168,6.141625,5.8370814,5.364649,4.892216,4.4197836,3.9473507,3.474918,3.541293,3.611572,3.677947,3.7443218,3.8106966,4.466636,5.1225758,5.7785153,6.434455,7.08649,6.610153,6.133816,5.6535745,5.1772375,4.7009,4.661856,4.618908,4.579864,4.5408196,4.5017757,4.2597027,4.0215344,3.7794614,3.541293,3.2992198,2.639376,1.979532,1.319688,0.659844,0.0,0.46071947,0.92143893,1.3782539,1.8389735,2.2996929,3.0727646,3.8458362,4.618908,5.388075,6.1611466,6.0244927,5.8878384,5.7511845,5.610626,5.473972,5.5989127,5.7199492,5.840986,5.9659266,6.086963,6.3329406,6.578918,6.8209906,7.066968,7.3129454,6.7819467,6.250948,5.7238536,5.192855,4.661856,4.806319,4.950782,5.099149,5.2436123,5.388075,5.661383,5.938596,6.211904,6.4891167,6.7624245,7.2582836,7.7541428,8.246098,8.741957,9.237816,9.475985,9.714153,9.948417,10.186585,10.424754,10.295909,10.163159,10.034314,9.905469,9.776623,9.983557,10.19049,10.397423,10.604357,10.81129,10.865952,10.920613,10.979179,11.033841,11.088503,11.154878,11.221252,11.291532,11.357906,11.424281,11.545318,11.666354,11.783486,11.904523,12.025558,16.008049,19.99054,23.97303,27.95552,31.938011,40.633114,49.332123,58.03113,66.726234,75.42524,74.38277,73.340294,72.29781,71.25534,70.21287,64.653,59.09313,53.53326,47.97339,42.41352,40.2661,38.11868,35.971256,33.823837,31.676416,26.811531,21.946646,17.08176,12.212971,7.348085,7.406651,7.465217,7.523783,7.578445,7.6370106,11.92014,16.20327,20.486399,24.765623,29.048752,29.790588,30.53633,31.278166,32.020004,32.76184,33.671566,34.58129,35.491016,36.40074,37.314373,32.25427,27.198067,22.13796,17.08176,12.025558,14.832824,17.640089,20.447355,23.25462,26.061886,27.014559,27.967234,28.919907,29.872581,30.825256,28.748114,26.674877,24.601639,22.524496,20.45126,26.436708,32.41825,38.4037,44.38915,50.3746,43.756638,37.13477,30.512903,23.894941,17.273075,19.682093,22.091108,24.49622,26.905235,29.314253,24.464985,19.615717,14.770353,9.921086,5.0757227,5.883934,6.6960497,7.504261,8.316377,9.124588,9.600925,10.081166,10.557504,11.033841,11.514082,10.307622,9.101162,7.898606,6.6921453,5.4856853,6.192382,6.899079,7.601871,8.308568,9.01136,7.7814736,6.551587,5.3217,4.0918136,2.8619268,8.640442,14.418958,20.19357,25.972084,31.750599,29.493855,27.241014,24.98427,22.73143,20.474686,19.010534,17.550287,16.086138,14.625891,13.16174,12.435521,11.713207,10.986988,10.260769,9.538455,7.676055,5.813655,3.951255,2.0888553,0.22645533,2.194274,4.1581883,6.126007,8.093826,10.061645,10.662923,11.2642,11.861574,12.4628525,13.06413,14.141745,15.223265,16.300879,17.382399,18.463919,18.12033,17.776743,17.433157,17.093473,16.749886,16.199366,15.644939,15.0944195,14.539994,13.985569,11.66245,9.339331,7.012306,4.689187,2.3621633,3.4788225,4.591577,5.708236,6.8209906,7.9376497,8.921559,9.901564,10.885473,11.869383,12.849388,12.470661,12.091934,11.709302,11.330575,10.951848,9.913278,8.874706,7.8361354,6.801469,5.7628975,5.270943,4.7828927,4.290938,3.802888,3.310933,7.676055,12.041177,16.406298,20.77142,25.136541,21.528873,17.921206,14.313539,10.705871,7.098203,6.871748,6.6413884,6.4110284,6.180669,5.950309,5.196759,4.4393053,3.6857557,2.9283018,2.174752,2.4441557,2.7096553,2.979059,3.2445583,3.513962,3.9356375,4.357313,4.7789884,5.2006636,5.6262436,5.9268827,6.2314262,6.532065,6.8366084,7.137247,6.8951745,6.6531014,6.4110284,6.168956,5.9268827,6.1221027,6.321227,6.5164475,6.715572,6.910792,9.413514,11.916236,14.418958,16.921679,19.4244,17.538574,15.656653,13.770826,11.885,9.999174,9.030883,8.058686,7.0903945,6.1181984,5.1499066,4.8219366,4.493967,4.165997,3.8419318,3.513962,4.041056,4.5681505,5.095245,5.6223392,6.1494336,6.2314262,6.3134184,6.3993154,6.481308,6.5633,5.938596,5.3177958,4.6930914,4.0722914,3.4514916,2.7838387,2.1200905,1.456342,0.78868926,0.12494087,0.5661383,1.0112402,1.4524376,1.893635,2.338737,3.611572,4.8883114,6.1611466,7.437886,8.710721,7.4964523,6.278279,5.0601053,3.8419318,2.6237583,2.1005683,1.5734742,1.0502841,0.5231899,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.15617609,0.23816854,0.3240654,0.40605783,0.48805028,1.0268579,1.5656652,2.1083772,2.6471848,3.1859922,3.6935644,4.1972322,4.7009,5.2084727,5.7121406,6.785851,7.8556576,8.929368,10.003078,11.076789,10.475512,9.878138,9.280765,8.683391,8.086017,7.843944,7.5979667,7.3519893,7.1060123,6.8639393,7.098203,7.336372,7.57454,7.812709,8.050878,6.8873653,5.7238536,4.564246,3.4007344,2.2372224,2.0498111,1.8623998,1.6749885,1.4875772,1.3001659,1.2103647,1.1205635,1.0307622,0.94096094,0.8511597,0.8784905,0.9097257,0.94096094,0.96829176,0.999527,0.9058213,0.8160201,0.7223144,0.62860876,0.5388075,0.5505207,0.5622339,0.57394713,0.58566034,0.60127795,0.698888,0.79649806,0.8941081,0.9917182,1.0893283,1.1986516,1.3118792,1.4251068,1.5383345,1.6515622,1.5773785,1.5031948,1.4329157,1.358732,1.2884527,1.1947471,1.1010414,1.0112402,0.91753453,0.8238289,0.7145056,0.60518235,0.4958591,0.38653582,0.27330816,0.26549935,0.25378615,0.24597734,0.23426414,0.22645533,0.23426414,0.23816854,0.24597734,0.25378615,0.26159495,0.24597734,0.23426414,0.21864653,0.20302892,0.18741131,0.20693332,0.22645533,0.24597734,0.26940376,0.28892577,0.3240654,0.3631094,0.39824903,0.43729305,0.47633708,0.5622339,0.6481308,0.737932,0.8238289,0.9136301,0.97610056,1.038571,1.1010414,1.1635119,1.2259823,1.1205635,1.0151446,0.9097257,0.80430686,0.698888,0.59737355,0.4958591,0.39434463,0.28892577,0.18741131,0.21083772,0.23426414,0.25378615,0.27721256,0.30063897,0.60908675,0.9136301,1.2220778,1.5305257,1.8389735,3.1898966,4.5408196,5.8956475,7.2465706,8.601398,9.390087,10.178777,10.971371,11.760059,12.548749,13.501423,14.454097,15.406772,16.359446,17.31212,15.851873,14.391626,12.93138,11.471134,10.010887,9.655587,9.304191,8.94889,8.59359,8.238289,9.0465,9.850807,10.6590185,11.46723,12.27544,1.5383345,1.6086137,1.6827974,1.7530766,1.8272603,1.901444,1.9365835,1.9756275,2.0107672,2.0498111,2.0888553,2.1669433,2.2489357,2.3270237,2.4090161,2.4871042,2.5573835,2.6276627,2.697942,2.7682211,2.8385005,3.0259118,3.213323,3.4007344,3.5881457,3.775557,4.123049,4.4705405,4.8180323,5.165524,5.5130157,6.165051,6.817086,7.4691215,8.121157,8.773191,7.309041,5.840986,4.3729305,2.9048753,1.43682,1.2884527,1.1361811,0.9878138,0.8355421,0.6871748,0.60127795,0.5114767,0.42557985,0.3357786,0.24988174,0.21864653,0.19131571,0.16008049,0.12884527,0.10151446,0.10932326,0.12103647,0.12884527,0.14055848,0.14836729,0.14836729,0.14836729,0.14836729,0.14836729,0.14836729,0.13665408,0.12103647,0.10541886,0.08980125,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.058566034,0.113227665,0.1717937,0.23035973,0.28892577,0.28111696,0.27721256,0.27330816,0.26940376,0.26159495,0.37482262,0.48805028,0.60127795,0.7106012,0.8238289,1.7257458,2.6237583,3.5256753,4.423688,5.3256044,5.8370814,6.348558,6.8639393,7.375416,7.8868923,7.480835,7.0708723,6.6648145,6.2587566,5.8487945,5.4583545,5.0718184,4.6813784,4.290938,3.900498,3.7833657,3.6662338,3.5491016,3.4280653,3.310933,4.193328,5.0757227,5.958118,6.844417,7.726812,7.3519893,6.9810715,6.606249,6.2353306,5.8644123,5.840986,5.8175592,5.794133,5.7707067,5.7511845,5.1772375,4.60329,4.0332475,3.4593005,2.8892577,2.3114061,1.7335546,1.1557031,0.57785153,0.0,0.31625658,0.62860876,0.94486535,1.261122,1.5734742,2.5534792,3.5295796,4.50568,5.4856853,6.461786,6.239235,6.012779,5.786324,5.563773,5.337318,5.4271193,5.5169206,5.606722,5.6965227,5.786324,6.067441,6.348558,6.6257706,6.9068875,7.1880045,6.715572,6.2470436,5.7785153,5.3060827,4.8375545,5.169429,5.4973984,5.8292727,6.1572423,6.4891167,6.575013,6.66091,6.7507114,6.8366084,6.9264097,7.4691215,8.011833,8.550641,9.093353,9.636065,9.823476,10.010887,10.198298,10.38571,10.573121,10.518459,10.459893,10.401327,10.346666,10.2881,10.4286585,10.573121,10.71368,10.858143,10.998701,11.307149,11.615597,11.924045,12.228588,12.537036,12.658072,12.779109,12.89624,13.017277,13.138313,13.103174,13.0719385,13.040704,13.005564,12.974329,16.730364,20.486399,24.23853,27.994564,31.750599,41.253914,50.753326,60.25664,69.75996,79.26327,78.74399,78.220795,77.70151,77.18222,76.66294,70.49789,64.33283,58.167786,52.002735,45.83768,42.21049,38.5833,34.956112,31.328924,27.701735,23.4147,19.13157,14.844538,10.561408,6.2743745,6.453977,6.6335793,6.813182,6.996689,7.1762915,10.61607,14.059752,17.503435,20.943214,24.386896,26.33129,28.27568,30.223978,32.16837,34.112762,34.089336,34.06591,34.046387,34.02296,33.999535,29.78278,25.566027,21.349272,17.128613,12.911859,15.356014,17.796265,20.240421,22.680674,25.124828,25.671444,26.218061,26.768581,27.315199,27.861814,26.41328,24.960844,23.51231,22.063778,20.61134,26.2532,31.891157,37.53302,43.170975,48.812836,42.370575,35.92831,29.486046,23.043781,16.601519,18.94416,21.2868,23.629442,25.96818,28.310822,23.785618,19.256512,14.73131,10.202203,5.6730967,6.914696,8.156297,9.393991,10.6355915,11.873287,12.373051,12.86891,13.368673,13.864532,14.364296,12.790822,11.221252,9.651682,8.082112,6.5125427,6.5828223,6.6531014,6.7233806,6.79366,6.8639393,6.3173227,5.7707067,5.2279944,4.6813784,4.138666,8.898132,13.657599,18.417065,23.176533,27.935999,25.815908,23.695818,21.575727,19.455637,17.335546,16.800642,16.261835,15.723028,15.188125,14.649317,13.224211,11.799104,10.373997,8.94889,7.523783,6.0518236,4.575959,3.1000953,1.6242313,0.14836729,2.3699722,4.591577,6.8092775,9.030883,11.248583,12.8767185,14.50095,16.125181,17.749413,19.373644,20.209187,21.040823,21.872461,22.7041,23.535736,23.078922,22.622107,22.16529,21.708477,21.251661,19.525915,17.804073,16.082233,14.360392,12.63855,10.424754,8.210958,6.001066,3.78727,1.5734742,3.5725281,5.571582,7.5667315,9.565785,11.560935,12.716639,13.872341,15.028045,16.183748,17.33945,17.155943,16.972437,16.788929,16.609327,16.42582,14.13784,11.849861,9.561881,7.2739015,4.985922,4.6267166,4.267512,3.9083066,3.5491016,3.1859922,7.6721506,12.158309,16.644466,21.12672,25.612879,21.618675,17.628376,13.634172,9.643873,5.64967,5.7316628,5.8097506,5.891743,5.969831,6.0518236,5.2045684,4.3612175,3.513962,2.6706111,1.8233559,2.2840753,2.7408905,3.1977055,3.6545205,4.1113358,4.552533,4.9937305,5.4310236,5.872221,6.3134184,6.5867267,6.8561306,7.1294384,7.4027467,7.676055,7.266093,6.860035,6.453977,6.044015,5.6379566,5.9542136,6.266566,6.5828223,6.899079,7.211431,9.846903,12.482374,15.117846,17.753317,20.388788,18.51077,16.632753,14.754736,12.8767185,10.998701,9.8429985,8.691199,7.535496,6.379793,5.22409,5.0913405,4.9546866,4.8219366,4.6852827,4.548629,4.8102236,5.0718184,5.3295093,5.591104,5.8487945,5.7668023,5.6848097,5.602817,5.520825,5.4388323,5.0601053,4.6813784,4.3065557,3.9278288,3.5491016,2.8775444,2.2059872,1.53443,0.8589685,0.18741131,0.71841,1.2533131,1.7843118,2.3192148,2.8502135,3.9629683,5.0757227,6.1884775,7.3012323,8.413987,7.3051367,6.196286,5.0913405,3.9824903,2.87364,2.2996929,1.7257458,1.1517987,0.57394713,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.1678893,0.28502136,0.40215343,0.5192855,0.63641757,1.4212024,2.2059872,2.9907722,3.7794614,4.564246,4.493967,4.4275923,4.3612175,4.290938,4.224563,5.45445,6.6804323,7.9064145,9.136301,10.362284,9.421323,8.484266,7.5433054,6.602344,5.661383,5.5091114,5.3529353,5.196759,5.040583,4.8883114,5.0640097,5.2358036,5.4115014,5.5871997,5.7628975,4.9234514,4.087909,3.2484627,2.4129205,1.5734742,1.43682,1.3001659,1.1635119,1.0268579,0.8862993,0.8277333,0.76916724,0.7066968,0.6481308,0.58566034,0.6559396,0.7262188,0.79649806,0.8667773,0.93705654,0.8550641,0.77307165,0.6910792,0.60908675,0.5231899,0.5622339,0.60127795,0.63641757,0.6754616,0.7106012,0.76526284,0.8160201,0.8706817,0.92143893,0.97610056,1.0268579,1.0737107,1.1244678,1.175225,1.2259823,1.1596074,1.0932326,1.0307622,0.96438736,0.9019169,0.8433509,0.78478485,0.7262188,0.6715572,0.61299115,0.5466163,0.48414588,0.41777104,0.3513962,0.28892577,0.28502136,0.28111696,0.28111696,0.27721256,0.27330816,0.28111696,0.28502136,0.28892577,0.29673457,0.30063897,0.27721256,0.25378615,0.23426414,0.21083772,0.18741131,0.21864653,0.24597734,0.27721256,0.30844778,0.3357786,0.39824903,0.46071947,0.5231899,0.58566034,0.6481308,0.78868926,0.92534333,1.0619974,1.1986516,1.33921,1.43682,1.5383345,1.6359446,1.737459,1.8389735,1.678893,1.5227169,1.3665408,1.2064602,1.0502841,0.8902037,0.7301232,0.5700427,0.40996224,0.24988174,0.25378615,0.25378615,0.25769055,0.26159495,0.26159495,0.48024148,0.698888,0.9136301,1.1322767,1.3509232,2.2957885,3.2445583,4.193328,5.138193,6.086963,6.984976,7.882988,8.781001,9.679013,10.573121,11.736633,12.89624,14.055848,15.215456,16.375063,15.059279,13.743496,12.431617,11.115833,9.80005,9.554072,9.308095,9.066022,8.8200445,8.574067,9.343235,10.108498,10.877665,11.6468315,12.412095,1.5500476,1.6164225,1.6867018,1.7530766,1.8194515,1.8858263,1.9248703,1.9639144,1.999054,2.0380979,2.0732377,2.1513257,2.2294137,2.3075018,2.3855898,2.463678,2.5456703,2.631567,2.717464,2.803361,2.8892577,3.1000953,3.310933,3.5256753,3.736513,3.951255,4.2284675,4.5095844,4.7907014,5.0718184,5.349031,6.2587566,7.164578,8.074304,8.980125,9.885946,8.136774,6.3836975,4.630621,2.8775444,1.1244678,0.97610056,0.8238289,0.6754616,0.5231899,0.37482262,0.3513962,0.3240654,0.30063897,0.27330816,0.24988174,0.22255093,0.19522011,0.1678893,0.14055848,0.113227665,0.12884527,0.14836729,0.1639849,0.1835069,0.19912452,0.19912452,0.19912452,0.19912452,0.19912452,0.19912452,0.1796025,0.16008049,0.14055848,0.12103647,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.07418364,0.14446288,0.21864653,0.28892577,0.3631094,0.359205,0.359205,0.3553006,0.3513962,0.3513962,0.4997635,0.6481308,0.80040246,0.94876975,1.1010414,2.260649,3.4241607,4.5876727,5.7511845,6.910792,7.211431,7.5120697,7.812709,8.113348,8.413987,7.90251,7.3910336,6.883461,6.3719845,5.8644123,5.5559645,5.2475166,4.939069,4.630621,4.3260775,4.0215344,3.7208953,3.416352,3.1157131,2.8111696,3.9239242,5.0327744,6.141625,7.2543793,8.36323,8.093826,7.8283267,7.558923,7.2934237,7.0240197,7.0201154,7.016211,7.008402,7.0044975,7.000593,6.094772,5.1889505,4.283129,3.3812122,2.475391,1.979532,1.4836729,0.9917182,0.4958591,0.0,0.1717937,0.339683,0.5114767,0.679366,0.8511597,2.0341935,3.213323,4.396357,5.579391,6.7624245,6.4500723,6.13772,5.825368,5.5130157,5.2006636,5.2592297,5.3138914,5.3724575,5.4310236,5.4856853,5.801942,6.1181984,6.434455,6.746807,7.0630636,6.6531014,6.2431393,5.833177,5.423215,5.0132523,5.5286336,6.044015,6.559396,7.0708723,7.5862536,7.4886436,7.387129,7.2856145,7.1880045,7.08649,7.676055,8.265619,8.859089,9.448653,10.0382185,10.174872,10.311526,10.44818,10.588739,10.725393,10.741011,10.756628,10.768341,10.783959,10.799577,10.877665,10.955752,11.033841,11.111929,11.186112,11.748346,12.306676,12.86891,13.427239,13.985569,14.161267,14.33306,14.504854,14.676648,14.848442,14.664935,14.481428,14.294017,14.11051,13.923099,17.452679,20.978354,24.507933,28.033607,31.563189,41.87081,52.178432,62.486053,72.79368,83.101295,83.101295,83.1052,83.10911,83.10911,83.113014,76.34278,69.57254,62.80231,56.032078,49.261845,44.154884,39.047928,33.940968,28.834011,23.723148,20.021774,16.316498,12.611219,8.905942,5.2006636,5.5013027,5.805846,6.1064854,6.4110284,6.7116675,9.315904,11.916236,14.520472,17.120804,5052.0,22.871988,26.018936,29.165884,32.31674,35.463684,34.507107,33.554432,32.597855,31.641275,30.688602,27.311295,23.933987,20.556679,17.17937,13.798158,15.879204,17.956347,20.033487,22.11063,24.187773,24.328331,24.472794,24.613352,24.757814,24.898373,24.074545,23.250715,22.426888,21.599154,20.775324,26.069695,31.364063,36.658432,41.956707,47.251076,40.984512,34.721848,28.455284,22.188719,15.926057,18.202324,20.47859,22.75876,25.035027,27.311295,23.106253,18.897306,14.688361,10.48332,6.2743745,7.9454584,9.616543,11.283723,12.954806,14.625891,15.141272,15.660558,16.175938,16.695225,17.210606,15.277926,13.341343,11.408664,9.47208,7.5394006,6.9732623,6.407124,5.840986,5.278752,4.7126136,4.853172,4.9937305,5.134289,5.270943,5.4115014,9.155824,12.89624,16.640562,20.38098,24.125301,22.13796,20.154524,18.171087,16.183748,14.200311,14.586847,14.973383,15.363823,15.750359,16.136894,14.012899,11.888905,9.761005,7.6370106,5.5130157,4.423688,3.338264,2.2489357,1.1635119,0.07418364,2.5495746,5.0210614,7.492548,9.964035,12.439425,15.086611,17.7377,20.388788,23.035973,25.687063,26.272722,26.858383,27.444044,28.025799,28.61146,28.041416,27.46747,26.893522,26.32348,25.749533,22.85637,19.96321,17.073952,14.180789,11.287627,9.187058,7.08649,4.985922,2.8892577,0.78868926,3.6662338,6.547683,9.4291315,12.306676,15.188125,16.515621,17.843119,19.170614,20.498112,21.82561,21.841227,21.856844,21.868557,21.884174,21.899792,18.362404,14.825015,11.287627,7.7502384,4.21285,3.9824903,3.7521305,3.521771,3.2914112,3.0610514,7.6682463,12.271536,16.87873,21.482021,26.089216,21.708477,17.331642,12.954806,8.577971,4.2011366,4.591577,4.9781127,5.368553,5.758993,6.1494336,5.2162814,4.279225,3.3460727,2.4090161,1.475864,2.1239948,2.7682211,3.416352,4.0644827,4.7126136,5.169429,5.6262436,6.086963,6.5437784,7.000593,7.2426662,7.4847393,7.726812,7.968885,8.210958,7.6409154,7.066968,6.4969254,5.9229784,5.349031,5.7824197,6.2158084,6.649197,7.0786815,7.5120697,10.280292,13.048512,15.816733,18.58105,21.349272,19.479063,17.608854,15.738646,13.868437,11.998228,10.6590185,9.319808,7.9805984,6.6413884,5.298274,5.35684,5.4154058,5.473972,5.5286336,5.5871997,5.579391,5.571582,5.563773,5.5559645,5.548156,5.3021784,5.056201,4.806319,4.560342,4.3143644,4.181615,4.0488653,3.9161155,3.7833657,3.6506162,2.97125,2.2918842,1.6086137,0.92924774,0.24988174,0.8706817,1.4953861,2.1161861,2.7408905,3.3616903,4.3143644,5.263134,6.211904,7.1606736,8.113348,7.113821,6.1181984,5.1186714,4.123049,3.1235218,2.4988174,1.8741131,1.2494087,0.62470436,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.1756981,0.3318742,0.48414588,0.63641757,0.78868926,1.8194515,2.8463092,3.8770714,4.9078336,5.938596,5.298274,4.657952,4.01763,3.377308,2.736986,4.1191444,5.5013027,6.883461,8.265619,9.651682,8.367134,7.08649,5.801942,4.521298,3.2367494,3.174279,3.1079042,3.0415294,2.979059,2.912684,3.0259118,3.1391394,3.2484627,3.3616903,3.474918,2.9634414,2.4519646,1.9365835,1.4251068,0.9136301,0.8238289,0.737932,0.6481308,0.5622339,0.47633708,0.44510186,0.41386664,0.38653582,0.3553006,0.3240654,0.43338865,0.5466163,0.6559396,0.76526284,0.8745861,0.80430686,0.7301232,0.6559396,0.58566034,0.5114767,0.57394713,0.63641757,0.698888,0.76135844,0.8238289,0.8316377,0.8394465,0.8472553,0.8550641,0.8628729,0.8511597,0.8394465,0.8238289,0.81211567,0.80040246,0.7418364,0.6832704,0.62860876,0.5700427,0.5114767,0.48805028,0.46852827,0.44510186,0.42167544,0.39824903,0.37872702,0.359205,0.339683,0.32016098,0.30063897,0.30454338,0.30844778,0.31625658,0.32016098,0.3240654,0.3279698,0.3318742,0.3318742,0.3357786,0.3357786,0.30844778,0.27721256,0.24597734,0.21864653,0.18741131,0.22645533,0.26940376,0.30844778,0.3474918,0.38653582,0.47633708,0.5622339,0.6481308,0.737932,0.8238289,1.0112402,1.1986516,1.3860629,1.5734742,1.7608855,1.901444,2.0380979,2.174752,2.3114061,2.4480603,2.241127,2.0302892,1.8194515,1.6086137,1.4016805,1.183034,0.96438736,0.74574083,0.5309987,0.31235218,0.29673457,0.27721256,0.26159495,0.24207294,0.22645533,0.3513962,0.48024148,0.60908675,0.7340276,0.8628729,1.4055848,1.9482968,2.4910088,3.0337205,3.5764325,4.579864,5.5832953,6.590631,7.5940623,8.601398,9.967939,11.334479,12.70102,14.0714655,15.438006,14.2666855,13.09927,11.927949,10.756628,9.589212,9.452558,9.315904,9.183154,9.0465,8.913751,9.639969,10.366188,11.096312,11.82253,12.548749,1.5617609,1.6242313,1.6867018,1.7491722,1.8116426,1.8741131,1.9131571,1.9482968,1.9873407,2.0263848,2.0615244,2.135708,2.2137961,2.2879796,2.3621633,2.436347,2.5378613,2.639376,2.736986,2.8385005,2.9361105,3.174279,3.4124475,3.6506162,3.8887846,4.123049,4.337791,4.548629,4.7633705,4.9742084,5.1889505,6.348558,7.5120697,8.675582,9.839094,10.998701,8.960603,6.9264097,4.8883114,2.8502135,0.81211567,0.6637484,0.5114767,0.3631094,0.21083772,0.062470436,0.10151446,0.13665408,0.1756981,0.21083772,0.24988174,0.22645533,0.19912452,0.1756981,0.14836729,0.12494087,0.14836729,0.1756981,0.19912452,0.22645533,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.22645533,0.19912452,0.1756981,0.14836729,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.43729305,0.43729305,0.43729305,0.43729305,0.43729305,0.62470436,0.81211567,0.999527,1.1869383,1.3743496,2.7994564,4.224563,5.64967,7.0747766,8.499884,8.58578,8.675582,8.761478,8.85128,8.937177,8.324185,7.7111945,7.098203,6.4891167,5.8761253,5.64967,5.423215,5.2006636,4.9742084,4.7516575,4.263607,3.775557,3.2875066,2.7994564,2.3114061,3.6506162,4.985922,6.3251314,7.6643414,8.999647,8.835662,8.675582,8.511597,8.351517,8.187531,8.1992445,8.210958,8.226576,8.238289,8.250002,7.012306,5.774611,4.5369153,3.2992198,2.0615244,1.6515622,1.2376955,0.8238289,0.41386664,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,1.5110037,2.900971,4.2870336,5.6730967,7.0630636,6.66091,6.262661,5.8644123,5.462259,5.0640097,5.087436,5.1108627,5.138193,5.1616197,5.1889505,5.5364423,5.8878384,6.239235,6.5867267,6.9381227,6.5867267,6.239235,5.8878384,5.5364423,5.1889505,5.8878384,6.5867267,7.2856145,7.988407,8.687295,8.398369,8.113348,7.824422,7.5394006,7.250475,7.8868923,8.52331,9.163632,9.80005,10.436467,10.526268,10.612165,10.698062,10.787864,10.87376,10.963562,11.0494585,11.139259,11.225157,11.311053,11.326671,11.338385,11.350098,11.361811,11.373524,12.185639,13.001659,13.813775,14.625891,15.438006,15.660558,15.8870125,16.113468,16.33602,16.562475,16.226696,15.8870125,15.551234,15.211552,14.875772,18.174992,21.474213,24.773432,28.076557,31.375776,42.487705,53.599632,64.71156,75.823494,86.93932,87.46252,87.9857,88.5128,89.03599,89.56308,82.18767,74.81225,67.43684,60.06142,52.686005,46.099277,39.51255,32.925823,26.339098,19.748466,16.624945,13.501423,10.373997,7.250475,4.123049,4.548629,4.9742084,5.3997884,5.825368,6.250948,8.011833,9.776623,11.537509,13.298394,15.063184,19.412687,23.762192,28.111696,32.4612,36.810703,34.924877,33.03905,31.14932,29.263494,27.373764,24.835903,22.301945,19.764084,17.226223,14.688361,16.398489,18.112522,19.826555,21.536682,23.250715,22.98912,22.723621,22.462027,22.200432,21.938837,21.735807,21.536682,21.337559,21.138433,20.93931,25.886187,30.83697,35.78775,40.738533,45.689316,39.598446,33.511486,27.424522,21.337559,15.250595,17.464392,19.674282,21.888079,24.101875,26.311768,22.426888,18.538101,14.649317,10.760532,6.8756523,8.976221,11.076789,13.173453,15.274021,17.37459,17.913397,18.448301,18.987108,19.525915,20.06082,17.761126,15.461433,13.16174,10.862047,8.562354,7.363703,6.1611466,4.9624953,3.7638438,2.5612879,3.3890212,4.21285,5.036679,5.8644123,6.688241,9.413514,12.138786,14.864059,17.589333,20.310701,18.463919,16.613232,14.762545,12.911859,11.061172,12.376955,13.688834,15.000713,16.312593,17.624472,14.801589,11.974802,9.148014,6.3251314,3.4983444,2.7994564,2.1005683,1.4016805,0.698888,0.0,2.7252727,5.4505453,8.175818,10.901091,13.626364,17.300406,20.97445,24.64849,28.326439,32.00048,32.336258,32.67594,33.011723,33.351402,33.687183,33.000008,32.31283,31.625658,30.938484,30.251308,26.186827,22.126247,18.061766,14.001186,9.936704,7.9493628,5.9620223,3.9746814,1.9873407,0.0,3.7638438,7.523783,11.287627,15.051471,18.81141,20.310701,21.813896,23.313187,24.812477,26.311768,26.526508,26.737347,26.948185,27.162926,27.373764,22.586967,17.800169,13.013372,8.226576,3.435874,3.338264,3.2367494,3.1391394,3.0376248,2.9361105,7.6643414,12.388668,17.112995,21.837322,26.56165,21.798277,17.03881,12.27544,7.5120697,2.7486992,3.4514916,4.1503797,4.8492675,5.548156,6.250948,5.22409,4.2011366,3.174279,2.1513257,1.1244678,1.9639144,2.7994564,3.638903,4.474445,5.3138914,5.786324,6.262661,6.7389984,7.211431,7.687768,7.898606,8.113348,8.324185,8.538928,8.749765,8.011833,7.2739015,6.5359693,5.7980375,5.0640097,5.610626,6.1611466,6.7116675,7.262188,7.812709,10.71368,13.610746,16.511717,19.412687,22.31366,20.45126,18.58886,16.72646,14.864059,13.001659,11.475039,9.948417,8.4257,6.899079,5.376362,5.6262436,5.8761253,6.126007,6.375889,6.6257706,6.348558,6.0752497,5.801942,5.5247293,5.251421,4.8375545,4.423688,4.0137253,3.5998588,3.1859922,3.2992198,3.4124475,3.5256753,3.638903,3.7482262,3.0610514,2.3738766,1.6867018,0.999527,0.31235218,1.0268579,1.737459,2.4519646,3.1625657,3.873167,4.661856,5.4505453,6.239235,7.0240197,7.812709,6.9264097,6.036206,5.1499066,4.263607,3.3734035,2.7018464,2.0263848,1.3509232,0.6754616,0.0,0.0,0.0,0.0,0.0,0.0,0.18741131,0.37482262,0.5622339,0.74964523,0.93705654,2.2137961,3.4866312,4.7633705,6.036206,7.3129454,6.098676,4.8883114,3.6740425,2.463678,1.2494087,2.787743,4.3260775,5.8644123,7.3988423,8.937177,7.3129454,5.688714,4.0605783,2.436347,0.81211567,0.8394465,0.8628729,0.8862993,0.9136301,0.93705654,0.9878138,1.038571,1.0893283,1.1361811,1.1869383,0.999527,0.81211567,0.62470436,0.43729305,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.21083772,0.3631094,0.5114767,0.6637484,0.81211567,0.74964523,0.6871748,0.62470436,0.5622339,0.4997635,0.58566034,0.6754616,0.76135844,0.8511597,0.93705654,0.9019169,0.8628729,0.8238289,0.78868926,0.74964523,0.6754616,0.60127795,0.5231899,0.44900626,0.37482262,0.3240654,0.27330816,0.22645533,0.1756981,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.21083772,0.23816854,0.26159495,0.28892577,0.31235218,0.3240654,0.3357786,0.3513962,0.3631094,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.3357786,0.30063897,0.26159495,0.22645533,0.18741131,0.23816854,0.28892577,0.3357786,0.38653582,0.43729305,0.5505207,0.6637484,0.77307165,0.8862993,0.999527,1.2376955,1.475864,1.7140326,1.9482968,2.1864653,2.3621633,2.5378613,2.7135596,2.8892577,3.0610514,2.7994564,2.5378613,2.2762666,2.0107672,1.7491722,1.475864,1.1986516,0.92534333,0.6481308,0.37482262,0.3357786,0.30063897,0.26159495,0.22645533,0.18741131,0.22645533,0.26159495,0.30063897,0.3357786,0.37482262,0.5114767,0.6481308,0.78868926,0.92534333,1.0619974,2.174752,3.2875066,4.4002614,5.5130157,6.6257706,8.1992445,9.776623,11.350098,12.923572,14.50095,13.4740925,12.4511385,11.424281,10.401327,9.37447,9.351044,9.323712,9.300286,9.276859,9.249529,9.936704,10.6238785,11.311053,11.998228,12.689307,1.5617609,1.6242313,1.6827974,1.7413634,1.8038338,1.8623998,1.901444,1.9443923,1.9834363,2.0224805,2.0615244,2.135708,2.2137961,2.2879796,2.3621633,2.436347,2.5534792,2.6706111,2.7916477,2.9087796,3.0259118,3.232845,3.4397783,3.6467118,3.853645,4.0605783,4.318269,4.572055,4.825841,5.083532,5.337318,6.27047,7.2036223,8.136774,9.066022,9.999174,8.207053,6.4149327,4.6228123,2.8306916,1.038571,0.8511597,0.6676528,0.48414588,0.29673457,0.113227665,0.13274968,0.15227169,0.1717937,0.19131571,0.21083772,0.19912452,0.18741131,0.1756981,0.1639849,0.14836729,0.1639849,0.1796025,0.19522011,0.21083772,0.22645533,0.22255093,0.21864653,0.21864653,0.21474212,0.21083772,0.19131571,0.1678893,0.14446288,0.12103647,0.10151446,0.093705654,0.08589685,0.078088045,0.07027924,0.062470436,0.06637484,0.06637484,0.07027924,0.07418364,0.07418364,0.1678893,0.26159495,0.3513962,0.44510186,0.5388075,0.5466163,0.5583295,0.5661383,0.57785153,0.58566034,1.2494087,1.9092526,2.5690966,3.2289407,3.8887846,5.114767,6.3407493,7.570636,8.796618,10.0265045,9.956225,9.885946,9.815667,9.745388,9.675109,8.831758,7.984503,7.141152,6.2938967,5.4505453,5.270943,5.095245,4.9156423,4.7399445,4.564246,4.1581883,3.7521305,3.3460727,2.9439192,2.5378613,3.638903,4.743849,5.84489,6.9459314,8.050878,7.957172,7.8634663,7.773665,7.6799593,7.5862536,7.7541428,7.9220324,8.089922,8.257811,8.4257,7.1216297,5.813655,4.5095844,3.2055142,1.901444,1.5188124,1.1400855,0.76135844,0.37872702,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,1.5890918,3.0805733,4.5681505,6.0596323,7.551114,6.89127,6.2314262,5.571582,4.911738,4.251894,4.4900627,4.728231,4.970304,5.2084727,5.4505453,5.7511845,6.0518236,6.348558,6.649197,6.949836,6.606249,6.2587566,5.9151692,5.571582,5.22409,5.786324,6.348558,6.910792,7.47693,8.039165,7.882988,7.726812,7.570636,7.4183645,7.262188,7.843944,8.421796,9.0035515,9.581403,10.163159,10.108498,10.05774,10.003078,9.952321,9.901564,10.085071,10.268578,10.455989,10.639496,10.826907,10.881569,10.936231,10.990892,11.045554,11.100216,11.927949,12.755682,13.583415,14.411149,15.238882,15.410676,15.586374,15.762072,15.93777,16.113468,15.863586,15.617609,15.371632,15.12175,14.875772,17.854832,20.83389,23.816854,26.795912,29.774971,40.07869,50.38631,60.69003,70.993744,81.30137,82.94512,84.588875,86.236534,87.88029,89.52404,82.07444,74.62093,67.167435,59.71393,52.264328,45.029472,37.79852,30.563662,23.332708,16.101755,13.708356,11.314958,8.921559,6.5281606,4.138666,4.5017757,4.8687897,5.2318993,5.5989127,5.9620223,7.656533,9.351044,11.0494585,12.743969,14.438479,18.58886,22.739239,26.885714,31.036093,35.186474,32.67594,30.169315,27.658785,25.148254,22.637724,20.954927,19.27213,17.589333,15.906535,14.223738,15.293544,16.359446,17.429253,18.495153,19.561056,19.354122,19.147188,18.940256,18.733322,18.526388,20.462973,22.399555,24.33614,26.276627,28.213211,32.05124,35.889267,39.72339,43.561417,47.399445,41.101643,34.79994,28.498232,22.200432,15.8987255,17.929016,19.9554,21.981785,24.00817,26.038458,22.551826,19.069101,15.582469,12.095839,8.6131115,10.049932,11.486752,12.923572,14.364296,15.801116,16.277452,16.75379,17.234032,17.71037,18.186707,16.41801,14.653222,12.884527,11.115833,9.351044,8.160201,6.969358,5.7785153,4.591577,3.4007344,4.6384296,5.8800297,7.1216297,8.359325,9.600925,11.881096,14.161267,16.441439,18.72161,21.00178,18.9793,16.960724,14.938243,12.919667,10.901091,13.345247,15.789403,18.233559,20.68162,23.125774,19.514202,15.906535,12.294963,8.683391,5.0757227,4.5993857,4.126953,3.6506162,3.174279,2.7018464,4.985922,7.2739015,9.561881,11.849861,14.13784,17.366781,20.591818,23.820759,27.045794,30.274734,31.301594,32.32845,33.359215,34.38607,35.41293,34.514915,33.616905,32.71889,31.820879,30.926771,26.874,22.825136,18.77627,14.723501,10.674636,8.542832,6.4110284,4.279225,2.1435168,0.011713207,3.6467118,7.277806,10.9089,14.543899,18.174992,5052.0,21.275087,22.825136,24.375183,25.925232,26.054077,26.186827,26.315672,26.444517,26.573362,22.07549,17.581524,13.083652,8.58578,4.087909,3.9434462,3.7989833,3.6506162,3.506153,3.3616903,7.08649,10.807385,14.528281,18.25308,21.973976,18.073479,14.176885,10.276386,6.375889,2.475391,3.533484,4.591577,5.645766,6.703859,7.7619514,7.0513506,6.3407493,5.6340523,4.9234514,4.21285,4.9820175,5.7511845,6.524256,7.2934237,8.062591,8.105539,8.148487,8.191436,8.234385,8.273428,8.488171,8.699008,8.913751,9.124588,9.339331,8.433509,7.531592,6.629675,5.727758,4.825841,5.3529353,5.8800297,6.407124,6.9342184,7.461313,9.788337,12.111456,14.438479,16.761599,19.088623,17.491722,15.8987255,14.301826,12.708829,11.111929,9.897659,8.683391,7.4691215,6.250948,5.036679,5.290465,5.5442514,5.794133,6.0479193,6.3017054,5.930787,5.559869,5.1889505,4.8219366,4.4510183,4.21285,3.9746814,3.736513,3.4983444,3.2640803,3.2289407,3.1977055,3.1664703,3.1313305,3.1000953,2.5612879,2.018576,1.4797685,0.94096094,0.39824903,0.97219616,1.5461433,2.1161861,2.690133,3.2640803,3.8614538,4.4588275,5.056201,5.6535745,6.250948,5.6926184,5.134289,4.575959,4.0215344,3.4632049,2.8345962,2.2059872,1.5812829,0.95267415,0.3240654,0.26940376,0.21083772,0.15227169,0.093705654,0.039044023,0.77697605,1.5188124,2.2567444,2.998581,3.736513,4.165997,4.591577,5.0210614,5.446641,5.8761253,5.267039,4.661856,4.0527697,3.4436827,2.8385005,3.7794614,4.7243266,5.6652875,6.606249,7.551114,6.168956,4.7907014,3.408543,2.0302892,0.6481308,0.6754616,0.698888,0.7262188,0.74964523,0.77307165,0.8160201,0.8550641,0.8941081,0.93315214,0.97610056,0.97610056,0.97610056,0.97610056,0.97610056,0.97610056,0.98390937,0.9917182,0.9956226,1.0034313,1.0112402,0.92924774,0.8433509,0.75745404,0.6715572,0.58566034,0.7418364,0.8980125,1.0541886,1.2064602,1.3626363,1.2650263,1.1674163,1.0698062,0.97219616,0.8745861,0.8706817,0.8706817,0.8667773,0.8667773,0.8628729,0.8277333,0.79259366,0.75745404,0.7223144,0.6871748,0.62079996,0.5544251,0.48414588,0.41777104,0.3513962,0.30844778,0.26549935,0.22255093,0.1796025,0.13665408,0.16008049,0.1835069,0.20693332,0.22645533,0.24988174,0.28111696,0.30844778,0.339683,0.3709182,0.39824903,0.39824903,0.39434463,0.39434463,0.39044023,0.38653582,0.41386664,0.44119745,0.46852827,0.4958591,0.5231899,0.5544251,0.58175594,0.60908675,0.63641757,0.6637484,0.8160201,0.97219616,1.1283722,1.2806439,1.43682,1.53443,1.6281357,1.7218413,1.815547,1.9131571,2.2684577,2.6276627,2.9868677,3.3421683,3.7013733,3.8458362,3.9902992,4.134762,4.279225,4.423688,4.185519,3.9434462,3.7052777,3.4632049,3.2250361,3.0883822,2.951728,2.8111696,2.6745155,2.5378613,2.5651922,2.592523,2.619854,2.6471848,2.6745155,2.4597735,2.2450314,2.0302892,1.815547,1.6008049,1.5070993,1.4133936,1.3235924,1.2298868,1.1361811,2.069333,2.998581,3.9278288,4.8570766,5.786324,7.1841,8.581876,9.979652,11.377428,12.775204,11.924045,11.06898,10.217821,9.366661,8.511597,8.597494,8.683391,8.769287,8.85128,8.937177,9.643873,10.354475,11.061172,11.767868,12.4745655,1.5617609,1.620327,1.678893,1.7335546,1.7921207,1.8506867,1.893635,1.9365835,1.9756275,2.018576,2.0615244,2.135708,2.2137961,2.2879796,2.3621633,2.436347,2.5730011,2.7057507,2.8424048,2.979059,3.1118085,3.2914112,3.4671092,3.6467118,3.8224099,3.998108,4.298747,4.5954814,4.892216,5.1889505,5.4856853,6.1884775,6.89127,7.5940623,8.296855,8.999647,7.453504,5.903456,4.357313,2.8111696,1.261122,1.0424755,0.8238289,0.60127795,0.38263142,0.1639849,0.1639849,0.1678893,0.1717937,0.1717937,0.1756981,0.1756981,0.1756981,0.1756981,0.1756981,0.1756981,0.1796025,0.1835069,0.19131571,0.19522011,0.19912452,0.19522011,0.19131571,0.1835069,0.1796025,0.1756981,0.15617609,0.13665408,0.113227665,0.093705654,0.07418364,0.07418364,0.07027924,0.06637484,0.06637484,0.062470436,0.078088045,0.09761006,0.113227665,0.13274968,0.14836729,0.24597734,0.3435874,0.44119745,0.5388075,0.63641757,0.6559396,0.679366,0.698888,0.71841,0.737932,1.8702087,3.0024853,4.134762,5.267039,6.3993154,7.4300776,8.460839,9.491602,10.518459,11.549222,11.322766,11.096312,10.865952,10.639496,10.413041,9.335425,8.257811,7.180196,6.1025805,5.024966,4.8961205,4.7633705,4.6345253,4.50568,4.376835,4.0527697,3.7287042,3.408543,3.084478,2.7643168,3.631094,4.4978714,5.364649,6.2314262,7.098203,7.0786815,7.055255,7.0318284,7.008402,6.98888,7.309041,7.633106,7.9532676,8.277332,8.601398,7.2270484,5.8566036,4.482254,3.1118085,1.737459,1.3899672,1.0424755,0.6949836,0.3474918,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,1.6671798,3.260176,4.853172,6.446168,8.039165,7.1177254,6.196286,5.278752,4.357313,3.435874,3.892689,4.3455997,4.802415,5.2592297,5.7121406,5.9620223,6.211904,6.461786,6.7116675,6.9615493,6.621866,6.282183,5.9425,5.602817,5.263134,5.688714,6.114294,6.5359693,6.9615493,7.387129,7.363703,7.3441806,7.320754,7.297328,7.2739015,7.7970915,8.320281,8.843472,9.366661,9.885946,9.694631,9.503315,9.308095,9.116779,8.925464,9.20658,9.491602,9.772718,10.053836,10.338858,10.436467,10.534078,10.631687,10.729298,10.826907,11.666354,12.509705,13.353056,14.196406,15.035853,15.160794,15.285735,15.410676,15.535617,15.660558,15.504381,15.348206,15.188125,15.031949,14.875772,17.53467,20.19357,22.85637,25.515268,28.174168,37.673576,47.169083,56.668495,66.164,75.663414,78.42773,81.19205,83.95636,86.72068,89.4889,81.957306,74.42962,66.898026,59.366436,51.83875,43.959663,36.084484,28.205402,20.326319,12.4511385,10.791768,9.128492,7.4691215,5.8097506,4.1503797,4.454923,4.759466,5.0640097,5.368553,5.6730967,7.3012323,8.929368,10.557504,12.185639,13.813775,17.761126,21.712381,25.663635,29.610987,33.56224,30.430912,27.295675,24.164345,21.033014,17.901684,17.073952,16.246218,15.418485,14.590752,13.763018,14.184693,14.606369,15.028045,15.453624,15.875299,15.723028,15.570756,15.418485,15.266212,15.113941,19.186234,23.262428,27.338625,31.410915,35.487114,38.212383,40.937656,43.66293,46.388203,49.113476,42.600933,36.08839,29.575848,23.063305,16.55076,18.393639,20.236517,22.079395,23.918367,25.761246,22.680674,19.596195,16.515621,13.431144,10.350571,11.123642,11.900618,12.67369,13.450665,14.223738,14.641508,15.059279,15.477051,15.894821,16.312593,15.078801,13.841106,12.607315,11.373524,10.135828,8.956698,7.7775693,6.5984397,5.4193106,4.2362766,5.891743,7.5472097,9.202676,10.858143,12.513609,14.348679,16.183748,18.018816,19.853886,21.688955,19.498585,17.308216,15.117846,12.927476,10.737106,14.313539,17.893875,21.470308,25.04674,28.623173,24.23072,19.834364,15.438006,11.045554,6.649197,6.3993154,6.1494336,5.899552,5.64967,5.3997884,7.250475,9.101162,10.951848,12.798631,14.649317,17.429253,20.209187,22.98912,25.769054,28.548988,30.266926,31.984863,33.7028,35.42074,37.138676,36.029823,34.920975,33.81603,32.707176,31.598328,27.561176,23.524023,19.486872,15.449719,11.412568,9.136301,6.8561306,4.579864,2.3035975,0.023426414,3.5295796,7.0318284,10.534078,14.036326,17.538574,19.13938,20.73628,22.337086,23.937891,25.538694,25.585548,25.6324,25.679255,25.726107,25.776863,21.567919,17.358973,13.153932,8.944985,4.73604,4.548629,4.357313,4.165997,3.978586,3.78727,6.5086384,9.226103,11.947471,14.668839,17.386303,14.348679,11.311053,8.273428,5.2358036,2.1981785,3.6154766,5.02887,6.446168,7.859562,9.276859,8.878611,8.484266,8.089922,7.6955767,7.3012323,8.0040245,8.706817,9.405705,10.108498,10.81129,10.42085,10.034314,9.643873,9.253433,8.862993,9.073831,9.288573,9.499411,9.714153,9.924991,8.859089,7.7892823,6.7233806,5.6535745,4.5876727,5.0913405,5.5989127,6.1025805,6.606249,7.113821,8.862993,10.612165,12.361338,14.114414,15.863586,14.53609,13.208592,11.881096,10.553599,9.226103,8.320281,7.4144597,6.5086384,5.606722,4.7009,4.9546866,5.2084727,5.466163,5.7199492,5.9737353,5.5091114,5.044488,4.579864,4.11524,3.6506162,3.5881457,3.5256753,3.4632049,3.4007344,3.338264,3.1586614,2.9829633,2.803361,2.6276627,2.4480603,2.05762,1.6632754,1.2728351,0.8784905,0.48805028,0.92143893,1.3509232,1.7843118,2.2177005,2.6510892,3.057147,3.4632049,3.873167,4.279225,4.689187,4.4588275,4.2323723,4.0059166,3.775557,3.5491016,2.97125,2.3894942,1.8116426,1.2298868,0.6481308,0.5349031,0.42167544,0.30454338,0.19131571,0.07418364,1.3665408,2.6588979,3.951255,5.2436123,6.5359693,6.1181984,5.6965227,5.278752,4.8570766,4.4393053,4.435401,4.4314966,4.4314966,4.4275923,4.423688,4.7711797,5.1186714,5.466163,5.813655,6.1611466,5.02887,3.892689,2.7565079,1.6242313,0.48805028,0.5114767,0.5388075,0.5622339,0.58566034,0.61299115,0.6442264,0.6715572,0.7027924,0.7340276,0.76135844,0.94876975,1.1361811,1.3235924,1.5110037,1.698415,1.7530766,1.8038338,1.8584955,1.9092526,1.9639144,1.7921207,1.6242313,1.4524376,1.2806439,1.1127546,1.2728351,1.4329157,1.5929961,1.7530766,1.9131571,1.7804074,1.6476578,1.5149081,1.3821584,1.2494087,1.1557031,1.0659018,0.97219616,0.8784905,0.78868926,0.75354964,0.7223144,0.6910792,0.6559396,0.62470436,0.5661383,0.5036679,0.44510186,0.38653582,0.3240654,0.28892577,0.25378615,0.21864653,0.1835069,0.14836729,0.1835069,0.21474212,0.24597734,0.28111696,0.31235218,0.3474918,0.38263142,0.41777104,0.45291066,0.48805028,0.46852827,0.45291066,0.43338865,0.41777104,0.39824903,0.45681506,0.5114767,0.5661383,0.62079996,0.6754616,0.76916724,0.8589685,0.95267415,1.0463798,1.1361811,1.397776,1.6593709,1.9170616,2.1786566,2.436347,2.514435,2.592523,2.6706111,2.7486992,2.8267872,3.3031244,3.7794614,4.2557983,4.73604,5.212377,5.3256044,5.4427366,5.5559645,5.6730967,5.786324,5.571582,5.3529353,5.134289,4.9156423,4.7009,4.7009,4.7009,4.7009,4.7009,4.7009,4.7907014,4.884407,4.9781127,5.0718184,5.1616197,4.6930914,4.2284675,3.7599394,3.2914112,2.8267872,2.5027218,2.1786566,1.8584955,1.53443,1.2142692,1.9600099,2.7057507,3.455396,4.2011366,4.950782,6.168956,7.3910336,8.609207,9.8312845,11.0494585,10.370092,9.690726,9.01136,8.32809,7.648724,7.843944,8.039165,8.234385,8.429605,8.624825,9.351044,10.081166,10.807385,11.533605,12.263727,1.5617609,1.6164225,1.6710842,1.7257458,1.7843118,1.8389735,1.8819219,1.9287747,1.9717231,2.018576,2.0615244,2.135708,2.2137961,2.2879796,2.3621633,2.436347,2.5886188,2.7408905,2.893162,3.049338,3.2016098,3.3460727,3.49444,3.6428072,3.7911747,3.9356375,4.279225,4.618908,4.958591,5.298274,5.6379566,6.1103897,6.5828223,7.055255,7.5276875,8.00012,6.6960497,5.395884,4.0918136,2.7916477,1.4875772,1.2337911,0.97610056,0.7223144,0.46852827,0.21083772,0.19912452,0.1835069,0.1678893,0.15227169,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.19912452,0.19522011,0.19131571,0.1835069,0.1796025,0.1756981,0.1678893,0.16008049,0.15227169,0.14446288,0.13665408,0.12103647,0.10151446,0.08589685,0.06637484,0.05075723,0.05075723,0.05466163,0.058566034,0.058566034,0.062470436,0.093705654,0.12884527,0.16008049,0.19131571,0.22645533,0.3279698,0.42948425,0.5309987,0.63641757,0.737932,0.76916724,0.79649806,0.8277333,0.8589685,0.8862993,2.4910088,4.095718,5.704332,7.309041,8.913751,9.745388,10.577025,11.408664,12.244205,13.075843,12.689307,12.306676,11.92014,11.533605,11.150972,9.839094,8.531119,7.2192397,5.911265,4.5993857,4.5173936,4.435401,4.3534083,4.271416,4.1894236,3.9473507,3.7091823,3.4671092,3.2289407,2.9868677,3.619381,4.251894,4.884407,5.5169206,6.1494336,6.196286,6.2431393,6.2938967,6.3407493,6.387602,6.8639393,7.3441806,7.8205175,8.296855,8.773191,7.336372,5.8956475,4.454923,3.0141985,1.5734742,1.261122,0.94486535,0.62860876,0.31625658,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,1.7452679,3.4397783,5.134289,6.8287997,8.52331,7.3441806,6.165051,4.985922,3.8067923,2.6237583,3.2953155,3.9668727,4.6345253,5.3060827,5.9737353,6.1767645,6.375889,6.575013,6.774138,6.9732623,6.6413884,6.3056097,5.969831,5.6340523,5.298274,5.5871997,5.8761253,6.1611466,6.4500723,6.7389984,6.8483214,6.957645,7.066968,7.1762915,7.2856145,7.7541428,8.218767,8.683391,9.148014,9.612638,9.280765,8.94889,8.6131115,8.281238,7.9493628,8.32809,8.710721,9.089449,9.468176,9.850807,9.991365,10.131924,10.268578,10.409137,10.549695,11.408664,12.263727,13.122696,13.981665,14.836729,14.9109125,14.989,15.063184,15.137367,15.211552,15.145176,15.078801,15.008522,14.942147,14.875772,17.21451,19.553246,21.895887,24.234625,26.573362,35.26456,43.95576,52.64696,61.334255,70.02545,73.91033,77.79521,81.68009,85.56497,89.44985,81.84408,74.2344,66.628624,59.018944,51.41317,42.88986,34.36655,25.843239,17.323833,8.800523,7.871275,6.9459314,6.016684,5.0913405,4.1620927,4.40807,4.6540475,4.8961205,5.142098,5.388075,6.9459314,8.507692,10.069453,11.62731,13.189071,16.937298,20.685524,24.437654,28.18588,31.938011,28.181976,24.425941,20.67381,16.917774,13.16174,13.189071,13.216402,13.243732,13.271063,13.298394,13.075843,12.853292,12.630741,12.408191,12.185639,12.08803,11.994324,11.896713,11.799104,11.701493,17.913397,24.125301,30.337206,36.54911,42.761013,44.37353,45.98605,47.598568,49.211086,50.823605,44.100224,37.376842,30.649557,23.926178,17.198893,18.858263,20.51373,22.1731,23.828568,25.487938,22.805614,20.127193,17.448774,14.766449,12.08803,12.201257,12.31058,12.423808,12.537036,12.650263,13.005564,13.364769,13.723974,14.079274,14.438479,13.735687,13.032895,12.330102,11.62731,10.924518,9.753197,8.58578,7.4144597,6.2431393,5.0757227,7.1450562,9.21439,11.283723,13.35696,15.426293,16.816261,18.206228,19.596195,20.986162,22.37613,20.013966,17.655706,15.293544,12.935285,10.573121,15.285735,19.994444,24.707058,29.415766,34.124477,28.943335,23.766096,18.584955,13.403813,8.226576,8.1992445,8.175818,8.148487,8.125061,8.101635,9.511124,10.924518,12.337912,13.751305,15.160794,17.495626,19.826555,22.161386,24.492315,26.823244,29.23226,31.641275,34.046387,36.455402,38.86442,37.54473,36.228947,34.90926,33.593475,32.27379,28.24835,24.226816,20.201378,16.175938,12.150499,9.725866,7.3051367,4.8805027,2.4597735,0.039044023,3.408543,6.7819467,10.155351,13.528754,16.898252,18.549814,20.201378,21.849035,23.500597,25.148254,25.113115,25.08188,25.04674,25.0116,24.976461,21.056442,17.140326,13.224211,9.304191,5.388075,5.153811,4.9156423,4.6813784,4.447114,4.21285,5.930787,7.648724,9.366661,11.080693,12.798631,10.6238785,8.449126,6.2743745,4.0996222,1.9248703,3.697469,5.4700675,7.2426662,9.0152645,10.787864,10.705871,10.627783,10.545791,10.467703,10.38571,11.022127,11.6585455,12.291059,12.927476,13.563893,12.740065,11.916236,11.096312,10.272482,9.448653,9.663396,9.874233,10.088976,10.299813,10.510651,9.280765,8.046973,6.813182,5.5832953,4.349504,4.83365,5.3138914,5.7980375,6.278279,6.7624245,7.9376497,9.112875,10.2881,11.4633255,12.63855,11.576552,10.518459,9.456462,8.398369,7.336372,6.7429028,6.1494336,5.55206,4.958591,4.3612175,4.618908,4.8765984,5.134289,5.3919797,5.64967,5.0913405,4.5291066,3.970777,3.408543,2.8502135,2.9634414,3.076669,3.1859922,3.2992198,3.4124475,3.0883822,2.7682211,2.4441557,2.1239948,1.7999294,1.5539521,1.3118792,1.0659018,0.8199245,0.57394713,0.8667773,1.1596074,1.4524376,1.7452679,2.0380979,2.2567444,2.4714866,2.690133,2.9087796,3.1235218,3.2289407,3.330455,3.4319696,3.533484,3.638903,3.1039999,2.5730011,2.0380979,1.5070993,0.97610056,0.80430686,0.62860876,0.45681506,0.28502136,0.113227665,1.9561055,3.802888,5.645766,7.492548,9.339331,8.070399,6.801469,5.5364423,4.267512,2.998581,3.6037633,4.2050414,4.806319,5.4115014,6.012779,5.7668023,5.5169206,5.270943,5.0210614,4.775084,3.8848803,2.9946766,2.1044729,1.2142692,0.3240654,0.3513962,0.37482262,0.39824903,0.42557985,0.44900626,0.46852827,0.48805028,0.5114767,0.5309987,0.5505207,0.92534333,1.3001659,1.6749885,2.0498111,2.4246337,2.522244,2.619854,2.717464,2.815074,2.912684,2.6588979,2.4012074,2.1474214,1.893635,1.6359446,1.8038338,1.9678187,2.1318035,2.2957885,2.463678,2.2957885,2.1278992,1.9600099,1.7921207,1.6242313,1.4407244,1.261122,1.077615,0.8941081,0.7106012,0.6832704,0.6520352,0.62079996,0.59346914,0.5622339,0.5114767,0.45681506,0.40605783,0.3513962,0.30063897,0.27330816,0.24597734,0.21864653,0.19131571,0.1639849,0.20693332,0.24597734,0.28892577,0.3318742,0.37482262,0.41386664,0.45681506,0.4958591,0.5349031,0.57394713,0.5427119,0.5114767,0.47633708,0.44510186,0.41386664,0.4958591,0.57785153,0.659844,0.7418364,0.8238289,0.98390937,1.1400855,1.2962615,1.456342,1.6125181,1.9756275,2.3426414,2.7057507,3.0727646,3.435874,3.4983444,3.5569105,3.619381,3.677947,3.736513,4.3338866,4.93126,5.5286336,6.126007,6.7233806,6.8092775,6.8951745,6.9810715,7.0630636,7.1489606,6.9537406,6.75852,6.5633,6.36808,6.1767645,6.3134184,6.4500723,6.5867267,6.7233806,6.8639393,7.0201154,7.1762915,7.336372,7.492548,7.648724,6.930314,6.2079997,5.4895897,4.7711797,4.0488653,3.4983444,2.9439192,2.3933985,1.8389735,1.2884527,1.8506867,2.416825,2.9829633,3.5491016,4.1113358,5.153811,6.196286,7.238762,8.281238,9.323712,8.81614,8.308568,7.800996,7.2934237,6.785851,7.094299,7.3988423,7.703386,8.007929,8.312472,9.058213,9.807858,10.553599,11.303245,12.0489855,1.5617609,1.6164225,1.6671798,1.7218413,1.7725986,1.8233559,1.8741131,1.9209659,1.9678187,2.0146716,2.0615244,2.135708,2.2137961,2.2879796,2.3621633,2.436347,2.6081407,2.77603,2.9478238,3.1157131,3.2875066,3.4046388,3.521771,3.638903,3.7560349,3.873167,4.2557983,4.6384296,5.0210614,5.4036927,5.786324,6.028397,6.2743745,6.5164475,6.75852,7.000593,5.9425,4.884407,3.8263142,2.7682211,1.7140326,1.4212024,1.1322767,0.8433509,0.5544251,0.26159495,0.23035973,0.19912452,0.1639849,0.13274968,0.10151446,0.12494087,0.14836729,0.1756981,0.19912452,0.22645533,0.21083772,0.19522011,0.1796025,0.1639849,0.14836729,0.14055848,0.12884527,0.12103647,0.10932326,0.10151446,0.08589685,0.07027924,0.05466163,0.039044023,0.023426414,0.031235218,0.039044023,0.046852827,0.05466163,0.062470436,0.10932326,0.15617609,0.20693332,0.25378615,0.30063897,0.40605783,0.5153811,0.62079996,0.7301232,0.8394465,0.8784905,0.91753453,0.95657855,0.9956226,1.038571,3.1157131,5.192855,7.269997,9.347139,11.424281,12.0606985,12.693212,13.329629,13.966047,14.59856,14.055848,13.513136,12.974329,12.431617,11.888905,10.346666,8.804427,7.2582836,5.716045,4.173806,4.138666,4.1035266,4.068387,4.0332475,3.998108,3.8419318,3.6857557,3.5256753,3.3694992,3.213323,3.611572,4.0059166,4.4041657,4.802415,5.2006636,5.3177958,5.434928,5.55206,5.6691923,5.786324,6.4188375,7.0513506,7.6838636,8.316377,8.94889,7.4417906,5.9346914,4.4275923,2.920493,1.4133936,1.1283722,0.8472553,0.5661383,0.28111696,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,1.8233559,3.619381,5.4193106,7.2153354,9.01136,7.570636,6.133816,4.6930914,3.252367,1.8116426,2.697942,3.5842414,4.466636,5.3529353,6.239235,6.387602,6.5359693,6.688241,6.8366084,6.98888,6.657006,6.329036,5.997162,5.6691923,5.337318,5.4856853,5.6379566,5.786324,5.938596,6.086963,6.329036,6.571109,6.813182,7.0591593,7.3012323,7.70729,8.113348,8.52331,8.929368,9.339331,8.866898,8.3944645,7.918128,7.445695,6.9732623,7.453504,7.929841,8.406178,8.886419,9.362757,9.546264,9.725866,9.909373,10.09288,10.276386,11.147068,12.021654,12.892336,13.766922,14.637604,14.661031,14.688361,14.711788,14.739119,14.762545,14.785972,14.809398,14.828919,14.852346,14.875772,16.894348,18.916828,20.935406,22.953981,24.976461,32.855545,40.738533,48.62152,56.50451,64.3875,69.392944,74.398384,79.40383,84.40927,89.41081,81.72695,74.04308,66.35922,58.67145,50.98759,41.820053,32.652515,23.48498,14.317443,5.1499066,4.9546866,4.759466,4.564246,4.369026,4.173806,4.3612175,4.5447245,4.728231,4.9156423,5.099149,6.590631,8.086017,9.577498,11.06898,12.564366,16.113468,19.662569,23.211672,26.760773,30.31378,25.936945,21.556206,17.17937,12.802535,8.4257,9.308095,10.19049,11.072885,11.955279,12.837675,11.970898,11.10412,10.2334385,9.366661,8.499884,8.456935,8.413987,8.371038,8.32809,8.289046,16.636658,24.988174,33.33969,41.6873,50.03882,50.53858,51.038345,51.53811,52.037872,52.537636,45.599514,38.661392,31.723269,24.78905,17.850927,19.322887,20.794846,22.266806,23.738766,25.210726,22.93446,20.658192,18.378021,16.101755,13.825488,13.274967,12.724447,12.173926,11.623405,11.076789,11.373524,11.6702585,11.966993,12.263727,12.564366,12.392572,12.220779,12.05289,11.881096,11.713207,10.553599,9.393991,8.234385,7.0708723,5.911265,8.398369,10.881569,13.368673,15.851873,18.338978,19.283842,20.228708,21.173573,22.118439,23.063305,20.53325,18.003199,15.473146,12.943093,10.413041,16.254026,22.098917,27.939903,33.780888,39.62578,33.65985,27.693926,21.727999,15.765976,9.80005,9.999174,10.198298,10.401327,10.600452,10.799577,11.775677,12.751778,13.723974,14.700074,15.676175,17.562002,19.443924,21.32975,23.215576,25.101402,28.197594,31.293783,34.39388,37.49007,40.58626,39.05964,37.53302,36.006397,34.475872,32.94925,28.935526,24.925705,20.911978,16.898252,12.888432,10.319335,7.7541428,5.185046,2.6159496,0.05075723,3.2914112,6.5359693,9.776623,13.021181,16.261835,17.964155,19.662569,21.360985,23.063305,24.761719,24.644587,24.527454,24.410322,24.29319,24.17606,20.548868,16.921679,13.2905855,9.663396,6.036206,5.758993,5.477876,5.196759,4.9156423,4.6384296,5.3529353,6.067441,6.7819467,7.4964523,8.210958,6.899079,5.5871997,4.2753205,2.9634414,1.6515622,3.7794614,5.911265,8.039165,10.170968,12.298867,12.533132,12.771299,13.005564,13.239828,13.4740925,14.044135,14.610273,15.176412,15.746454,16.312593,15.059279,13.802062,12.548749,11.291532,10.0382185,10.249056,10.4637985,10.674636,10.889378,11.100216,9.702439,8.304664,6.9068875,5.5091114,4.1113358,4.572055,5.0327744,5.493494,5.9542136,6.4110284,7.012306,7.6135845,8.210958,8.812236,9.413514,8.62092,7.8283267,7.0357327,6.2431393,5.4505453,5.165524,4.8805027,4.5954814,4.31046,4.025439,4.283129,4.5447245,4.806319,5.0640097,5.3256044,4.6696653,4.0137253,3.3616903,2.7057507,2.0498111,2.338737,2.6237583,2.912684,3.2016098,3.4866312,3.018103,2.5534792,2.084951,1.6164225,1.1517987,1.0541886,0.95657855,0.8589685,0.76135844,0.6637484,0.8160201,0.96829176,1.1205635,1.2728351,1.4251068,1.4524376,1.4797685,1.5070993,1.53443,1.5617609,1.9951496,2.4285383,2.8619268,3.2914112,3.7247996,3.240654,2.7565079,2.2684577,1.7843118,1.3001659,1.0698062,0.8394465,0.60908675,0.37872702,0.14836729,2.5495746,4.942973,7.3441806,9.741484,12.138786,10.0226,7.9064145,5.794133,3.677947,1.5617609,2.7682211,3.978586,5.185046,6.3915067,7.601871,6.75852,5.9151692,5.0718184,4.2284675,3.3890212,2.7408905,2.096664,1.4524376,0.80821127,0.1639849,0.18741131,0.21083772,0.23816854,0.26159495,0.28892577,0.29673457,0.30844778,0.31625658,0.3279698,0.3357786,0.9019169,1.4641509,2.0263848,2.5886188,3.1508527,3.2914112,3.435874,3.5764325,3.7208953,3.8614538,3.521771,3.182088,2.8424048,2.5027218,2.1630387,2.330928,2.5027218,2.6706111,2.8424048,3.0141985,2.8111696,2.6081407,2.4051118,2.2020829,1.999054,1.7257458,1.456342,1.183034,0.9097257,0.63641757,0.60908675,0.58175594,0.5544251,0.5270943,0.4997635,0.45681506,0.40996224,0.3631094,0.32016098,0.27330816,0.25378615,0.23426414,0.21474212,0.19522011,0.1756981,0.22645533,0.28111696,0.3318742,0.38653582,0.43729305,0.48414588,0.5270943,0.57394713,0.61689556,0.6637484,0.61689556,0.5661383,0.5192855,0.47243267,0.42557985,0.5349031,0.6442264,0.75354964,0.8667773,0.97610056,1.1986516,1.4212024,1.6437533,1.8663043,2.0888553,2.5573835,3.0259118,3.4983444,3.9668727,4.4393053,4.478349,4.521298,4.564246,4.607195,4.650143,5.368553,6.086963,6.801469,7.519879,8.238289,8.292951,8.347612,8.402273,8.456935,8.511597,8.339804,8.16801,7.996216,7.824422,7.648724,7.9259367,8.1992445,8.476458,8.749765,9.023073,9.245625,9.468176,9.690726,9.913278,10.135828,9.163632,8.191436,7.2192397,6.2470436,5.2748475,4.493967,3.7091823,2.9283018,2.1435168,1.3626363,1.7452679,2.1278992,2.5105307,2.893162,3.2757936,4.138666,5.0054436,5.8683167,6.735094,7.601871,7.266093,6.930314,6.5945354,6.2587566,5.9268827,6.3407493,6.754616,7.168483,7.5862536,8.00012,8.769287,9.534551,10.303718,11.06898,11.838148,1.5617609,1.6125181,1.6632754,1.7140326,1.7608855,1.8116426,1.8623998,1.9131571,1.9639144,2.0107672,2.0615244,2.135708,2.2137961,2.2879796,2.3621633,2.436347,2.6237583,2.8111696,2.998581,3.1859922,3.3734035,3.4632049,3.5491016,3.638903,3.7247996,3.8106966,4.2362766,4.661856,5.087436,5.5130157,5.938596,5.950309,5.9620223,5.9737353,5.989353,6.001066,5.1889505,4.376835,3.5608149,2.7486992,1.9365835,1.6125181,1.2884527,0.96438736,0.63641757,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.10151446,0.13665408,0.1756981,0.21083772,0.24988174,0.22645533,0.19912452,0.1756981,0.14836729,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.37482262,0.48805028,0.60127795,0.7106012,0.8238289,0.93705654,0.9878138,1.038571,1.0893283,1.1361811,1.1869383,3.736513,6.2860875,8.835662,11.389141,13.938716,14.376009,14.813302,15.250595,15.687888,16.125181,15.426293,14.723501,14.024612,13.325725,12.626837,10.850334,9.073831,7.3012323,5.5247293,3.7482262,3.7638438,3.775557,3.78727,3.7989833,3.8106966,3.736513,3.6623292,3.5881457,3.513962,3.435874,3.5998588,3.7638438,3.9239242,4.087909,4.251894,4.4393053,4.6267166,4.814128,5.001539,5.1889505,5.9737353,6.7624245,7.551114,8.335898,9.124588,7.551114,5.9737353,4.4002614,2.8267872,1.2494087,0.999527,0.74964523,0.4997635,0.24988174,0.0,0.0,0.0,0.0,0.0,0.0,1.901444,3.7989833,5.700427,7.601871,9.499411,7.800996,6.098676,4.4002614,2.7018464,0.999527,2.1005683,3.2016098,4.298747,5.3997884,6.5008297,6.5984397,6.699954,6.801469,6.899079,7.000593,6.676528,6.348558,6.0244927,5.700427,5.376362,5.388075,5.3997884,5.4115014,5.423215,5.4388323,5.813655,6.1884775,6.5633,6.9381227,7.3129454,7.6643414,8.011833,8.36323,8.710721,9.062118,8.449126,7.8361354,7.223144,6.6140575,6.001066,6.575013,7.1489606,7.726812,8.300759,8.874706,9.101162,9.323712,9.550168,9.776623,9.999174,10.889378,11.775677,12.661977,13.548276,14.438479,14.411149,14.387722,14.364296,14.336966,14.313539,14.426766,14.53609,14.649317,14.762545,14.875772,16.574188,18.276506,19.974922,21.673336,23.375656,30.450434,37.52521,44.599987,51.674763,58.749542,64.87555,71.00156,77.12366,83.249664,89.37567,81.61372,73.85177,66.085915,58.32396,50.562008,40.750248,30.938484,21.122816,11.311053,1.4992905,2.0380979,2.5769055,3.1118085,3.6506162,4.1894236,4.3143644,4.4393053,4.564246,4.689187,4.814128,6.239235,7.6643414,9.089449,10.510651,11.935758,15.285735,18.635712,21.98569,25.335667,28.685644,23.68801,18.68647,13.688834,8.687295,3.6857557,5.423215,7.1606736,8.898132,10.6355915,12.373051,10.862047,9.351044,7.8361354,6.3251314,4.814128,4.825841,4.8375545,4.8492675,4.860981,4.8765984,15.363823,25.851048,36.338272,46.825497,57.31272,56.69973,56.08674,55.473747,54.860756,54.25167,47.098804,39.949844,32.800884,25.648018,18.499058,19.78751,21.075964,22.364416,23.648964,24.937418,23.063305,21.189192,19.311174,17.437061,15.562947,14.348679,13.138313,11.924045,10.71368,9.499411,9.737579,9.975748,10.213917,10.44818,10.686349,11.0494585,11.412568,11.775677,12.138786,12.501896,11.350098,10.198298,9.050405,7.898606,6.7507114,9.651682,12.548749,15.449719,18.35069,21.251661,21.751425,22.251188,22.750952,23.250715,23.750479,21.048632,18.35069,15.648844,12.950902,10.249056,17.226223,24.199486,31.176653,38.149914,45.123177,38.37637,31.625658,24.874947,18.124235,11.373524,11.799104,12.224684,12.650263,13.075843,13.501423,14.036326,14.575133,15.113941,15.648844,16.187653,17.624472,19.061293,20.498112,21.938837,23.375656,27.162926,30.950197,34.73747,38.52474,42.312008,40.574547,38.83709,37.09963,35.36217,33.624714,29.626604,25.624592,21.626484,17.624472,13.626364,10.912805,8.1992445,5.4856853,2.77603,0.062470436,3.174279,6.2860875,9.4018,12.513609,15.625418,17.37459,19.123762,20.876839,22.62601,24.375183,24.17606,23.976934,23.773905,23.574781,23.375656,20.037392,16.69913,13.360865,10.0265045,6.688241,6.364176,6.036206,5.7121406,5.388075,5.0640097,4.775084,4.4861584,4.2011366,3.912211,3.6232853,3.174279,2.7252727,2.2762666,1.8233559,1.3743496,3.8614538,6.348558,8.835662,11.326671,13.813775,14.364296,14.9109125,15.461433,16.011953,16.562475,17.062239,17.562002,18.061766,18.56153,19.061293,17.37459,15.687888,14.001186,12.31058,10.6238785,10.838621,11.0494585,11.2642,11.475039,11.685876,10.124115,8.562354,7.000593,5.4388323,3.873167,4.3143644,4.7516575,5.1889505,5.6262436,6.0635366,6.086963,6.114294,6.13772,6.1611466,6.1884775,5.661383,5.138193,4.6110992,4.087909,3.5608149,3.5881457,3.611572,3.638903,3.6623292,3.6857557,3.951255,4.21285,4.474445,4.73604,5.001539,4.251894,3.4983444,2.7486992,1.999054,1.2494087,1.7140326,2.174752,2.639376,3.1000953,3.5608149,2.951728,2.338737,1.7257458,1.1127546,0.4997635,0.5505207,0.60127795,0.6481308,0.698888,0.74964523,0.76135844,0.77307165,0.78868926,0.80040246,0.81211567,0.6481308,0.48805028,0.3240654,0.1639849,0.0,0.76135844,1.5266213,2.2879796,3.049338,3.8106966,3.3734035,2.9361105,2.4988174,2.0615244,1.6242313,1.33921,1.0502841,0.76135844,0.47633708,0.18741131,3.1391394,6.086963,9.0386915,11.986515,14.938243,11.974802,9.01136,6.0518236,3.0883822,0.12494087,1.9365835,3.7482262,5.563773,7.375416,9.187058,7.7502384,6.3134184,4.8765984,3.435874,1.999054,1.6008049,1.1986516,0.80040246,0.39824903,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.8745861,1.6242313,2.3738766,3.1235218,3.873167,4.0605783,4.251894,4.4393053,4.6267166,4.814128,4.388548,3.9629683,3.5373883,3.1118085,2.6862288,2.8619268,3.0376248,3.213323,3.3890212,3.5608149,3.3265507,3.0883822,2.8502135,2.612045,2.3738766,2.0107672,1.6515622,1.2884527,0.92534333,0.5622339,0.5388075,0.5114767,0.48805028,0.46071947,0.43729305,0.39824903,0.3631094,0.3240654,0.28892577,0.24988174,0.23816854,0.22645533,0.21083772,0.19912452,0.18741131,0.24988174,0.31235218,0.37482262,0.43729305,0.4997635,0.5505207,0.60127795,0.6481308,0.698888,0.74964523,0.6871748,0.62470436,0.5622339,0.4997635,0.43729305,0.57394713,0.7106012,0.8511597,0.9878138,1.1244678,1.4133936,1.698415,1.9873407,2.2762666,2.5612879,3.1391394,3.7130866,4.2870336,4.860981,5.4388323,5.462259,5.4856853,5.5130157,5.5364423,5.563773,6.3993154,7.238762,8.074304,8.913751,9.749292,9.776623,9.80005,9.823476,9.850807,9.874233,9.725866,9.573594,9.425227,9.276859,9.124588,9.538455,9.948417,10.362284,10.77615,11.186112,11.475039,11.763964,12.0489855,12.337912,12.626837,11.400854,10.174872,8.94889,7.726812,6.5008297,5.4856853,4.474445,3.4632049,2.4519646,1.43682,1.6359446,1.8389735,2.0380979,2.2372224,2.436347,3.1235218,3.8106966,4.5017757,5.1889505,5.8761253,5.7121406,5.548156,5.388075,5.22409,5.0640097,5.5871997,6.114294,6.6374836,7.1606736,7.687768,8.476458,9.261242,10.049932,10.838621,11.623405,1.5266213,1.5773785,1.6281357,1.6827974,1.7335546,1.7882162,1.8389735,1.893635,1.9443923,1.999054,2.0498111,2.1278992,2.2059872,2.2840753,2.358259,2.436347,2.6237583,2.8111696,2.998581,3.1859922,3.3734035,3.4788225,3.5842414,3.68966,3.795079,3.900498,4.283129,4.6696653,5.056201,5.4388323,5.825368,5.7707067,5.7199492,5.6691923,5.6145306,5.563773,4.841459,4.123049,3.4007344,2.6823244,1.9639144,1.6281357,1.2962615,0.96438736,0.63251317,0.30063897,0.25378615,0.20693332,0.15617609,0.10932326,0.062470436,0.09761006,0.13274968,0.1678893,0.20302892,0.23816854,0.21474212,0.19131571,0.1717937,0.14836729,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.06637484,0.06637484,0.07027924,0.07418364,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.13665408,0.19131571,0.24207294,0.29673457,0.3474918,0.39824903,0.58566034,0.76916724,0.95657855,1.1400855,1.3235924,1.5578566,1.7882162,2.0224805,2.2567444,2.4871042,4.5681505,6.6531014,8.734148,10.819098,12.900145,13.583415,14.27059,14.95386,15.641035,16.324306,15.570756,14.821111,14.067561,13.314012,12.564366,10.924518,9.288573,7.648724,6.012779,4.376835,4.165997,3.959064,3.7521305,3.5451972,3.338264,3.3070288,3.2757936,3.2484627,3.2172275,3.1859922,3.3460727,3.506153,3.6662338,3.8263142,3.9863946,4.3026514,4.618908,4.93126,5.2475166,5.563773,6.250948,6.942027,7.633106,8.324185,9.01136,7.5003567,5.989353,4.474445,2.9634414,1.4485333,1.2064602,0.96438736,0.7223144,0.48024148,0.23816854,0.21474212,0.19131571,0.1717937,0.14836729,0.12494087,1.620327,3.1157131,4.6110992,6.1064854,7.601871,6.4383593,5.278752,4.1191444,2.959537,1.7999294,2.494913,3.1898966,3.8848803,4.579864,5.2748475,5.364649,5.45445,5.5442514,5.6340523,5.7238536,5.6535745,5.579391,5.5091114,5.434928,5.3607445,5.466163,5.571582,5.677001,5.7824197,5.8878384,6.1494336,6.407124,6.6687193,6.9264097,7.1880045,7.445695,7.70729,7.968885,8.226576,8.488171,8.101635,7.7111945,7.3246584,6.9381227,6.551587,7.2075267,7.8634663,8.52331,9.17925,9.839094,9.975748,10.116306,10.256865,10.397423,10.537982,11.361811,12.181735,13.005564,13.829392,14.649317,14.914817,15.180316,15.445815,15.711315,15.976814,16.894348,17.811884,18.729418,19.646952,20.560583,22.40346,24.242434,26.081408,27.924286,29.763258,35.53787,41.31248,47.08709,52.861702,58.636314,63.286457,67.93269,72.57893,77.22908,81.87531,74.79273,67.710144,60.62756,53.54497,46.462387,37.58768,28.712975,19.838268,10.963562,2.0888553,2.893162,3.7013733,4.5095844,5.3177958,6.126007,6.211904,6.3017054,6.387602,6.473499,6.5633,7.2934237,8.023546,8.75367,9.483793,10.213917,13.700547,17.18718,20.67381,24.164345,27.650976,22.914936,18.178898,13.446761,8.710721,3.9746814,5.4310236,6.883461,8.339804,9.796145,11.248583,10.249056,9.245625,8.242193,7.238762,6.239235,5.938596,5.6379566,5.337318,5.036679,4.73604,14.313539,23.891037,33.468536,43.046036,52.623535,53.40051,54.17358,54.950558,55.72363,56.500607,49.394592,42.28858,35.186474,28.080462,20.97445,21.962263,22.950077,23.937891,24.925705,25.913517,23.891037,21.868557,19.846077,17.823597,15.801116,14.376009,12.950902,11.525795,10.100689,8.675582,9.101162,9.526741,9.948417,10.373997,10.799577,10.955752,11.111929,11.2642,11.420377,11.576552,10.58093,9.589212,8.597494,7.605776,6.6140575,8.898132,11.182208,13.466284,15.754263,18.038338,19.022247,20.006157,20.99397,21.97788,22.96179,20.712854,18.463919,16.211079,13.962143,11.713207,17.226223,22.739239,28.24835,33.761368,39.274384,34.046387,28.81449,23.586494,18.354595,13.1266,13.438952,13.755209,14.0714655,14.383818,14.700074,15.21936,15.734741,16.254026,16.769407,17.288692,18.346786,19.400974,20.459068,21.51716,22.575254,25.936945,29.29473,32.65642,36.014206,39.375896,37.689194,35.99859,34.311886,32.625187,30.938484,27.393286,23.84809,20.30289,16.757694,13.212498,10.865952,8.519405,6.168956,3.8224099,1.475864,4.5564375,7.633106,10.71368,13.794253,16.874826,18.307743,19.740658,21.173573,22.60649,24.039404,23.79733,23.559164,23.317091,23.078922,22.83685,19.619621,16.402393,13.185166,9.967939,6.7507114,6.3836975,6.016684,5.645766,5.278752,4.911738,4.630621,4.3534083,4.0722914,3.7911747,3.513962,3.2016098,2.8892577,2.5769055,2.260649,1.9482968,5.1186714,8.285142,11.4516115,14.621986,17.788456,18.046146,18.303837,18.56153,18.81922,19.07691,19.073006,19.069101,19.069101,19.065197,19.061293,17.351164,15.637131,13.923099,12.212971,10.498938,10.61607,10.733202,10.8542385,10.971371,11.088503,9.80005,8.511597,7.223144,5.938596,4.650143,5.0483923,5.4505453,5.8487945,6.250948,6.649197,6.407124,6.165051,5.9229784,5.6809053,5.4388323,5.0522966,4.6657605,4.283129,3.8965936,3.513962,3.4983444,3.4827268,3.4671092,3.4514916,3.435874,3.7013733,3.9629683,4.224563,4.4861584,4.7516575,4.009821,3.2718892,2.5300527,1.7882162,1.0502841,1.4212024,1.796025,2.1669433,2.541766,2.912684,2.4129205,1.9131571,1.4133936,0.9136301,0.41386664,0.5153811,0.61689556,0.71841,0.8238289,0.92534333,0.8784905,0.8355421,0.78868926,0.74574083,0.698888,0.5583295,0.42167544,0.28111696,0.14055848,0.0,0.62079996,1.2455044,1.8663043,2.4910088,3.1118085,2.7526035,2.3933985,2.0341935,1.6710842,1.3118792,1.0854238,0.8589685,0.62860876,0.40215343,0.1756981,2.5808098,4.985922,7.3910336,9.796145,12.201257,9.784432,7.3715115,4.9546866,2.541766,0.12494087,1.6008049,3.076669,4.548629,6.0244927,7.5003567,6.379793,5.2592297,4.138666,3.018103,1.901444,1.5266213,1.1557031,0.78088045,0.40996224,0.039044023,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.1678893,0.1717937,0.1756981,0.1835069,0.18741131,0.79259366,1.397776,2.0029583,2.6081407,3.213323,3.357786,3.5022488,3.6467118,3.7911747,3.9356375,3.5998588,3.2640803,2.9243972,2.5886188,2.2489357,2.6940374,3.135235,3.5764325,4.0215344,4.462732,4.251894,4.041056,3.8341231,3.6232853,3.4124475,2.87364,2.338737,1.7999294,1.261122,0.7262188,0.6832704,0.64032197,0.59737355,0.5544251,0.5114767,0.45681506,0.40215343,0.3474918,0.29283017,0.23816854,0.24207294,0.24597734,0.25378615,0.25769055,0.26159495,0.31625658,0.3709182,0.42557985,0.48414588,0.5388075,0.5622339,0.58566034,0.61299115,0.63641757,0.6637484,0.7418364,0.8160201,0.8941081,0.97219616,1.0502841,1.1205635,1.1947471,1.2689307,1.33921,1.4133936,1.7686942,2.1239948,2.4792955,2.8306916,3.1859922,3.8497405,4.513489,5.173333,5.8370814,6.5008297,6.4891167,6.473499,6.461786,6.4500723,6.4383593,7.250475,8.062591,8.874706,9.686822,10.498938,10.729298,10.955752,11.182208,11.408664,11.639023,11.45942,11.283723,11.10412,10.928422,10.748819,10.783959,10.819098,10.8542385,10.889378,10.924518,10.986988,11.0494585,11.111929,11.174399,11.23687,10.401327,9.565785,8.734148,7.898606,7.0630636,6.2314262,5.395884,4.564246,3.7326086,2.900971,3.0024853,3.1039999,3.2094188,3.310933,3.4124475,3.7833657,4.154284,4.521298,4.892216,5.263134,5.1225758,4.9820175,4.841459,4.7009,4.564246,5.1030536,5.6418614,6.180669,6.7233806,7.262188,8.03526,8.8083315,9.581403,10.350571,11.123642,1.4875772,1.542239,1.5969005,1.6515622,1.7062237,1.7608855,1.815547,1.8741131,1.9287747,1.9834363,2.0380979,2.1161861,2.1981785,2.2762666,2.358259,2.436347,2.6237583,2.8111696,2.998581,3.1859922,3.3734035,3.4983444,3.619381,3.7443218,3.8653584,3.9863946,4.3338866,4.677474,5.0210614,5.368553,5.7121406,5.5950084,5.477876,5.3607445,5.2436123,5.12648,4.4978714,3.8692627,3.240654,2.6159496,1.9873407,1.6476578,1.3079748,0.96829176,0.62860876,0.28892577,0.24207294,0.19912452,0.15227169,0.10932326,0.062470436,0.093705654,0.12884527,0.16008049,0.19131571,0.22645533,0.20693332,0.1835069,0.1639849,0.14446288,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.078088045,0.09761006,0.113227665,0.13274968,0.14836729,0.1639849,0.1756981,0.18741131,0.19912452,0.21083772,0.25378615,0.29673457,0.339683,0.38263142,0.42557985,0.6832704,0.94096094,1.1986516,1.456342,1.7140326,2.1278992,2.541766,2.9556324,3.3734035,3.78727,5.4036927,7.016211,8.632633,10.249056,11.861574,12.794726,13.727879,14.661031,15.594183,16.52343,15.719124,14.914817,14.11051,13.306203,12.501896,10.998701,9.499411,8.00012,6.5008297,5.001539,4.572055,4.1464753,3.716991,3.2914112,2.8619268,2.8775444,2.893162,2.9087796,2.9243972,2.9361105,3.096191,3.252367,3.408543,3.5686235,3.7247996,4.165997,4.6110992,5.0522966,5.493494,5.938596,6.5281606,7.1216297,7.715099,8.308568,8.898132,7.4495993,6.001066,4.548629,3.1000953,1.6515622,1.4133936,1.1791295,0.94486535,0.7106012,0.47633708,0.42948425,0.38653582,0.339683,0.29673457,0.24988174,1.33921,2.4285383,3.521771,4.6110992,5.700427,5.0796275,4.4588275,3.8380275,3.2211318,2.6003318,2.8892577,3.1781836,3.4710135,3.7599394,4.0488653,4.1308575,4.2089458,4.290938,4.369026,4.4510183,4.630621,4.8102236,4.989826,5.169429,5.349031,5.548156,5.743376,5.9425,6.141625,6.336845,6.481308,6.6257706,6.774138,6.918601,7.0630636,7.230953,7.4027467,7.570636,7.7424297,7.914223,7.7502384,7.5862536,7.426173,7.262188,7.098203,7.8400397,8.581876,9.319808,10.061645,10.799577,10.8542385,10.9089,10.963562,11.018223,11.076789,11.834243,12.591698,13.349152,14.106606,14.864059,15.418485,15.97291,16.527334,17.08176,17.636185,19.36193,21.083773,22.805614,24.527454,26.249296,28.228828,30.20836,32.191795,34.17133,36.15086,40.625305,45.09975,49.574196,54.04864,58.523087,61.69346,64.86384,68.03421,71.20458,74.37496,67.97174,61.56852,55.169205,48.765984,42.362766,34.425114,26.487465,18.549814,10.612165,2.6745155,3.7521305,4.829746,5.9073606,6.984976,8.062591,8.113348,8.164105,8.210958,8.261715,8.312472,8.347612,8.382751,8.4178915,8.453031,8.488171,12.111456,15.738646,19.36193,22.98912,26.612406,22.141865,17.671324,13.200784,8.734148,4.263607,5.434928,6.606249,7.7814736,8.952794,10.124115,9.63216,9.140205,8.648251,8.156297,7.6643414,7.0513506,6.4383593,5.825368,5.212377,4.5993857,13.2671585,21.934933,30.602705,39.270477,47.93825,50.101288,52.264328,54.423462,56.586502,58.749542,51.69038,44.63122,37.568157,30.508999,23.44984,24.137014,24.82419,25.511364,26.19854,26.885714,24.718771,22.547922,20.377075,18.206228,16.039284,14.399435,12.763491,11.123642,9.487698,7.8517528,8.460839,9.073831,9.686822,10.299813,10.912805,10.858143,10.807385,10.756628,10.701966,10.651209,9.815667,8.980125,8.144583,7.309041,6.473499,8.144583,9.815667,11.486752,13.153932,14.825015,16.296974,17.76503,19.233086,20.705046,22.1731,20.37317,18.573242,16.773312,14.973383,13.173453,17.226223,21.275087,25.323954,29.376722,33.425587,29.716406,26.003319,22.294136,18.584955,14.875772,15.078801,15.285735,15.488764,15.695697,15.8987255,16.398489,16.894348,17.394112,17.88997,18.38583,19.065197,19.740658,20.420023,21.09939,21.77485,24.707058,27.639263,30.57147,33.503677,36.435883,34.79994,33.163994,31.524143,29.888199,28.24835,25.159967,22.071587,18.9793,15.890917,12.798631,10.819098,8.835662,6.852226,4.8687897,2.8892577,5.9346914,8.98403,12.029464,15.078801,18.124235,19.240894,20.35365,21.470308,22.586967,23.699722,23.418604,23.141392,22.860275,22.579159,22.301945,19.20185,16.10566,13.005564,9.909373,6.813182,6.4032197,5.9932575,5.5832953,5.173333,4.7633705,4.4900627,4.2167544,3.9434462,3.6740425,3.4007344,3.2250361,3.049338,2.87364,2.7018464,2.5261483,6.3719845,10.221725,14.067561,17.913397,21.763138,21.727999,21.69286,21.657719,21.62258,21.58744,21.083773,20.5762,20.072533,19.568865,19.061293,17.323833,15.586374,13.848915,12.111456,10.373997,10.397423,10.42085,10.444276,10.4637985,10.487225,9.475985,8.460839,7.4495993,6.4383593,5.423215,5.786324,6.1494336,6.5125427,6.8756523,7.238762,6.727285,6.2158084,5.708236,5.196759,4.689187,4.4432096,4.1972322,3.951255,3.7091823,3.4632049,3.408543,3.3538816,3.2992198,3.240654,3.1859922,3.4514916,3.7130866,3.9746814,4.2362766,4.5017757,3.7716527,3.0415294,2.3114061,1.5812829,0.8511597,1.1322767,1.4133936,1.698415,1.979532,2.260649,1.8741131,1.4875772,1.1010414,0.7106012,0.3240654,0.48024148,0.63641757,0.78868926,0.94486535,1.1010414,0.9956226,0.8941081,0.79259366,0.6910792,0.58566034,0.46852827,0.3513962,0.23426414,0.11713207,0.0,0.48414588,0.96438736,1.4485333,1.9287747,2.4129205,2.1318035,1.8467822,1.5656652,1.2806439,0.999527,0.8316377,0.6637484,0.4958591,0.3318742,0.1639849,2.0224805,3.8809757,5.743376,7.601871,9.464272,7.5940623,5.727758,3.8614538,1.9912452,0.12494087,1.261122,2.4012074,3.5373883,4.6735697,5.813655,5.009348,4.2089458,3.4046388,2.6042364,1.7999294,1.456342,1.1088502,0.76526284,0.42167544,0.07418364,0.10151446,0.12494087,0.14836729,0.1756981,0.19912452,0.21083772,0.21864653,0.23035973,0.23816854,0.24988174,0.7106012,1.1713207,1.6281357,2.0888553,2.5495746,2.6510892,2.7565079,2.8580225,2.959537,3.0610514,2.8111696,2.5612879,2.3114061,2.0615244,1.8116426,2.522244,3.232845,3.9434462,4.6540475,5.3607445,5.181142,4.997635,4.814128,4.630621,4.4510183,3.736513,3.0259118,2.3114061,1.6008049,0.8862993,0.8277333,0.76916724,0.7066968,0.6481308,0.58566034,0.5153811,0.44119745,0.3709182,0.29673457,0.22645533,0.24597734,0.26940376,0.29283017,0.31625658,0.3357786,0.38653582,0.43338865,0.48024148,0.5270943,0.57394713,0.57394713,0.57394713,0.57394713,0.57394713,0.57394713,0.79259366,1.0112402,1.2259823,1.4446288,1.6632754,1.6710842,1.678893,1.6867018,1.6906061,1.698415,2.1239948,2.5456703,2.9673457,3.3890212,3.8106966,4.564246,5.3138914,6.0635366,6.813182,7.562827,7.5120697,7.461313,7.4105554,7.363703,7.3129454,8.101635,8.886419,9.675109,10.4637985,11.248583,11.681972,12.111456,12.54094,12.970425,13.399908,13.196879,12.989946,12.786918,12.579984,12.376955,12.033368,11.68978,11.346193,11.00651,10.662923,10.498938,10.338858,10.174872,10.010887,9.850807,9.405705,8.960603,8.515501,8.070399,7.6252975,6.9732623,6.321227,5.6691923,5.0132523,4.3612175,4.369026,4.3729305,4.376835,4.380739,4.388548,4.4393053,4.493967,4.5447245,4.5993857,4.650143,4.533011,4.415879,4.298747,4.181615,4.0605783,4.618908,5.173333,5.727758,6.282183,6.8366084,7.5940623,8.351517,9.108971,9.866425,10.6238785,1.4485333,1.5070993,1.5656652,1.6242313,1.678893,1.737459,1.796025,1.8506867,1.9092526,1.9678187,2.0263848,2.1083772,2.1903696,2.2723622,2.3543546,2.436347,2.6237583,2.8111696,2.998581,3.1859922,3.3734035,3.513962,3.6545205,3.795079,3.9356375,4.0761957,4.380739,4.6852827,4.989826,5.2943697,5.5989127,5.4193106,5.2358036,5.0522966,4.8687897,4.689187,4.154284,3.619381,3.0805733,2.5456703,2.0107672,1.6632754,1.3157835,0.96829176,0.62079996,0.27330816,0.23426414,0.19131571,0.14836729,0.10541886,0.062470436,0.093705654,0.12103647,0.15227169,0.1835069,0.21083772,0.19522011,0.1756981,0.16008049,0.14055848,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.093705654,0.12884527,0.16008049,0.19131571,0.22645533,0.23816854,0.24988174,0.26159495,0.27330816,0.28892577,0.32016098,0.3513962,0.38653582,0.41777104,0.44900626,0.78088045,1.1088502,1.4407244,1.7686942,2.1005683,2.697942,3.2953155,3.892689,4.4900627,5.087436,6.2353306,7.3832245,8.531119,9.679013,10.826907,12.006037,13.185166,14.364296,15.543426,16.72646,15.867491,15.008522,14.153459,13.29449,12.439425,11.076789,9.714153,8.351517,6.98888,5.6262436,4.9781127,4.3299823,3.6818514,3.0337205,2.3855898,2.4480603,2.5066261,2.5690966,2.6276627,2.6862288,2.8424048,2.998581,3.1508527,3.3070288,3.4632049,4.0332475,4.60329,5.173333,5.743376,6.3134184,6.8092775,7.3012323,7.7970915,8.292951,8.78881,7.3988423,6.012779,4.6267166,3.2367494,1.8506867,1.6242313,1.3938715,1.1674163,0.94096094,0.7106012,0.6442264,0.57785153,0.5114767,0.44119745,0.37482262,1.0580931,1.7452679,2.4285383,3.1157131,3.7989833,3.7208953,3.638903,3.5608149,3.4788225,3.4007344,3.2836022,3.1703746,3.0532427,2.9400148,2.8267872,2.893162,2.9634414,3.0337205,3.1039999,3.174279,3.6076677,4.041056,4.474445,4.903929,5.337318,5.6262436,5.919074,6.2079997,6.4969254,6.785851,6.817086,6.8483214,6.8756523,6.9068875,6.9381227,7.016211,7.098203,7.1762915,7.2582836,7.336372,7.3988423,7.461313,7.523783,7.5862536,7.648724,8.472553,9.296382,10.116306,10.940135,11.763964,11.732729,11.701493,11.674163,11.642927,11.611692,12.306676,12.997755,13.688834,14.383818,15.074897,15.918248,16.765503,17.608854,18.45611,19.29946,21.82561,24.355661,26.88181,29.411861,31.938011,34.0581,36.178192,38.298283,40.418373,42.538464,45.71274,48.88702,52.0613,55.239483,58.41376,60.10437,61.798878,63.489487,65.184,66.8746,61.15075,55.430798,49.706944,43.983093,38.26314,31.262548,24.261955,17.261362,10.260769,3.2640803,4.6110992,5.958118,7.3051367,8.652155,9.999174,10.010887,10.0265045,10.0382185,10.049932,10.061645,9.4018,8.741957,8.082112,7.422269,6.7624245,10.526268,14.286208,18.05005,21.813896,25.573835,21.368793,17.163752,12.958711,8.75367,4.548629,5.4388323,6.329036,7.2192397,8.109444,8.999647,9.019169,9.034787,9.054309,9.069926,9.089449,8.164105,7.238762,6.3134184,5.388075,4.462732,12.220779,19.978827,27.736874,35.491016,43.249065,46.798164,50.351173,53.900272,57.449375,60.998478,53.98617,46.96996,39.953747,32.94144,25.925232,26.311768,26.698303,27.088743,27.475279,27.861814,25.546503,23.22729,20.908073,18.592764,16.273548,14.426766,12.576079,10.725393,8.874706,7.0240197,7.824422,8.624825,9.425227,10.22563,11.0260315,10.764437,10.506746,10.2451515,9.983557,9.725866,9.0465,8.371038,7.6916723,7.016211,6.336845,7.3910336,8.449126,9.503315,10.557504,11.611692,13.567798,15.523903,17.476105,19.43221,21.388315,20.037392,18.68647,17.335546,15.988527,14.637604,17.226223,19.810938,22.399555,24.988174,27.576794,25.386423,23.196054,21.005684,18.815315,16.624945,16.71865,16.816261,16.909966,17.003672,17.101282,17.57762,18.053955,18.534197,19.010534,19.486872,19.783606,20.084246,20.38098,20.677715,20.97445,23.481075,25.983797,28.490423,30.993145,33.49977,31.910679,30.325493,28.7364,27.151213,25.562122,22.926651,20.291178,17.655706,15.024139,12.388668,10.768341,9.151918,7.535496,5.919074,4.298747,7.3168497,10.331048,13.345247,16.359446,19.373644,20.174046,20.970545,21.767042,22.563541,23.363943,23.043781,22.723621,22.40346,22.0833,21.763138,18.784079,15.808925,12.829865,9.850807,6.8756523,6.422742,5.969831,5.5169206,5.0640097,4.6110992,4.3455997,4.084005,3.8185053,3.5530062,3.2875066,3.2484627,3.213323,3.174279,3.1391394,3.1000953,7.629202,12.154405,16.683512,21.208714,25.73782,25.40985,25.08188,24.75391,24.425941,24.101875,23.090635,22.0833,21.075964,20.068628,19.061293,17.300406,15.535617,13.774731,12.013845,10.249056,10.178777,10.104593,10.034314,9.96013,9.885946,9.148014,8.413987,7.676055,6.9381227,6.2001905,6.524256,6.8483214,7.1762915,7.5003567,7.824422,7.0474463,6.27047,5.493494,4.716518,3.9356375,3.8341231,3.7287042,3.6232853,3.5178664,3.4124475,3.3187418,3.2211318,3.1274261,3.0337205,2.9361105,3.2016098,3.4632049,3.7247996,3.9863946,4.251894,3.5295796,2.8111696,2.0888553,1.3704453,0.6481308,0.8433509,1.0346665,1.2259823,1.4212024,1.6125181,1.33921,1.0619974,0.78868926,0.5114767,0.23816854,0.44510186,0.6520352,0.8589685,1.0659018,1.2767396,1.116659,0.95657855,0.79649806,0.63641757,0.47633708,0.37872702,0.28502136,0.19131571,0.093705654,0.0,0.3435874,0.6832704,1.0268579,1.3704453,1.7140326,1.5070993,1.3040704,1.097137,0.8941081,0.6871748,0.58175594,0.47243267,0.3631094,0.25769055,0.14836729,1.4641509,2.7799344,4.095718,5.4115014,6.7233806,5.4036927,4.084005,2.7643168,1.4446288,0.12494087,0.92534333,1.7257458,2.5261483,3.3265507,4.123049,3.638903,3.154757,2.6706111,2.1864653,1.698415,1.3821584,1.0659018,0.74574083,0.42948425,0.113227665,0.13665408,0.1639849,0.18741131,0.21083772,0.23816854,0.25378615,0.26940376,0.28111696,0.29673457,0.31235218,0.62860876,0.94096094,1.2572175,1.5734742,1.8858263,1.9482968,2.0068626,2.069333,2.1278992,2.1864653,2.0263848,1.8623998,1.698415,1.5383345,1.3743496,2.3543546,3.330455,4.3065557,5.2865605,6.262661,6.1064854,5.9542136,5.7980375,5.6418614,5.4856853,4.5993857,3.7130866,2.8267872,1.9365835,1.0502841,0.97219616,0.8941081,0.8160201,0.7418364,0.6637484,0.57394713,0.48414588,0.39434463,0.30063897,0.21083772,0.25378615,0.29283017,0.3318742,0.3709182,0.41386664,0.45291066,0.49195468,0.5309987,0.57394713,0.61299115,0.58566034,0.5622339,0.5388075,0.5114767,0.48805028,0.8433509,1.2025559,1.5617609,1.9170616,2.2762666,2.2177005,2.1591344,2.1005683,2.0459068,1.9873407,2.4792955,2.9673457,3.4593005,3.9473507,4.4393053,5.2748475,6.114294,6.949836,7.7892823,8.624825,8.538928,8.449126,8.36323,8.273428,8.187531,8.94889,9.714153,10.475512,11.23687,11.998228,12.630741,13.263254,13.895767,14.528281,15.160794,14.930434,14.69617,14.465811,14.231546,14.001186,13.2788725,12.560462,11.838148,11.119738,10.401327,10.010887,9.6243515,9.237816,8.85128,8.460839,8.406178,8.351517,8.296855,8.242193,8.187531,7.715099,7.2426662,6.7702336,6.297801,5.825368,5.7316628,5.6418614,5.548156,5.45445,5.3607445,5.099149,4.83365,4.5681505,4.3026514,4.037152,3.9434462,3.8458362,3.7521305,3.6584249,3.5608149,4.1308575,4.7009,5.270943,5.840986,6.4110284,7.1567693,7.898606,8.640442,9.382278,10.124115,1.4133936,1.4719596,1.53443,1.5929961,1.6515622,1.7140326,1.7725986,1.8311646,1.893635,1.9522011,2.0107672,2.096664,2.182561,2.2684577,2.3543546,2.436347,2.6237583,2.8111696,2.998581,3.1859922,3.3734035,3.533484,3.68966,3.8458362,4.0059166,4.1620927,4.4275923,4.6930914,4.958591,5.22409,5.4856853,5.239708,4.9937305,4.743849,4.4978714,4.251894,3.8067923,3.3655949,2.9243972,2.4792955,2.0380979,1.6827974,1.3274968,0.97219616,0.61689556,0.26159495,0.22255093,0.1835069,0.14055848,0.10151446,0.062470436,0.08980125,0.11713207,0.14446288,0.1717937,0.19912452,0.1835069,0.1717937,0.15617609,0.14055848,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.10932326,0.15617609,0.20693332,0.25378615,0.30063897,0.31235218,0.3240654,0.3357786,0.3513962,0.3631094,0.38653582,0.40605783,0.42948425,0.45291066,0.47633708,0.8784905,1.2806439,1.6827974,2.084951,2.4871042,3.2679846,4.0488653,4.825841,5.606722,6.387602,7.066968,7.746334,8.4257,9.108971,9.788337,11.213444,12.642454,14.0714655,15.4965725,16.925583,16.015858,15.1061325,14.196406,13.286681,12.373051,11.150972,9.924991,8.699008,7.47693,6.250948,5.3841705,4.513489,3.6467118,2.7799344,1.9131571,2.018576,2.1239948,2.2294137,2.330928,2.436347,2.5886188,2.7408905,2.893162,3.049338,3.2016098,3.8965936,4.5954814,5.2943697,5.989353,6.688241,7.08649,7.480835,7.8790836,8.277332,8.675582,7.348085,6.0244927,4.7009,3.3734035,2.0498111,1.8311646,1.6086137,1.3899672,1.1713207,0.94876975,0.8589685,0.76916724,0.679366,0.58956474,0.4997635,0.78088045,1.0580931,1.33921,1.620327,1.901444,2.358259,2.8189783,3.279698,3.7404175,4.2011366,3.6818514,3.1586614,2.639376,2.1200905,1.6008049,1.6593709,1.7218413,1.7804074,1.8389735,1.901444,2.5847144,3.2718892,3.9551594,4.6384296,5.3256044,5.708236,6.0908675,6.473499,6.8561306,7.238762,7.152865,7.066968,6.9810715,6.899079,6.813182,6.801469,6.79366,6.7819467,6.774138,6.7624245,7.0513506,7.336372,7.6252975,7.914223,8.1992445,9.105066,10.010887,10.916709,11.818625,12.724447,12.611219,12.494087,12.380859,12.263727,12.150499,12.779109,13.403813,14.032422,14.661031,15.285735,16.421915,17.558098,18.694279,19.826555,20.962736,24.29319,27.62755,30.96191,34.292366,37.626724,39.88347,42.14412,44.404766,46.665417,48.926064,50.80018,52.67429,54.548405,56.426422,58.300533,58.515278,58.73002,58.94476,59.159504,59.374245,54.33366,49.289173,44.248592,39.2041,34.16352,28.099983,22.036446,15.97291,9.913278,3.8497405,5.466163,7.08649,8.702912,10.319335,11.935758,11.912332,11.888905,11.861574,11.838148,11.810817,10.455989,9.101162,7.746334,6.3915067,5.036679,8.937177,12.837675,16.738173,20.63867,24.539167,20.595722,16.65618,12.716639,8.777096,4.8375545,5.446641,6.0518236,6.66091,7.266093,7.8751793,8.402273,8.929368,9.456462,9.983557,10.510651,9.276859,8.039165,6.801469,5.563773,4.3260775,11.170495,18.018816,24.867138,31.71546,38.56378,43.498947,48.438015,53.377083,58.31225,63.251316,56.28196,49.308697,42.339336,35.36998,28.400621,28.486519,28.57632,28.662216,28.748114,28.837915,26.374237,23.906654,21.442978,18.9793,16.511717,14.450192,12.388668,10.323239,8.261715,6.2001905,7.1880045,8.175818,9.163632,10.151445,11.139259,10.670732,10.202203,9.733675,9.269051,8.800523,8.281238,7.7619514,7.238762,6.719476,6.2001905,6.6413884,7.0786815,7.519879,7.9610763,8.398369,10.838621,13.2788725,15.719124,18.159374,20.599627,19.701614,18.799696,17.901684,16.999767,16.101755,17.226223,18.35069,19.475159,20.599627,21.724094,21.056442,20.384884,19.713327,19.045673,18.374117,18.3585,18.346786,18.33117,18.315552,18.299932,18.756748,19.213564,19.674282,20.131098,20.587914,20.50592,20.423927,20.341936,20.256039,20.174046,22.251188,24.328331,26.409376,28.486519,30.563662,29.025326,27.486992,25.948658,24.414227,22.875893,20.693333,18.514675,16.33602,14.153459,11.974802,10.721489,9.468176,8.218767,6.9654536,5.7121406,8.695104,11.678067,14.661031,17.643993,20.623053,21.103294,21.583536,22.063778,22.544018,23.02426,22.665054,22.305851,21.946646,21.583536,21.22433,18.366308,15.5082855,12.654168,9.796145,6.9381227,6.4422636,5.9464045,5.4505453,4.958591,4.462732,4.2050414,3.9473507,3.68966,3.4319696,3.174279,3.2757936,3.3734035,3.474918,3.5764325,3.6740425,8.882515,14.090988,19.29946,24.504028,29.712502,29.091702,28.470901,27.854006,27.233206,26.612406,25.101402,23.594303,22.0833,20.572296,19.061293,17.273075,15.488764,13.700547,11.912332,10.124115,9.956225,9.788337,9.6243515,9.456462,9.288573,8.823949,8.36323,7.898606,7.437886,6.9732623,7.262188,7.551114,7.8361354,8.125061,8.413987,7.367607,6.321227,5.278752,4.2323723,3.1859922,3.2211318,3.2562714,3.2914112,3.3265507,3.3616903,3.2289407,3.0922866,2.9556324,2.822883,2.6862288,2.951728,3.213323,3.474918,3.736513,3.998108,3.2914112,2.5808098,1.8702087,1.1596074,0.44900626,0.5544251,0.6559396,0.75745404,0.8589685,0.96438736,0.80040246,0.63641757,0.47633708,0.31235218,0.14836729,0.40996224,0.6715572,0.92924774,1.1908426,1.4485333,1.2337911,1.0151446,0.79649806,0.58175594,0.3631094,0.28892577,0.21864653,0.14446288,0.07418364,0.0,0.20302892,0.40605783,0.60908675,0.80821127,1.0112402,0.8862993,0.75745404,0.62860876,0.5036679,0.37482262,0.3279698,0.28111696,0.23426414,0.1835069,0.13665408,0.9058213,1.678893,2.4480603,3.2172275,3.9863946,3.213323,2.4441557,1.6710842,0.8980125,0.12494087,0.58566034,1.0502841,1.5110037,1.9756275,2.436347,2.2684577,2.1005683,1.9365835,1.7686942,1.6008049,1.3118792,1.0190489,0.7301232,0.44119745,0.14836729,0.1756981,0.19912452,0.22645533,0.24988174,0.27330816,0.29673457,0.31625658,0.3357786,0.3553006,0.37482262,0.5466163,0.7145056,0.8862993,1.0541886,1.2259823,1.2415999,1.261122,1.2767396,1.2962615,1.3118792,1.2376955,1.1635119,1.0893283,1.0112402,0.93705654,2.182561,3.4280653,4.6735697,5.919074,7.1606736,7.0357327,6.9068875,6.7780423,6.6531014,6.524256,5.462259,4.4002614,3.338264,2.2762666,1.2142692,1.116659,1.0229534,0.92924774,0.8316377,0.737932,0.62860876,0.5231899,0.41386664,0.30844778,0.19912452,0.25769055,0.31625658,0.3709182,0.42948425,0.48805028,0.5192855,0.5544251,0.58566034,0.61689556,0.6481308,0.60127795,0.5505207,0.4997635,0.44900626,0.39824903,0.8980125,1.3938715,1.893635,2.3894942,2.8892577,2.7643168,2.6432803,2.5183394,2.397303,2.2762666,2.8306916,3.3890212,3.9473507,4.50568,5.0640097,5.989353,6.910792,7.8361354,8.761478,9.686822,9.561881,9.43694,9.311999,9.187058,9.062118,9.80005,10.537982,11.275913,12.013845,12.751778,13.583415,14.418958,15.254499,16.090042,16.925583,16.663988,16.406298,16.144703,15.883108,15.625418,14.528281,13.431144,12.334006,11.23687,10.135828,9.526741,8.913751,8.300759,7.687768,7.0747766,7.4105554,7.746334,8.078208,8.413987,8.749765,8.456935,8.164105,7.871275,7.578445,7.2856145,7.098203,6.9068875,6.715572,6.5281606,6.336845,5.755089,5.173333,4.591577,4.0059166,3.4241607,3.3538816,3.279698,3.2094188,3.135235,3.0610514,3.6467118,4.2323723,4.8180323,5.4036927,5.989353,6.715572,7.4417906,8.171914,8.898132,9.6243515,1.3743496,1.43682,1.4992905,1.5617609,1.6242313,1.6867018,1.7491722,1.8116426,1.8741131,1.9365835,1.999054,2.0888553,2.174752,2.260649,2.35045,2.436347,2.6237583,2.8111696,2.998581,3.1859922,3.3734035,3.5491016,3.7247996,3.900498,4.0761957,4.251894,4.474445,4.7009,4.9234514,5.1499066,5.376362,5.0640097,4.7516575,4.4393053,4.123049,3.8106966,3.4632049,3.1118085,2.7643168,2.4129205,2.0615244,1.698415,1.33921,0.97610056,0.61299115,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.37482262,0.38653582,0.39824903,0.41386664,0.42557985,0.43729305,0.44900626,0.46071947,0.47633708,0.48805028,0.4997635,0.97610056,1.4485333,1.9248703,2.4012074,2.87364,3.8380275,4.7985106,5.7628975,6.7233806,7.687768,7.898606,8.113348,8.324185,8.538928,8.749765,10.424754,12.099743,13.774731,15.449719,17.124708,16.164225,15.199838,14.239355,13.274967,12.31058,11.225157,10.135828,9.050405,7.9610763,6.8756523,5.786324,4.7009,3.611572,2.5261483,1.43682,1.5890918,1.737459,1.8858263,2.0380979,2.1864653,2.338737,2.4871042,2.639376,2.787743,2.9361105,3.7638438,4.5876727,5.4115014,6.239235,7.0630636,7.363703,7.6643414,7.9610763,8.261715,8.562354,7.3012323,6.036206,4.775084,3.513962,2.2489357,2.0380979,1.8233559,1.6125181,1.4016805,1.1869383,1.0737107,0.96438736,0.8511597,0.737932,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.0,0.999527,1.999054,2.998581,3.998108,5.001539,4.0761957,3.1508527,2.2255092,1.3001659,0.37482262,0.42557985,0.47633708,0.5231899,0.57394713,0.62470436,1.5617609,2.4988174,3.435874,4.376835,5.3138914,5.786324,6.262661,6.7389984,7.211431,7.687768,7.4886436,7.2856145,7.08649,6.8873653,6.688241,6.5867267,6.4891167,6.387602,6.2860875,6.1884775,6.699954,7.211431,7.726812,8.238289,8.749765,9.737579,10.725393,11.713207,12.70102,13.688834,13.4858055,13.286681,13.087557,12.888432,12.689307,13.251541,13.813775,14.376009,14.938243,15.500477,16.925583,18.35069,19.775797,21.200905,22.62601,26.760773,30.899439,35.038105,39.176773,43.311535,45.71274,48.11395,50.511253,52.91246,55.313667,55.887615,56.46156,57.039413,57.61336,58.187305,56.926186,55.66116,54.400036,53.138916,51.87389,47.512672,43.151455,38.78633,34.425114,30.063898,24.937418,19.810938,14.688361,9.561881,4.4393053,6.3251314,8.210958,10.100689,11.986515,13.8762455,13.813775,13.751305,13.688834,13.626364,13.563893,11.514082,9.464272,7.4105554,5.3607445,3.310933,7.348085,11.389141,15.426293,19.463446,23.500597,19.826555,16.148607,12.4745655,8.800523,5.12648,5.4505453,5.774611,6.098676,6.426646,6.7507114,7.7892823,8.823949,9.86252,10.901091,11.935758,10.38571,8.835662,7.2856145,5.735567,4.1894236,10.124115,16.062712,22.001307,27.935999,33.874596,40.199726,46.524857,52.84999,59.17512,65.50025,58.57384,51.651337,44.724926,37.79852,30.876013,30.66127,30.450434,30.235691,30.024853,29.814016,27.201971,24.586021,21.973976,19.36193,16.749886,14.473619,12.201257,9.924991,7.648724,5.376362,6.551587,7.726812,8.898132,10.073358,11.248583,10.573121,9.901564,9.226103,8.550641,7.8751793,7.5120697,7.1489606,6.785851,6.426646,6.0635366,5.8878384,5.7121406,5.5364423,5.3607445,5.1889505,8.113348,11.037745,13.962143,16.88654,19.810938,19.36193,18.912924,18.463919,18.011007,17.562002,17.226223,16.88654,16.55076,16.211079,15.875299,16.72646,17.573715,18.424873,19.276033,20.12329,19.998348,19.873407,19.748466,19.623526,19.498585,19.935879,20.37317,20.81437,21.251661,21.688955,21.22433,20.76361,20.298986,19.838268,19.373644,21.025206,22.67677,24.324427,25.975988,27.623646,26.136068,24.64849,23.160913,21.673336,20.18576,18.463919,16.738173,15.012426,13.286681,11.560935,10.674636,9.788337,8.898132,8.011833,7.125534,10.073358,13.025085,15.976814,18.924637,21.876366,22.036446,22.200432,22.364416,22.524496,22.688482,22.286327,21.888079,21.485926,21.087677,20.689428,17.948538,15.211552,12.4745655,9.737579,7.000593,6.461786,5.9268827,5.388075,4.8492675,4.3143644,4.0605783,3.8106966,3.5608149,3.310933,3.0610514,3.2992198,3.5373883,3.775557,4.0137253,4.251894,10.139732,16.023666,21.911505,27.799343,33.687183,32.773552,31.863827,30.950197,30.036566,29.12684,27.11217,25.101402,23.086731,21.075964,19.061293,17.24965,15.438006,13.626364,11.810817,9.999174,9.737579,9.475985,9.21439,8.94889,8.687295,8.499884,8.312472,8.125061,7.9376497,7.7502384,8.00012,8.250002,8.499884,8.749765,8.999647,7.687768,6.375889,5.0640097,3.7482262,2.436347,2.612045,2.787743,2.9634414,3.1391394,3.310933,3.1391394,2.9634414,2.787743,2.612045,2.436347,2.7018464,2.9634414,3.2250361,3.4866312,3.7482262,3.049338,2.35045,1.6515622,0.94876975,0.24988174,0.26159495,0.27330816,0.28892577,0.30063897,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.37482262,0.6871748,0.999527,1.3118792,1.6242313,1.3509232,1.0737107,0.80040246,0.5231899,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.3513962,0.57394713,0.80040246,1.0268579,1.2494087,1.0268579,0.80040246,0.57394713,0.3513962,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,0.74964523,0.9019169,1.0502841,1.1986516,1.3509232,1.4992905,1.2376955,0.97610056,0.7106012,0.44900626,0.18741131,0.21083772,0.23816854,0.26159495,0.28892577,0.31235218,0.3357786,0.3631094,0.38653582,0.41386664,0.43729305,0.46071947,0.48805028,0.5114767,0.5388075,0.5622339,0.5388075,0.5114767,0.48805028,0.46071947,0.43729305,0.44900626,0.46071947,0.47633708,0.48805028,0.4997635,2.0107672,3.5256753,5.036679,6.551587,8.062591,7.9610763,7.8634663,7.7619514,7.6643414,7.562827,6.3251314,5.087436,3.8497405,2.612045,1.3743496,1.261122,1.1517987,1.038571,0.92534333,0.81211567,0.6871748,0.5622339,0.43729305,0.31235218,0.18741131,0.26159495,0.3357786,0.41386664,0.48805028,0.5622339,0.58566034,0.61299115,0.63641757,0.6637484,0.6871748,0.61299115,0.5388075,0.46071947,0.38653582,0.31235218,0.94876975,1.5890918,2.2255092,2.8619268,3.4983444,3.310933,3.1235218,2.9361105,2.7486992,2.5612879,3.1859922,3.8106966,4.4393053,5.0640097,5.688714,6.699954,7.7111945,8.726339,9.737579,10.748819,10.588739,10.424754,10.260769,10.100689,9.936704,10.651209,11.361811,12.076316,12.786918,13.501423,14.53609,15.57466,16.613232,17.651802,18.68647,18.401447,18.112522,17.823597,17.538574,17.24965,15.773785,14.297921,12.825961,11.350098,9.874233,9.0386915,8.1992445,7.363703,6.524256,5.688714,6.4110284,7.137247,7.8634663,8.58578,9.311999,9.198771,9.085544,8.976221,8.862993,8.749765,8.460839,8.175818,7.8868923,7.601871,7.3129454,6.4110284,5.5130157,4.6110992,3.7130866,2.8111696,2.7643168,2.7135596,2.6628022,2.612045,2.5612879,3.1625657,3.7638438,4.3612175,4.9624953,5.563773,6.2743745,6.98888,7.699481,8.413987,9.124588,1.3626363,1.43682,1.5070993,1.5812829,1.6515622,1.7257458,1.7491722,1.7686942,1.7921207,1.815547,1.8389735,1.901444,1.9639144,2.0263848,2.0888553,2.1513257,2.3738766,2.5964274,2.8189783,3.0415294,3.2640803,3.4632049,3.6662338,3.8692627,4.0722914,4.2753205,4.4705405,4.6657605,4.860981,5.056201,5.251421,5.017157,4.786797,4.552533,4.318269,4.087909,3.6857557,3.2875066,2.8892577,2.4871042,2.0888553,1.7140326,1.33921,0.96438736,0.58566034,0.21083772,0.23426414,0.25769055,0.28111696,0.30063897,0.3240654,0.40996224,0.4958591,0.58175594,0.6637484,0.74964523,0.6754616,0.60127795,0.5231899,0.44900626,0.37482262,0.3240654,0.27330816,0.22645533,0.1756981,0.12494087,0.1678893,0.21083772,0.25378615,0.29673457,0.3357786,0.5114767,0.6832704,0.8550641,1.0268579,1.1986516,1.261122,1.319688,1.3782539,1.4407244,1.4992905,1.9443923,2.3855898,2.8267872,3.2718892,3.7130866,4.513489,5.3177958,6.1181984,6.9225054,7.726812,8.19534,8.663869,9.136301,9.60483,10.073358,11.393045,12.708829,14.028518,15.344301,16.663988,15.664462,14.668839,13.6693125,12.67369,11.674163,10.565312,9.456462,8.343708,7.2348576,6.126007,5.2358036,4.3455997,3.455396,2.5651922,1.6749885,1.7999294,1.9248703,2.0498111,2.174752,2.2996929,2.358259,2.416825,2.4714866,2.5300527,2.5886188,3.2757936,3.9668727,4.657952,5.349031,6.036206,6.481308,6.9225054,7.363703,7.8088045,8.250002,7.2739015,6.3017054,5.3256044,4.349504,3.3734035,2.8892577,2.4051118,1.9209659,1.43682,0.94876975,0.8706817,0.78868926,0.7106012,0.62860876,0.5505207,0.45291066,0.3553006,0.25769055,0.16008049,0.062470436,0.8511597,1.6359446,2.4246337,3.213323,3.998108,3.2718892,2.541766,1.8116426,1.0815194,0.3513962,0.38653582,0.42557985,0.46071947,0.4997635,0.5388075,1.6008049,2.6628022,3.7247996,4.786797,5.8487945,6.5008297,7.1567693,7.8088045,8.460839,9.112875,8.81614,8.52331,8.226576,7.9337454,7.6370106,7.605776,7.570636,7.5394006,7.5081654,7.47693,7.8361354,8.19534,8.554545,8.913751,9.276859,10.096785,10.916709,11.736633,12.556558,13.376482,13.306203,13.239828,13.173453,13.103174,13.036799,13.845011,14.653222,15.461433,16.26574,17.073952,18.54591,20.021774,21.493734,22.965694,24.437654,28.486519,32.53148,36.580345,40.62921,44.67417,45.92358,47.17689,48.4263,49.67571,50.925117,51.323368,51.721615,52.115963,52.51421,52.91246,51.30775,49.70304,48.09833,46.49362,44.888912,40.953274,37.01764,33.082,29.146362,25.210726,20.935406,16.65618,12.380859,8.101635,3.8263142,5.8683167,7.910319,9.952321,11.994324,14.036326,14.223738,14.407245,14.590752,14.778163,14.96167,12.654168,10.346666,8.039165,5.7316628,3.4241607,7.039637,10.655114,14.27059,17.886066,21.501543,18.354595,15.211552,12.064603,8.921559,5.774611,6.3407493,6.9068875,7.4691215,8.03526,8.601398,9.366661,10.135828,10.901091,11.6702585,12.439425,10.803481,9.171441,7.5394006,5.9073606,4.2753205,9.151918,14.028518,18.90902,23.785618,28.662216,34.284557,39.906895,45.529236,51.151573,56.773914,51.553726,46.329636,41.105545,35.88536,30.66127,30.551949,30.43872,30.325493,30.212265,30.099037,27.553368,25.0116,22.46593,19.92026,17.37459,14.95386,12.529227,10.108498,7.6838636,5.263134,6.2431393,7.223144,8.203149,9.183154,10.163159,9.749292,9.331521,8.917655,8.503788,8.086017,7.7385254,7.3910336,7.043542,6.6960497,6.348558,6.75852,7.164578,7.570636,7.9805984,8.386656,10.502842,12.619028,14.73131,16.847496,18.963682,18.600573,18.241367,17.882162,17.522957,17.163752,17.460487,17.757221,18.053955,18.35069,18.651329,19.229181,19.810938,20.388788,20.970545,21.548395,21.079868,20.61134,20.138906,19.670378,19.20185,19.311174,19.420496,19.52982,19.639143,19.748466,19.092527,18.436588,17.776743,17.120804,16.46096,17.99539,19.525915,21.060347,22.590872,24.125301,23.371752,22.618202,21.868557,21.115007,20.361458,19.393166,18.420969,17.452679,16.484386,15.51219,14.668839,13.821584,12.978233,12.130978,11.287627,13.610746,15.933866,18.256985,20.5762,22.899319,22.62601,22.356607,22.0833,21.809992,21.536682,21.06425,20.587914,20.111576,19.639143,19.162806,16.808453,14.454097,12.095839,9.741484,7.387129,7.8634663,8.335898,8.812236,9.288573,9.761005,10.510651,11.2642,12.013845,12.763491,13.513136,13.759113,14.008995,14.254972,14.50095,14.750832,17.874353,20.99397,24.117493,27.241014,30.360632,29.400148,28.435762,27.475279,26.510891,25.550407,24.086258,22.618202,21.15405,19.689901,18.22575,16.515621,14.809398,13.103174,11.393045,9.686822,9.237816,8.78881,8.335898,7.8868923,7.437886,7.355894,7.2739015,7.191909,7.1060123,7.0240197,7.5120697,8.00012,8.488171,8.976221,9.464272,8.101635,6.7389984,5.376362,4.0137253,2.6510892,2.6940374,2.7408905,2.7838387,2.8306916,2.87364,2.7447948,2.6159496,2.4831998,2.3543546,2.2255092,2.4441557,2.6588979,2.8775444,3.096191,3.310933,2.690133,2.069333,1.4446288,0.8238289,0.19912452,0.21083772,0.21864653,0.23035973,0.23816854,0.24988174,0.23426414,0.21864653,0.20693332,0.19131571,0.1756981,0.45291066,0.7301232,1.0073358,1.2845483,1.5617609,1.3157835,1.0737107,0.8277333,0.58175594,0.3357786,0.27721256,0.21864653,0.15617609,0.09761006,0.039044023,0.093705654,0.14836729,0.20302892,0.25769055,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.07418364,0.08199245,0.093705654,0.10151446,0.113227665,0.28892577,0.46852827,0.6442264,0.8238289,0.999527,0.8199245,0.64032197,0.46071947,0.28111696,0.10151446,0.21474212,0.3318742,0.44510186,0.5583295,0.6754616,1.116659,1.5617609,2.0029583,2.4441557,2.8892577,2.463678,2.0380979,1.6125181,1.1869383,0.76135844,0.7262188,0.6910792,0.6559396,0.62079996,0.58566034,0.7066968,0.8277333,0.94876975,1.0659018,1.1869383,1.3118792,1.43682,1.5617609,1.6867018,1.8116426,1.6086137,1.4055848,1.2064602,1.0034313,0.80040246,0.79649806,0.79649806,0.79259366,0.78868926,0.78868926,1.9561055,3.1235218,4.290938,5.4583545,6.6257706,6.6335793,6.6452928,6.6531014,6.6648145,6.676528,5.606722,4.5408196,3.4710135,2.4051118,1.33921,1.2259823,1.116659,1.0073358,0.8980125,0.78868926,0.6715572,0.5583295,0.44119745,0.3279698,0.21083772,0.28111696,0.3513962,0.42167544,0.49195468,0.5622339,0.5700427,0.57785153,0.58566034,0.59346914,0.60127795,0.5388075,0.47633708,0.41386664,0.3513962,0.28892577,0.9878138,1.6867018,2.3855898,3.0883822,3.78727,3.7794614,3.7716527,3.7638438,3.7560349,3.7482262,4.318269,4.8883114,5.4583545,6.028397,6.5984397,7.3988423,8.19534,8.991838,9.788337,10.588739,10.71368,10.838621,10.963562,11.088503,11.213444,12.341816,13.466284,14.594656,15.723028,16.8514,18.401447,19.9554,21.509352,23.0594,24.613352,23.648964,22.688482,21.724094,20.76361,19.799223,18.073479,16.351637,14.625891,12.900145,11.174399,10.397423,9.620447,8.843472,8.066495,7.2856145,7.9766936,8.667773,9.358852,10.046027,10.737106,10.553599,10.373997,10.19049,10.006983,9.823476,9.507219,9.190963,8.870802,8.554545,8.238289,7.3324676,6.426646,5.520825,4.618908,3.7130866,3.521771,3.3265507,3.135235,2.9439192,2.7486992,3.2094188,3.6662338,4.123049,4.579864,5.036679,5.7316628,6.426646,7.1216297,7.816613,8.511597,1.3509232,1.4329157,1.5149081,1.5969005,1.678893,1.7608855,1.7452679,1.7257458,1.7101282,1.6906061,1.6749885,1.7140326,1.7491722,1.7882162,1.8233559,1.8623998,2.1200905,2.377781,2.6354716,2.893162,3.1508527,3.3812122,3.611572,3.8419318,4.068387,4.298747,4.466636,4.630621,4.794606,4.958591,5.12648,4.9742084,4.8219366,4.6657605,4.513489,4.3612175,3.912211,3.4632049,3.0141985,2.5612879,2.1122816,1.7257458,1.33921,0.94876975,0.5622339,0.1756981,0.25769055,0.339683,0.42167544,0.5036679,0.58566034,0.7340276,0.8784905,1.0229534,1.1674163,1.3118792,1.175225,1.038571,0.9019169,0.76135844,0.62470436,0.5388075,0.44900626,0.3631094,0.27330816,0.18741131,0.21083772,0.23426414,0.25378615,0.27721256,0.30063897,0.63251317,0.96438736,1.2962615,1.6281357,1.9639144,2.069333,2.1786566,2.2840753,2.3933985,2.4988174,2.9087796,3.3187418,3.7287042,4.138666,4.548629,5.192855,5.833177,6.477403,7.1216297,7.7619514,8.488171,9.218294,9.944512,10.670732,11.400854,12.361338,13.32182,14.278399,15.238882,16.199366,15.168603,14.133936,13.103174,12.068507,11.037745,9.905469,8.773191,7.6409154,6.5086384,5.376362,4.6813784,3.9902992,3.2992198,2.6042364,1.9131571,2.0107672,2.1122816,2.2137961,2.3114061,2.4129205,2.377781,2.3426414,2.3075018,2.2723622,2.2372224,2.7916477,3.3460727,3.9044023,4.4588275,5.0132523,5.5989127,6.180669,6.7663293,7.3519893,7.9376497,7.250475,6.5633,5.8761253,5.1889505,4.5017757,3.7443218,2.9868677,2.2294137,1.4680552,0.7106012,0.6637484,0.61689556,0.5700427,0.5231899,0.47633708,0.40605783,0.3357786,0.26549935,0.19522011,0.12494087,0.698888,1.2767396,1.8506867,2.4246337,2.998581,2.463678,1.9287747,1.3938715,0.8589685,0.3240654,0.3513962,0.37482262,0.39824903,0.42557985,0.44900626,1.6359446,2.8267872,4.0137253,5.2006636,6.387602,7.2192397,8.046973,8.878611,9.706344,10.537982,10.147541,9.757101,9.366661,8.976221,8.58578,8.62092,8.65606,8.691199,8.726339,8.761478,8.968412,9.17925,9.386183,9.593117,9.80005,10.452085,11.10412,11.756155,12.408191,13.06413,13.1266,13.192975,13.25935,13.32182,13.388195,14.438479,15.492668,16.546856,17.597141,18.651329,20.170141,21.688955,23.211672,24.730484,26.249296,30.20836,34.16352,38.122585,42.081646,46.036808,46.13832,46.23593,46.337444,46.43896,46.53657,46.75912,46.977768,47.196415,47.418964,47.63761,45.689316,43.74102,41.796627,39.848328,37.900032,34.39388,30.883821,27.377668,23.871515,20.361458,16.933393,13.501423,10.073358,6.6413884,3.213323,5.4115014,7.605776,9.803954,12.002132,14.200311,14.633699,15.063184,15.4965725,15.929961,16.36335,13.798158,11.232965,8.667773,6.1025805,3.5373883,6.7311897,9.921086,13.114887,16.30869,19.498585,16.88654,14.27059,11.654641,9.0386915,6.426646,7.230953,8.03526,8.839567,9.643873,10.44818,10.947944,11.443803,11.943566,12.439425,12.939189,11.221252,9.507219,7.793187,6.0791545,4.3612175,8.179723,11.998228,15.816733,19.631334,23.44984,28.369387,33.288933,38.20848,43.13193,48.05148,44.52971,41.01184,37.49007,33.9683,30.450434,30.43872,30.423103,30.411388,30.399675,30.387962,27.908667,25.433277,22.953981,20.47859,17.999294,15.430198,12.861101,10.2881,7.719003,5.1499066,5.9346914,6.719476,7.504261,8.289046,9.073831,8.921559,8.765383,8.609207,8.456935,8.300759,7.968885,7.633106,7.3012323,6.969358,6.6374836,7.629202,8.617016,9.608734,10.596548,11.588266,12.892336,14.196406,15.504381,16.808453,18.112522,17.843119,17.573715,17.30431,17.031002,16.761599,17.694752,18.627903,19.561056,20.494207,21.423454,21.735807,22.044254,22.356607,22.665054,22.973503,22.161386,21.345367,20.529346,19.713327,18.90121,18.682566,18.463919,18.249176,18.030529,17.811884,16.960724,16.10566,15.254499,14.40334,13.548276,14.965574,16.378967,17.796265,19.20966,20.623053,20.607435,20.591818,20.572296,20.556679,20.537155,20.322414,20.107672,19.89293,19.678188,19.463446,18.659138,17.858736,17.054428,16.254026,15.449719,17.14423,18.838741,20.53325,22.231667,23.926178,23.215576,22.508879,21.802181,21.095486,20.388788,19.838268,19.287746,18.737226,18.186707,17.636185,15.664462,13.692739,11.721016,9.749292,7.773665,9.261242,10.748819,12.236397,13.723974,15.211552,16.960724,18.7138,20.462973,22.212145,23.961317,24.219007,24.476698,24.734388,24.992079,25.24977,25.608974,25.964275,26.32348,26.678782,27.037985,26.026745,25.0116,24.00036,22.98912,21.973976,21.056442,20.138906,19.221373,18.303837,17.386303,15.785499,14.180789,12.579984,10.979179,9.37447,8.738052,8.101635,7.461313,6.824895,6.1884775,6.211904,6.2314262,6.2548523,6.278279,6.3017054,7.0240197,7.7502384,8.476458,9.198771,9.924991,8.511597,7.098203,5.688714,4.2753205,2.8619268,2.77603,2.6940374,2.6081407,2.522244,2.436347,2.3543546,2.2684577,2.182561,2.096664,2.0107672,2.1864653,2.358259,2.5300527,2.7018464,2.87364,2.330928,1.7843118,1.2415999,0.6949836,0.14836729,0.15617609,0.1639849,0.1717937,0.1796025,0.18741131,0.20693332,0.22645533,0.24597734,0.26940376,0.28892577,0.5309987,0.77307165,1.0151446,1.2572175,1.4992905,1.2845483,1.0698062,0.8550641,0.64032197,0.42557985,0.3553006,0.28502136,0.21474212,0.14446288,0.07418364,0.12103647,0.1717937,0.21864653,0.26549935,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.07027924,0.078088045,0.08589685,0.093705654,0.10151446,0.23035973,0.359205,0.49195468,0.62079996,0.74964523,0.61689556,0.48024148,0.3435874,0.21083772,0.07418364,0.1796025,0.28502136,0.39044023,0.4958591,0.60127795,1.3353056,2.069333,2.803361,3.541293,4.2753205,3.6857557,3.1000953,2.514435,1.9248703,1.33921,1.2415999,1.1478943,1.0541886,0.95657855,0.8628729,1.077615,1.2923572,1.5070993,1.7218413,1.9365835,2.1630387,2.3855898,2.612045,2.8385005,3.0610514,2.6823244,2.3035975,1.9209659,1.542239,1.1635119,1.1439898,1.1283722,1.1088502,1.0932326,1.0737107,1.8975395,2.7213683,3.541293,4.365122,5.1889505,5.3060827,5.4271193,5.548156,5.6691923,5.786324,4.8883114,3.9942036,3.096191,2.1981785,1.3001659,1.1908426,1.0854238,0.97610056,0.8706817,0.76135844,0.6559396,0.5544251,0.44900626,0.3435874,0.23816854,0.30063897,0.3670138,0.43338865,0.4958591,0.5622339,0.5544251,0.5427119,0.5309987,0.5231899,0.5114767,0.46071947,0.41386664,0.3631094,0.31235218,0.26159495,1.0268579,1.7882162,2.5495746,3.310933,4.0761957,4.2479897,4.4197836,4.591577,4.7633705,4.939069,5.45445,5.9659266,6.481308,6.996689,7.5120697,8.093826,8.675582,9.261242,9.8429985,10.424754,10.838621,11.248583,11.66245,12.076316,12.486279,14.028518,15.570756,17.1169,18.659138,20.201378,22.266806,24.33614,26.401567,28.470901,30.53633,28.900385,27.260536,25.624592,23.988647,22.348799,20.37317,18.401447,16.42582,14.450192,12.4745655,11.756155,11.04165,10.323239,9.60483,8.886419,9.542359,10.198298,10.8542385,11.506273,12.162213,11.908427,11.6585455,11.404759,11.150972,10.901091,10.553599,10.206107,9.858616,9.511124,9.163632,8.253906,7.3441806,6.4305506,5.520825,4.6110992,4.279225,3.9434462,3.6076677,3.2718892,2.9361105,3.252367,3.5686235,3.8809757,4.1972322,4.513489,5.1889505,5.8683167,6.5437784,7.223144,7.898606,1.33921,1.4290112,1.5227169,1.6164225,1.7062237,1.7999294,1.7413634,1.6867018,1.6281357,1.5695697,1.5110037,1.5266213,1.5383345,1.5500476,1.5617609,1.5734742,1.8663043,2.1591344,2.4519646,2.7447948,3.0376248,3.2953155,3.5530062,3.8106966,4.068387,4.3260775,4.4588275,4.5954814,4.728231,4.8648853,5.001539,4.927356,4.853172,4.7828927,4.7087092,4.6384296,4.138666,3.638903,3.1391394,2.639376,2.135708,1.737459,1.33921,0.93705654,0.5388075,0.13665408,0.28111696,0.42167544,0.5661383,0.7066968,0.8511597,1.0541886,1.261122,1.4641509,1.6710842,1.8741131,1.6749885,1.475864,1.2767396,1.0737107,0.8745861,0.74964523,0.62470436,0.4997635,0.37482262,0.24988174,0.25378615,0.25378615,0.25769055,0.26159495,0.26159495,0.75354964,1.2494087,1.7413634,2.233318,2.7252727,2.8814487,3.0337205,3.1898966,3.3460727,3.4983444,3.8770714,4.2557983,4.630621,5.009348,5.388075,5.8683167,6.3524623,6.8366084,7.3168497,7.800996,8.784905,9.768814,10.756628,11.740538,12.724447,13.325725,13.930907,14.532186,15.133463,15.738646,14.668839,13.602938,12.533132,11.46723,10.401327,9.245625,8.089922,6.9342184,5.7785153,4.6267166,4.1308575,3.6349986,3.1391394,2.6432803,2.1513257,2.2255092,2.2996929,2.3738766,2.4480603,2.5261483,2.397303,2.2684577,2.1435168,2.0146716,1.8858263,2.3075018,2.7291772,3.1469483,3.5686235,3.9863946,4.716518,5.4427366,6.168956,6.899079,7.6252975,7.223144,6.824895,6.426646,6.0244927,5.6262436,4.5954814,3.5647192,2.533957,1.5031948,0.47633708,0.46071947,0.44510186,0.42948425,0.41386664,0.39824903,0.359205,0.31625658,0.27330816,0.23035973,0.18741131,0.5505207,0.9136301,1.2767396,1.6359446,1.999054,1.6593709,1.319688,0.98000497,0.64032197,0.30063897,0.31235218,0.3240654,0.3357786,0.3513962,0.3631094,1.6749885,2.9868677,4.298747,5.610626,6.9264097,7.9337454,8.941081,9.948417,10.955752,11.963089,11.478943,10.990892,10.506746,10.0226,9.538455,9.639969,9.741484,9.846903,9.948417,10.049932,10.104593,10.159255,10.213917,10.268578,10.323239,10.81129,11.295436,11.779582,12.263727,12.751778,12.946998,13.146122,13.341343,13.540467,13.735687,15.035853,16.332115,17.628376,18.928543,20.224804,21.794373,23.360039,24.925705,26.495274,28.06094,31.930202,35.79556,39.66482,43.534084,47.399445,46.34916,45.298874,44.248592,43.198307,42.14802,42.19097,42.23392,42.276867,42.319817,42.362766,40.07088,37.7829,35.491016,33.203037,30.911152,27.83058,24.75391,21.673336,18.592764,15.51219,12.93138,10.346666,7.7658563,5.181142,2.6003318,4.950782,7.3051367,9.659492,12.009941,14.364296,15.043662,15.723028,16.402393,17.08176,17.761126,14.938243,12.119265,9.296382,6.473499,3.6506162,6.4188375,9.190963,11.959184,14.73131,17.49953,15.41458,13.329629,11.2446785,9.159728,7.0747766,8.121157,9.163632,10.2100115,11.256392,12.298867,12.529227,12.755682,12.982138,13.208592,13.438952,11.639023,9.8429985,8.043069,6.2470436,4.4510183,7.2075267,9.964035,12.724447,15.480955,18.237463,22.454218,26.67097,30.89163,35.108383,39.325138,37.505688,35.69014,33.87069,32.05514,30.235691,30.325493,30.411388,30.50119,30.587088,30.67689,28.263968,25.854952,23.445936,21.036919,18.623999,15.906535,13.189071,10.471607,7.7541428,5.036679,5.6262436,6.2158084,6.8092775,7.3988423,7.988407,8.093826,8.1992445,8.300759,8.406178,8.511597,8.19534,7.8790836,7.558923,7.2426662,6.9264097,8.495979,10.069453,11.642927,13.216402,14.785972,15.281831,15.77769,16.273548,16.769407,17.261362,17.08176,16.902157,16.722555,16.542952,16.36335,17.929016,19.498585,21.06425,22.63382,24.199486,24.23853,24.281477,24.320522,24.359566,24.39861,23.239002,22.079395,20.919786,19.76018,18.600573,18.053955,17.511244,16.964628,16.421915,15.875299,14.828919,13.778636,12.732256,11.685876,10.6355915,11.935758,13.232019,14.528281,15.828446,17.124708,17.843119,18.56153,19.276033,19.994444,20.712854,21.251661,21.794373,22.333181,22.871988,23.410795,22.653341,21.891983,21.130625,20.37317,19.611813,20.68162,21.74752,22.813423,23.883228,24.949131,23.809046,22.665054,21.521065,20.38098,19.23699,18.612286,17.987581,17.362877,16.738173,16.113468,14.520472,12.93138,11.342289,9.753197,8.164105,10.662923,13.16174,15.664462,18.163279,20.662096,23.410795,26.163399,28.912098,31.660797,34.413403,34.6789,34.948303,35.213802,35.483208,35.748707,33.343594,30.93458,28.525562,26.120451,23.711435,22.649437,21.58744,20.525442,19.463446,18.401447,18.030529,17.65961,17.288692,16.921679,16.55076,15.051471,13.556085,12.056794,10.561408,9.062118,8.238289,7.4144597,6.5867267,5.7628975,4.939069,5.0640097,5.192855,5.3217,5.446641,5.575486,6.5359693,7.5003567,8.460839,9.425227,10.38571,8.925464,7.461313,6.001066,4.5369153,3.076669,2.8619268,2.6432803,2.4285383,2.2137961,1.999054,1.9600099,1.9209659,1.8819219,1.8389735,1.7999294,1.9287747,2.0537157,2.182561,2.3114061,2.436347,1.9717231,1.5031948,1.0346665,0.5661383,0.10151446,0.10541886,0.10932326,0.113227665,0.12103647,0.12494087,0.1796025,0.23426414,0.28892577,0.3435874,0.39824903,0.60908675,0.8160201,1.0229534,1.2298868,1.43682,1.2533131,1.0659018,0.8823949,0.698888,0.5114767,0.43338865,0.3513962,0.27330816,0.19131571,0.113227665,0.15227169,0.19131571,0.23426414,0.27330816,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.06637484,0.07418364,0.078088045,0.08199245,0.08589685,0.1717937,0.25378615,0.3357786,0.41777104,0.4997635,0.40996224,0.32016098,0.23035973,0.14055848,0.05075723,0.14446288,0.23816854,0.3357786,0.42948425,0.5231899,1.5539521,2.5808098,3.6076677,4.6345253,5.661383,4.911738,4.1620927,3.4124475,2.6628022,1.9131571,1.756981,1.6008049,1.4485333,1.2923572,1.1361811,1.4485333,1.756981,2.069333,2.377781,2.6862288,3.0141985,3.338264,3.6623292,3.9863946,4.3143644,3.7560349,3.1977055,2.639376,2.0810463,1.5266213,1.4914817,1.4602464,1.4290112,1.3938715,1.3626363,1.8389735,2.3192148,2.795552,3.2718892,3.7482262,3.978586,4.2089458,4.4393053,4.6696653,4.900025,4.173806,3.4436827,2.717464,1.9912452,1.261122,1.1557031,1.0541886,0.94876975,0.8433509,0.737932,0.6442264,0.5466163,0.45291066,0.359205,0.26159495,0.3240654,0.38263142,0.44119745,0.5036679,0.5622339,0.5349031,0.5075723,0.48024148,0.45291066,0.42557985,0.38653582,0.3513962,0.31235218,0.27330816,0.23816854,1.0619974,1.8858263,2.7135596,3.5373883,4.3612175,4.716518,5.067914,5.4193106,5.7707067,6.126007,6.5867267,7.043542,7.504261,7.9649806,8.4257,8.792714,9.159728,9.526741,9.893755,10.260769,10.963562,11.66245,12.361338,13.06413,13.763018,15.719124,17.679134,19.635239,21.591345,23.551353,26.132164,28.716879,31.297688,33.878498,36.46321,34.151806,31.836496,29.52509,27.213684,24.898373,22.67677,20.45126,18.22575,16.00024,13.774731,13.118792,12.458947,11.803008,11.143164,10.487225,11.108025,11.728825,12.34572,12.96652,13.58732,13.263254,12.943093,12.619028,12.298867,11.974802,11.596075,11.221252,10.8425255,10.4637985,10.088976,9.171441,8.257811,7.3441806,6.426646,5.5130157,5.036679,4.5564375,4.0801005,3.6037633,3.1235218,3.2992198,3.4710135,3.6428072,3.814601,3.9863946,4.646239,5.3060827,5.9659266,6.6257706,7.2856145,1.3235924,1.4290112,1.5305257,1.6320401,1.7335546,1.8389735,1.7413634,1.6437533,1.5461433,1.4485333,1.3509232,1.33921,1.3235924,1.3118792,1.3001659,1.2884527,1.6164225,1.9443923,2.2684577,2.5964274,2.9243972,3.2094188,3.49444,3.7794614,4.0644827,4.349504,4.454923,4.560342,4.6657605,4.7711797,4.8765984,4.884407,4.8883114,4.8961205,4.903929,4.911738,4.3612175,3.8106966,3.2640803,2.7135596,2.1630387,1.7491722,1.33921,0.92534333,0.5114767,0.10151446,0.30063897,0.5036679,0.7066968,0.9097257,1.1127546,1.3782539,1.6437533,1.9092526,2.1708477,2.436347,2.174752,1.9131571,1.6515622,1.3860629,1.1244678,0.96438736,0.80040246,0.63641757,0.47633708,0.31235218,0.29673457,0.27721256,0.26159495,0.24207294,0.22645533,0.8784905,1.5305257,2.182561,2.8345962,3.4866312,3.68966,3.892689,4.095718,4.298747,4.5017757,4.845363,5.1889505,5.5364423,5.8800297,6.223617,6.547683,6.871748,7.191909,7.5159745,7.8361354,9.081639,10.323239,11.564839,12.806439,14.051944,14.294017,14.539994,14.785972,15.031949,15.274021,14.17298,13.0719385,11.966993,10.865952,9.761005,8.58578,7.406651,6.2314262,5.0522966,3.873167,3.5764325,3.279698,2.9829633,2.6862288,2.3855898,2.436347,2.4871042,2.5378613,2.5886188,2.639376,2.416825,2.1981785,1.9756275,1.756981,1.5383345,1.8233559,2.1083772,2.3933985,2.67842,2.9634414,3.8341231,4.7009,5.571582,6.4422636,7.3129454,7.1997175,7.08649,6.9732623,6.8639393,6.7507114,5.446641,4.1464753,2.8424048,1.5383345,0.23816854,0.25378615,0.27330816,0.28892577,0.30844778,0.3240654,0.30844778,0.29673457,0.28111696,0.26549935,0.24988174,0.39824903,0.5505207,0.698888,0.8511597,0.999527,0.8550641,0.7106012,0.5661383,0.42167544,0.27330816,0.27330816,0.27330816,0.27330816,0.27330816,0.27330816,1.7140326,3.1508527,4.5876727,6.0244927,7.461313,8.648251,9.8312845,11.018223,12.201257,13.388195,12.806439,12.228588,11.6468315,11.06898,10.487225,10.6590185,10.826907,10.998701,11.166591,11.338385,11.240774,11.143164,11.045554,10.947944,10.850334,11.166591,11.486752,11.803008,12.119265,12.439425,12.767395,13.09927,13.427239,13.759113,14.087084,15.629322,17.17156,18.7138,20.256039,21.798277,23.4147,25.031122,26.64364,28.260063,29.876486,33.652042,37.431503,41.20706,44.986523,48.76208,46.5639,44.36182,42.16364,39.961555,37.76338,37.626724,37.493977,37.357323,37.220665,37.087917,34.45635,31.820879,29.189312,26.557745,23.926178,21.271183,18.620094,15.969006,13.314012,10.662923,8.929368,7.191909,5.4583545,3.7208953,1.9873407,4.493967,7.000593,9.511124,12.01775,14.524376,15.453624,16.378967,17.308216,18.233559,19.162806,16.082233,13.001659,9.921086,6.8405128,3.7638438,6.1103897,8.456935,10.803481,13.153932,15.500477,13.946525,12.388668,10.834716,9.280765,7.726812,9.01136,10.295909,11.580457,12.8650055,14.149553,14.106606,14.063657,14.020708,13.981665,13.938716,12.056794,10.178777,8.296855,6.4188375,4.5369153,6.2353306,7.9337454,9.628256,11.326671,13.025085,16.539047,20.053009,23.570877,27.084839,30.5988,30.485573,30.36844,30.255213,30.13808,30.024853,30.212265,30.399675,30.587088,30.774498,30.96191,28.619268,26.276627,23.933987,21.591345,19.248703,16.386776,13.520945,10.655114,7.7892823,4.9234514,5.3217,5.716045,6.1103897,6.504734,6.899079,7.266093,7.629202,7.996216,8.359325,8.726339,8.421796,8.121157,7.816613,7.5159745,7.211431,9.366661,11.521891,13.677121,15.832351,17.987581,17.671324,17.358973,17.042715,16.72646,16.414106,16.324306,16.2306,16.140799,16.050997,15.961197,18.163279,20.369267,22.57135,24.773432,26.975515,26.745155,26.514795,26.284435,26.054077,25.823717,24.320522,22.813423,21.310228,19.803127,18.299932,17.429253,16.554665,15.683984,14.809398,13.938716,12.693212,11.4516115,10.2100115,8.968412,7.726812,8.905942,10.085071,11.2642,12.44333,13.626364,15.078801,16.531239,17.983677,19.436115,20.888552,22.18091,23.47717,24.773432,26.06579,27.362051,26.64364,25.929136,25.210726,24.492315,23.773905,24.215103,24.6563,25.093594,25.53479,25.975988,24.39861,22.821232,21.243853,19.666473,18.089096,17.386303,16.687416,15.988527,15.285735,14.586847,13.380386,12.173926,10.963562,9.757101,8.550641,12.064603,15.57466,19.088623,22.59868,26.112642,29.860868,33.613,37.361225,41.113358,44.861584,45.138794,45.416008,45.69322,45.974335,46.25155,41.078217,35.904884,30.73155,25.558218,20.388788,19.276033,18.163279,17.050524,15.93777,14.825015,15.000713,15.180316,15.356014,15.535617,15.711315,14.321347,12.927476,11.533605,10.143637,8.749765,7.7385254,6.7233806,5.7121406,4.7009,3.6857557,3.9200199,4.154284,4.3846436,4.618908,4.8492675,6.0518236,7.250475,8.449126,9.651682,10.850334,9.339331,7.824422,6.3134184,4.7985106,3.2875066,2.9439192,2.5964274,2.25284,1.9092526,1.5617609,1.5656652,1.5734742,1.5773785,1.5812829,1.5890918,1.6710842,1.7530766,1.8350691,1.9170616,1.999054,1.6086137,1.2181735,0.8316377,0.44119745,0.05075723,0.05075723,0.05466163,0.058566034,0.058566034,0.062470436,0.15227169,0.24207294,0.3318742,0.42167544,0.5114767,0.6832704,0.8589685,1.0307622,1.2025559,1.3743496,1.2181735,1.0659018,0.9097257,0.75354964,0.60127795,0.5114767,0.42167544,0.3318742,0.23816854,0.14836729,0.1835069,0.21474212,0.24597734,0.28111696,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.06637484,0.06637484,0.07027924,0.07418364,0.07418364,0.10932326,0.14446288,0.1796025,0.21474212,0.24988174,0.20693332,0.16008049,0.113227665,0.07027924,0.023426414,0.10932326,0.19522011,0.28111696,0.3631094,0.44900626,1.7686942,3.0883822,4.4119744,5.7316628,7.0513506,6.13772,5.22409,4.3143644,3.4007344,2.4871042,2.2723622,2.05762,1.8428779,1.6281357,1.4133936,1.8194515,2.2216048,2.6276627,3.0337205,3.435874,3.8614538,4.2870336,4.7126136,5.138193,5.563773,4.825841,4.0918136,3.357786,2.6237583,1.8858263,1.8389735,1.7921207,1.7452679,1.698415,1.6515622,1.7843118,1.9131571,2.0459068,2.1786566,2.3114061,2.6510892,2.9907722,3.3343596,3.6740425,4.0137253,3.455396,2.8970666,2.338737,1.7843118,1.2259823,1.1205635,1.0190489,0.91753453,0.8160201,0.7106012,0.62860876,0.5427119,0.45681506,0.3709182,0.28892577,0.3435874,0.39824903,0.45291066,0.5075723,0.5622339,0.5192855,0.47243267,0.42557985,0.38263142,0.3357786,0.31235218,0.28892577,0.26159495,0.23816854,0.21083772,1.1010414,1.9873407,2.87364,3.7638438,4.650143,5.181142,5.716045,6.2470436,6.7780423,7.3129454,7.719003,8.121157,8.527214,8.933272,9.339331,9.491602,9.643873,9.796145,9.948417,10.100689,11.088503,12.076316,13.06413,14.048039,15.035853,17.409729,19.783606,22.153578,24.527454,26.90133,29.997522,33.09371,36.19381,39.29,42.386192,39.399323,36.412457,33.425587,30.43872,27.451853,24.976461,22.50107,20.025679,17.550287,15.074897,14.477524,13.88015,13.282777,12.685403,12.08803,12.67369,13.25935,13.841106,14.426766,15.012426,14.618082,14.227642,13.833297,13.442857,13.048512,12.642454,12.236397,11.826434,11.420377,11.014318,10.09288,9.171441,8.253906,7.3324676,6.4110284,5.794133,5.173333,4.552533,3.9317331,3.310933,3.3421683,3.3734035,3.4007344,3.4319696,3.4632049,4.1035266,4.747753,5.388075,6.0323014,6.676528,1.3118792,1.4251068,1.5383345,1.6515622,1.7608855,1.8741131,1.737459,1.6008049,1.4641509,1.3235924,1.1869383,1.1517987,1.1127546,1.0737107,1.038571,0.999527,1.3626363,1.7257458,2.0888553,2.4480603,2.8111696,3.1235218,3.435874,3.7482262,4.0605783,4.376835,4.4510183,4.5252023,4.5993857,4.6735697,4.7516575,4.8375545,4.9234514,5.0132523,5.099149,5.1889505,4.5876727,3.9863946,3.3890212,2.787743,2.1864653,1.7608855,1.33921,0.9136301,0.48805028,0.062470436,0.3240654,0.58566034,0.8511597,1.1127546,1.3743496,1.698415,2.0263848,2.35045,2.6745155,2.998581,2.6745155,2.35045,2.0263848,1.698415,1.3743496,1.175225,0.97610056,0.77307165,0.57394713,0.37482262,0.3357786,0.30063897,0.26159495,0.22645533,0.18741131,0.999527,1.8116426,2.6237583,3.435874,4.251894,4.5017757,4.7516575,5.001539,5.251421,5.5013027,5.813655,6.126007,6.4383593,6.7507114,7.0630636,7.223144,7.387129,7.551114,7.7111945,7.8751793,9.37447,10.87376,12.376955,13.8762455,15.375536,15.262308,15.14908,15.035853,14.92653,14.813302,13.673217,12.537036,11.400854,10.260769,9.124588,7.9259367,6.7233806,5.5247293,4.3260775,3.1235218,3.0259118,2.9243972,2.8267872,2.7252727,2.6237583,2.6510892,2.6745155,2.7018464,2.7252727,2.7486992,2.436347,2.1239948,1.8116426,1.4992905,1.1869383,1.33921,1.4875772,1.6359446,1.7882162,1.9365835,2.951728,3.9629683,4.9742084,5.989353,7.000593,7.1762915,7.348085,7.523783,7.699481,7.8751793,6.3017054,4.7243266,3.1508527,1.5734742,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.26159495,0.27330816,0.28892577,0.30063897,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.23816854,0.22645533,0.21083772,0.19912452,0.18741131,1.7491722,3.310933,4.8765984,6.4383593,8.00012,9.362757,10.725393,12.08803,13.450665,14.813302,14.13784,13.462379,12.786918,12.111456,11.435994,11.674163,11.912332,12.150499,12.388668,12.626837,12.376955,12.123169,11.873287,11.623405,11.373524,11.525795,11.674163,11.826434,11.974802,12.123169,12.587793,13.048512,13.513136,13.973856,14.438479,16.226696,18.011007,19.799223,21.58744,23.375656,25.03893,26.698303,28.361578,30.024853,31.68813,35.373886,39.063545,42.749302,46.43896,50.124718,46.77474,43.424763,40.074783,36.724808,33.374832,33.062477,32.750126,32.437775,32.125423,31.81307,28.837915,25.86276,22.887606,19.91245,16.937298,14.711788,12.486279,10.260769,8.039165,5.813655,4.9234514,4.037152,3.1508527,2.260649,1.3743496,4.037152,6.699954,9.362757,12.025558,14.688361,15.863586,17.03881,18.214037,19.389261,20.560583,17.226223,13.887959,10.549695,7.211431,3.873167,5.7980375,7.726812,9.651682,11.576552,13.501423,12.4745655,11.4516115,10.424754,9.4018,8.374943,9.901564,11.424281,12.950902,14.473619,16.00024,15.687888,15.375536,15.063184,14.750832,14.438479,12.4745655,10.510651,8.550641,6.5867267,4.6267166,5.263134,5.899552,6.5359693,7.1762915,7.812709,10.6238785,13.438952,16.250122,19.061293,21.876366,23.461554,25.050644,26.635832,28.224924,29.814016,30.099037,30.387962,30.67689,30.96191,31.250835,28.97457,26.698303,24.425941,22.149673,19.873407,16.863113,13.848915,10.838621,7.824422,4.814128,5.0132523,5.212377,5.4115014,5.610626,5.813655,6.4383593,7.0630636,7.687768,8.312472,8.937177,8.648251,8.36323,8.074304,7.7892823,7.5003567,10.237343,12.974329,15.711315,18.448301,21.189192,20.06082,18.936352,17.811884,16.687416,15.562947,15.562947,15.562947,15.562947,15.562947,15.562947,18.401447,21.236044,24.074545,26.913044,29.751545,29.251781,28.748114,28.24835,27.748587,27.248823,25.398136,23.551353,21.700668,19.849981,17.999294,16.800642,15.598087,14.399435,13.200784,11.998228,10.561408,9.124588,7.687768,6.250948,4.814128,5.8761253,6.9381227,8.00012,9.062118,10.124115,12.314485,14.50095,16.687416,18.87388,21.06425,23.114061,25.163872,27.213684,29.263494,31.313307,30.637844,29.962383,29.28692,28.61146,27.935999,27.748587,27.561176,27.373764,27.186354,26.998941,24.988174,22.973503,20.962736,18.948065,16.937298,16.164225,15.387249,14.614178,13.837202,13.06413,12.236397,11.412568,10.588739,9.761005,8.937177,13.462379,17.987581,22.512783,27.037985,31.563189,36.31094,41.0626,45.814255,50.562008,55.313667,55.598686,55.887615,56.17654,56.46156,56.75049,48.812836,40.875187,32.93754,24.999887,17.062239,15.8987255,14.739119,13.575606,12.412095,11.248583,11.974802,12.70102,13.423335,14.149553,14.875772,13.58732,12.298867,11.014318,9.725866,8.437413,7.238762,6.036206,4.8375545,3.638903,2.436347,2.77603,3.1118085,3.4514916,3.78727,4.123049,5.563773,7.000593,8.437413,9.874233,11.311053,9.749292,8.187531,6.6257706,5.0640097,3.4983444,3.0259118,2.5495746,2.0732377,1.6008049,1.1244678,1.175225,1.2259823,1.2767396,1.3235924,1.3743496,1.4133936,1.4485333,1.4875772,1.5266213,1.5617609,1.2494087,0.93705654,0.62470436,0.31235218,0.0,0.0,0.0,0.0,0.0,0.0,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,0.76135844,0.9019169,1.038571,1.175225,1.3118792,1.1869383,1.0619974,0.93705654,0.81211567,0.6871748,0.58566034,0.48805028,0.38653582,0.28892577,0.18741131,0.21083772,0.23816854,0.26159495,0.28892577,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,1.9873407,3.5998588,5.212377,6.824895,8.437413,7.363703,6.2860875,5.212377,4.138666,3.0610514,2.787743,2.514435,2.2372224,1.9639144,1.6867018,2.1864653,2.6862288,3.1859922,3.6857557,4.1894236,4.7126136,5.2358036,5.7628975,6.2860875,6.813182,5.899552,4.985922,4.0761957,3.1625657,2.2489357,2.1864653,2.1239948,2.0615244,1.999054,1.9365835,1.7257458,1.5110037,1.3001659,1.0893283,0.8745861,1.3235924,1.7765031,2.2255092,2.6745155,3.1235218,2.736986,2.35045,1.9639144,1.5734742,1.1869383,1.0893283,0.9878138,0.8862993,0.78868926,0.6871748,0.61299115,0.5388075,0.46071947,0.38653582,0.31235218,0.3631094,0.41386664,0.46071947,0.5114767,0.5622339,0.4997635,0.43729305,0.37482262,0.31235218,0.24988174,0.23816854,0.22645533,0.21083772,0.19912452,0.18741131,1.1361811,2.0888553,3.0376248,3.9863946,4.939069,5.64967,6.364176,7.0747766,7.7892823,8.499884,8.85128,9.198771,9.550168,9.901564,10.249056,10.186585,10.124115,10.061645,9.999174,9.936704,11.213444,12.486279,13.763018,15.035853,16.312593,19.100336,21.888079,24.675823,27.463566,30.251308,33.86288,37.474453,41.086025,44.7015,48.313072,44.650745,40.988415,37.326084,33.663757,30.001427,27.276154,24.55088,21.82561,19.100336,16.375063,15.836256,15.3013525,14.762545,14.223738,13.688834,14.239355,14.785972,15.336493,15.8870125,16.437534,15.976814,15.51219,15.051471,14.586847,14.126127,13.688834,13.251541,12.814248,12.376955,11.935758,11.014318,10.088976,9.163632,8.238289,7.3129454,6.551587,5.786324,5.024966,4.263607,3.4983444,3.3890212,3.2757936,3.1625657,3.049338,2.9361105,3.5608149,4.1894236,4.814128,5.4388323,6.0635366,1.2884527,1.4016805,1.5110037,1.6242313,1.737459,1.8506867,1.7023194,1.5539521,1.4055848,1.261122,1.1127546,1.0854238,1.0580931,1.0307622,1.0034313,0.97610056,1.2923572,1.6086137,1.9287747,2.2450314,2.5612879,2.8385005,3.1118085,3.3890212,3.6623292,3.9356375,4.037152,4.138666,4.2362766,4.337791,4.4393053,4.5954814,4.7516575,4.911738,5.067914,5.22409,4.728231,4.2362766,3.7404175,3.2445583,2.7486992,2.366068,1.9834363,1.6008049,1.2181735,0.8394465,1.0463798,1.2533131,1.4602464,1.6671798,1.8741131,2.069333,2.2645533,2.4597735,2.6549935,2.8502135,2.5495746,2.2489357,1.9482968,1.6515622,1.3509232,1.1557031,0.96438736,0.77307165,0.58175594,0.38653582,0.43338865,0.47633708,0.5231899,0.5661383,0.61299115,1.4914817,2.366068,3.2445583,4.123049,5.001539,5.1303844,5.2592297,5.388075,5.520825,5.64967,5.911265,6.1767645,6.4383593,6.699954,6.9615493,7.195813,7.426173,7.660437,7.890797,8.125061,9.280765,10.436467,11.588266,12.743969,13.899672,14.243259,14.590752,14.934339,15.281831,15.625418,14.204215,12.786918,11.365715,9.944512,8.52331,7.3246584,6.126007,4.9234514,3.7247996,2.5261483,2.7330816,2.9439192,3.154757,3.3655949,3.5764325,3.5725281,3.5686235,3.5686235,3.5647192,3.5608149,3.3343596,3.1039999,2.87364,2.6432803,2.4129205,2.4988174,2.5808098,2.6667068,2.7526035,2.8385005,3.8263142,4.8180323,5.805846,6.7975645,7.7892823,7.7892823,7.793187,7.793187,7.7970915,7.800996,6.239235,4.6813784,3.1196175,1.5617609,0.0,0.08589685,0.1717937,0.25378615,0.339683,0.42557985,0.5583295,0.6910792,0.8238289,0.95657855,1.0893283,0.8941081,0.698888,0.5036679,0.30844778,0.113227665,0.12884527,0.14836729,0.1639849,0.1835069,0.19912452,0.19131571,0.1796025,0.1717937,0.16008049,0.14836729,1.6320401,3.1157131,4.5993857,6.0791545,7.562827,8.925464,10.2881,11.650736,13.013372,14.376009,13.735687,13.09927,12.4628525,11.826434,11.186112,11.46723,11.748346,12.025558,12.306676,12.587793,12.552653,12.517513,12.482374,12.447234,12.412095,12.568271,12.724447,12.8767185,13.032895,13.189071,13.759113,14.329156,14.899199,15.469242,16.039284,17.882162,19.728945,21.571823,23.418604,25.261482,26.983324,28.701262,30.423103,32.14104,33.86288,37.146484,40.43399,43.71759,47.001194,50.2887,46.196888,42.10117,38.009357,33.91754,29.82573,29.849155,29.876486,29.899912,29.92334,29.95067,26.932568,23.914463,20.89636,17.878258,14.864059,12.978233,11.092407,9.20658,7.320754,5.4388323,4.872694,4.3065557,3.7443218,3.1781836,2.612045,4.8765984,7.137247,9.4018,11.66245,13.923099,15.035853,16.148607,17.261362,18.374117,19.486872,16.531239,13.571702,10.61607,7.656533,4.7009,5.997162,7.2934237,8.59359,9.889851,11.186112,10.721489,10.25296,9.784432,9.315904,8.85128,10.48332,12.119265,13.755209,15.391153,17.023193,17.003672,16.980246,16.95682,16.933393,16.91387,15.067088,13.224211,11.377428,9.530646,7.687768,7.4847393,7.28171,7.0786815,6.8756523,6.676528,9.14411,11.611692,14.079274,16.546856,19.014439,20.783133,22.555733,24.328331,26.10093,27.873528,28.27568,28.68174,29.083893,29.486046,29.888199,27.479183,25.074072,22.665054,20.256039,17.850927,15.551234,13.2554455,10.955752,8.659965,6.364176,6.168956,5.9776397,5.786324,5.591104,5.3997884,6.0205884,6.6413884,7.2582836,7.8790836,8.499884,8.265619,8.031356,7.793187,7.558923,7.3246584,10.2100115,13.095366,15.980719,18.866072,21.751425,20.076437,18.405352,16.734268,15.059279,13.388195,13.692739,13.997282,14.301826,14.606369,14.9109125,18.237463,21.564014,24.88666,28.213211,31.535856,32.94925,34.35874,35.76823,37.17772,38.587208,34.108856,29.634413,25.156063,20.677715,16.199366,15.277926,14.356487,13.431144,12.509705,11.588266,10.194394,8.804427,7.4105554,6.016684,4.6267166,5.4115014,6.196286,6.9810715,7.7658563,8.550641,10.249056,11.951375,13.64979,15.348206,17.050524,19.896833,22.743143,25.593357,28.439667,31.285975,30.161507,29.033134,27.904762,26.77639,25.651922,25.515268,25.378614,25.245865,25.109211,24.976461,23.153105,21.333654,19.514202,17.694752,15.875299,15.492668,15.110037,14.727406,14.344774,13.962143,13.091461,12.220779,11.354002,10.48332,9.612638,13.32182,17.031002,20.74409,24.453272,28.162453,32.16837,36.174286,40.1763,44.182217,48.188133,48.281837,48.375546,48.473152,48.56686,48.660564,42.585316,36.51397,30.43872,24.36347,18.28822,17.24184,16.191557,15.145176,14.098797,13.048512,13.134409,13.216402,13.298394,13.380386,13.462379,12.2793455,11.092407,9.909373,8.722435,7.5394006,6.5125427,5.4856853,4.462732,3.435874,2.4129205,2.7018464,2.9868677,3.2757936,3.5608149,3.8497405,5.1108627,6.36808,7.629202,8.890324,10.151445,8.683391,7.2192397,5.755089,4.290938,2.8267872,2.4480603,2.0732377,1.698415,1.3235924,0.94876975,1.0737107,1.1986516,1.3235924,1.4485333,1.5734742,1.5110037,1.4446288,1.3782539,1.3157835,1.2494087,0.999527,0.74964523,0.4997635,0.24988174,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.20693332,0.30844778,0.40996224,0.5114767,0.62470436,0.737932,0.8511597,0.96438736,1.0737107,0.9956226,0.92143893,0.8433509,0.76526284,0.6871748,0.6442264,0.59737355,0.5544251,0.5075723,0.46071947,0.42948425,0.39824903,0.3631094,0.3318742,0.30063897,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.10541886,0.21083772,0.31625658,0.42167544,0.5231899,1.8663043,3.2055142,4.5447245,5.883934,7.223144,6.3134184,5.4036927,4.493967,3.5842414,2.6745155,2.416825,2.1591344,1.901444,1.6437533,1.3860629,1.796025,2.2059872,2.6159496,3.0259118,3.435874,3.8458362,4.251894,4.661856,5.067914,5.473972,4.7516575,4.029343,3.3070288,2.5847144,1.8623998,1.8194515,1.7765031,1.7335546,1.6906061,1.6515622,1.4680552,1.2884527,1.1088502,0.92924774,0.74964523,1.1205635,1.4914817,1.8584955,2.2294137,2.6003318,2.2957885,1.9912452,1.6867018,1.3782539,1.0737107,0.9917182,0.9097257,0.8277333,0.74574083,0.6637484,0.58956474,0.5192855,0.44510186,0.3709182,0.30063897,0.339683,0.37872702,0.42167544,0.46071947,0.4997635,0.44900626,0.39824903,0.3513962,0.30063897,0.24988174,0.24597734,0.23816854,0.23426414,0.23035973,0.22645533,1.1674163,2.1083772,3.0532427,3.9942036,4.939069,5.704332,6.46569,7.230953,7.996216,8.761478,8.964508,9.167537,9.370565,9.573594,9.776623,9.725866,9.675109,9.6243515,9.573594,9.526741,10.994797,12.466757,13.934812,15.406772,16.874826,20.68162,24.492315,28.299107,32.1059,35.912693,43.990902,52.069107,60.143414,68.22162,76.29983,76.07337,75.85082,75.62437,75.40182,75.17536,71.618454,68.06154,64.500725,60.943813,57.386906,51.951977,46.517048,41.08212,35.647194,30.212265,28.888672,27.561176,26.237583,24.91399,23.586494,21.899792,20.21309,18.526388,16.835783,15.14908,14.586847,14.020708,13.45457,12.888432,12.326198,11.354002,10.38571,9.413514,8.445222,7.47693,6.7780423,6.083059,5.388075,4.6969957,3.998108,3.7794614,3.5608149,3.338264,3.1196175,2.900971,3.4710135,4.041056,4.6110992,5.181142,5.7511845,1.261122,1.3743496,1.4875772,1.6008049,1.7140326,1.8233559,1.6671798,1.5110037,1.3509232,1.1947471,1.038571,1.0190489,1.0034313,0.98390937,0.96829176,0.94876975,1.2220778,1.4953861,1.7686942,2.0380979,2.3114061,2.5495746,2.787743,3.0259118,3.2640803,3.4983444,3.6232853,3.7482262,3.873167,3.998108,4.123049,4.3534083,4.579864,4.806319,5.036679,5.263134,4.872694,4.482254,4.0918136,3.7013733,3.310933,2.97125,2.631567,2.2918842,1.9522011,1.6125181,1.7647898,1.9170616,2.069333,2.2216048,2.3738766,2.4402514,2.5066261,2.5690966,2.6354716,2.7018464,2.4246337,2.1513257,1.8741131,1.6008049,1.3235924,1.1400855,0.95657855,0.76916724,0.58566034,0.39824903,0.5270943,0.6559396,0.78088045,0.9097257,1.038571,1.979532,2.9243972,3.8653584,4.806319,5.7511845,5.758993,5.7707067,5.7785153,5.7902284,5.801942,6.012779,6.223617,6.4383593,6.649197,6.8639393,7.164578,7.4691215,7.7697606,8.074304,8.374943,9.183154,9.99527,10.803481,11.615597,12.423808,13.228115,14.028518,14.832824,15.633226,16.437534,14.735214,13.032895,11.330575,9.628256,7.9259367,6.7233806,5.5247293,4.3260775,3.1235218,1.9248703,2.4441557,2.9634414,3.4866312,4.0059166,4.5252023,4.493967,4.466636,4.435401,4.4041657,4.376835,4.2284675,4.0801005,3.9317331,3.7833657,3.638903,3.6584249,3.677947,3.697469,3.716991,3.736513,4.704805,5.6730967,6.6413884,7.605776,8.574067,8.406178,8.234385,8.066495,7.8947015,7.726812,6.180669,4.6345253,3.0883822,1.5461433,0.0,0.12103647,0.23816854,0.359205,0.48024148,0.60127795,0.8511597,1.1049459,1.358732,1.6086137,1.8623998,1.53443,1.2064602,0.8784905,0.5544251,0.22645533,0.21083772,0.19522011,0.1796025,0.1639849,0.14836729,0.14055848,0.13665408,0.12884527,0.12103647,0.113227665,1.5149081,2.9165885,4.318269,5.7238536,7.125534,8.488171,9.850807,11.213444,12.576079,13.938716,13.337439,12.73616,12.138786,11.537509,10.936231,11.260296,11.584361,11.904523,12.228588,12.548749,12.728352,12.911859,13.091461,13.271063,13.450665,13.610746,13.770826,13.930907,14.090988,14.251068,14.92653,15.605896,16.281357,16.960724,17.636185,19.541533,21.442978,23.344421,25.245865,27.151213,28.927717,30.70422,32.48072,34.26113,36.037632,38.919083,41.80053,44.685883,47.567333,50.44878,45.61513,40.781483,35.943928,31.110277,26.276627,26.635832,26.998941,27.362051,27.72516,28.08827,25.027218,21.966167,18.90902,15.847969,12.786918,11.240774,9.698535,8.152391,6.606249,5.0640097,4.8219366,4.575959,4.3338866,4.0918136,3.8497405,5.7121406,7.57454,9.43694,11.29934,13.16174,14.212025,15.262308,16.312593,17.362877,18.41316,15.836256,13.25935,10.67854,8.101635,5.5247293,6.196286,6.8639393,7.535496,8.203149,8.874706,8.964508,9.054309,9.14411,9.2339115,9.323712,11.06898,12.814248,14.559516,16.304783,18.05005,18.319456,18.584955,18.854359,19.119858,19.389261,17.65961,15.933866,14.204215,12.47847,10.748819,9.706344,8.663869,7.621393,6.578918,5.5364423,7.660437,9.780528,11.904523,14.028518,16.148607,18.108618,20.064724,22.020828,23.980839,25.936945,26.45623,26.971611,27.490896,28.006277,28.525562,25.983797,23.445936,20.90417,18.366308,15.824542,14.243259,12.661977,11.076789,9.495506,7.914223,7.328563,6.7429028,6.1572423,5.571582,4.985922,5.602817,6.2158084,6.832704,7.445695,8.062591,7.8790836,7.6955767,7.5159745,7.3324676,7.1489606,10.182681,13.216402,16.246218,19.279938,22.31366,20.092054,17.874353,15.652749,13.431144,11.213444,11.82253,12.431617,13.040704,13.653695,14.262781,18.073479,21.888079,25.698776,29.513376,33.324074,36.64672,39.96546,43.284203,46.60685,49.92559,42.81958,35.713566,28.61146,21.505447,14.399435,13.755209,13.110983,12.466757,11.818625,11.174399,9.82738,8.480362,7.1333427,5.786324,4.4393053,4.9468775,5.4505453,5.958118,6.46569,6.9732623,8.187531,9.4018,10.612165,11.826434,13.036799,16.683512,20.326319,23.97303,27.615837,31.262548,29.681267,28.103888,26.522604,24.941322,23.363943,23.278046,23.196054,23.114061,23.032068,22.950077,21.321941,19.693806,18.06567,16.441439,14.813302,14.821111,14.832824,14.840633,14.852346,14.864059,13.946525,13.032895,12.119265,11.20173,10.2881,13.181262,16.07833,18.97149,21.868557,24.761719,28.021894,31.28207,34.542248,37.80242,41.0626,40.96499,40.86738,40.769768,40.672157,40.574547,36.3617,32.14885,27.935999,23.723148,19.514202,18.58105,17.647898,16.714746,15.781594,14.848442,14.2901125,13.731783,13.169549,12.611219,12.0489855,10.967466,9.885946,8.800523,7.719003,6.6374836,5.786324,4.939069,4.087909,3.2367494,2.3855898,2.6237583,2.8619268,3.1000953,3.338264,3.5764325,4.657952,5.7394714,6.8209906,7.9064145,8.987934,7.621393,6.250948,4.884407,3.5178664,2.1513257,1.8741131,1.6008049,1.3235924,1.0502841,0.77307165,0.97610056,1.175225,1.3743496,1.5734742,1.7765031,1.6086137,1.4407244,1.2728351,1.1049459,0.93705654,0.74964523,0.5622339,0.37482262,0.18741131,0.0,0.0,0.0,0.0,0.0,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,0.48805028,0.57394713,0.6637484,0.74964523,0.8394465,0.80821127,0.77697605,0.74574083,0.71841,0.6871748,0.698888,0.7066968,0.71841,0.7262188,0.737932,0.6481308,0.5583295,0.46852827,0.37872702,0.28892577,0.23816854,0.18741131,0.13665408,0.08589685,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.13665408,0.26940376,0.40605783,0.5388075,0.6754616,1.7413634,2.8111696,3.8770714,4.9468775,6.012779,5.267039,4.521298,3.775557,3.0337205,2.2879796,2.0459068,1.8077383,1.5656652,1.3274968,1.0893283,1.4055848,1.7257458,2.0459068,2.366068,2.6862288,2.979059,3.2679846,3.5569105,3.8458362,4.138666,3.6037633,3.0727646,2.541766,2.0068626,1.475864,1.4524376,1.4290112,1.4055848,1.3860629,1.3626363,1.2142692,1.0659018,0.92143893,0.77307165,0.62470436,0.9136301,1.2064602,1.4953861,1.7843118,2.0732377,1.8506867,1.6281357,1.4055848,1.1869383,0.96438736,0.8980125,0.8316377,0.76916724,0.7027924,0.63641757,0.5661383,0.4958591,0.42557985,0.359205,0.28892577,0.31625658,0.3474918,0.37872702,0.40605783,0.43729305,0.39824903,0.3631094,0.3240654,0.28892577,0.24988174,0.25378615,0.25378615,0.25769055,0.26159495,0.26159495,1.1986516,2.1318035,3.06886,4.0020123,4.939069,5.755089,6.571109,7.3910336,8.207053,9.023073,9.081639,9.136301,9.190963,9.245625,9.300286,9.261242,9.226103,9.187058,9.151918,9.112875,10.77615,12.44333,14.106606,15.773785,17.437061,22.266806,27.092648,31.918488,36.748234,41.574074,54.11892,66.65986,79.204704,91.74564,104.28658,107.49991,110.713234,113.92655,117.13597,120.3493,115.96075,111.56829,107.17975,102.7912,98.39874,88.067696,77.73274,67.401695,57.07065,46.735695,43.53799,40.33638,37.138676,33.937065,30.739359,27.826675,24.91399,22.001307,19.088623,16.175938,15.480955,14.789876,14.098797,13.403813,12.712734,11.697589,10.682445,9.6673,8.652155,7.6370106,7.008402,6.3836975,5.755089,5.12648,4.5017757,4.173806,3.8458362,3.5178664,3.1898966,2.8619268,3.377308,3.892689,4.40807,4.9234514,5.4388323,1.2376955,1.3509232,1.4641509,1.5734742,1.6867018,1.7999294,1.6320401,1.4641509,1.2962615,1.1283722,0.96438736,0.95657855,0.94876975,0.94096094,0.93315214,0.92534333,1.1517987,1.3782539,1.6086137,1.8350691,2.0615244,2.260649,2.463678,2.6628022,2.8619268,3.0610514,3.213323,3.3616903,3.513962,3.6623292,3.8106966,4.1113358,4.40807,4.704805,5.001539,5.298274,5.0132523,4.728231,4.4432096,4.1581883,3.873167,3.5764325,3.279698,2.9829633,2.6862288,2.3855898,2.4831998,2.5808098,2.67842,2.77603,2.87364,2.8111696,2.7447948,2.67842,2.6159496,2.5495746,2.2996929,2.0498111,1.7999294,1.5500476,1.3001659,1.1205635,0.94486535,0.76916724,0.58956474,0.41386664,0.62079996,0.8316377,1.0424755,1.2533131,1.4641509,2.4714866,3.4788225,4.4861584,5.493494,6.5008297,6.3915067,6.278279,6.168956,6.0596323,5.950309,6.114294,6.2743745,6.4383593,6.5984397,6.7624245,7.1333427,7.5081654,7.8790836,8.253906,8.624825,9.089449,9.554072,10.018696,10.48332,10.951848,12.209065,13.470188,14.73131,15.988527,17.24965,15.266212,13.2788725,11.295436,9.308095,7.3246584,6.126007,4.9234514,3.7247996,2.5261483,1.3235924,2.15523,2.9868677,3.814601,4.646239,5.473972,5.4193106,5.3607445,5.3021784,5.2436123,5.1889505,5.1225758,5.056201,4.9937305,4.927356,4.860981,4.8180323,4.7711797,4.728231,4.6813784,4.6384296,5.5832953,6.5281606,7.473026,8.4178915,9.362757,9.019169,8.675582,8.335898,7.9923115,7.648724,6.1181984,4.591577,3.0610514,1.5305257,0.0,0.15617609,0.30844778,0.46462387,0.62079996,0.77307165,1.1478943,1.5188124,1.893635,2.2645533,2.639376,2.1786566,1.717937,1.2572175,0.79649806,0.3357786,0.28892577,0.24207294,0.19522011,0.14836729,0.10151446,0.093705654,0.08980125,0.08589685,0.078088045,0.07418364,1.397776,2.7213683,4.041056,5.364649,6.688241,8.050878,9.413514,10.77615,12.138786,13.501423,12.939189,12.376955,11.810817,11.248583,10.686349,11.053363,11.416472,11.783486,12.146595,12.513609,12.907954,13.302299,13.696643,14.090988,14.489237,14.653222,14.817206,14.981192,15.14908,15.313066,16.09785,16.882635,17.66742,18.452206,19.23699,21.197,23.15701,25.11702,27.07703,29.037039,30.872108,32.707176,34.542248,36.377316,38.212383,40.69168,43.170975,45.654175,48.133472,50.612766,45.033375,39.45789,33.878498,28.303013,22.723621,23.426414,24.125301,24.82419,25.523077,26.22587,23.12187,20.021774,16.917774,13.813775,10.71368,9.507219,8.300759,7.098203,5.891743,4.689187,4.7672753,4.8492675,4.927356,5.009348,5.087436,6.551587,8.011833,9.475985,10.936231,12.400381,13.388195,14.376009,15.363823,16.351637,17.335546,15.141272,12.943093,10.744915,8.546737,6.348558,6.3915067,6.434455,6.477403,6.520352,6.5633,7.211431,7.8556576,8.503788,9.151918,9.80005,11.654641,13.509232,15.363823,17.218414,19.07691,19.631334,20.189665,20.747993,21.306324,21.860748,20.252134,18.64352,17.031002,15.422389,13.813775,11.931853,10.046027,8.164105,6.282183,4.4002614,6.1767645,7.9532676,9.733675,11.510178,13.286681,15.430198,17.573715,19.713327,21.856844,24.00036,24.632874,25.265387,25.8979,26.530413,27.162926,24.48841,21.8178,19.143284,16.472673,13.798158,12.93138,12.064603,11.197825,10.331048,9.464272,8.484266,7.5081654,6.5281606,5.55206,4.575959,5.185046,5.794133,6.4032197,7.016211,7.6252975,7.4964523,7.363703,7.2348576,7.1060123,6.9732623,10.155351,13.333533,16.515621,19.693806,22.875893,20.107672,17.33945,14.571229,11.803008,9.0386915,9.952321,10.865952,11.783486,12.697116,13.610746,17.913397,22.212145,26.510891,30.813543,35.11229,40.34419,45.57218,50.80408,56.032078,61.263977,51.5303,41.796627,32.06295,22.333181,12.599506,12.232492,11.8654785,11.498465,11.131451,10.764437,9.460366,8.156297,6.8561306,5.55206,4.251894,4.478349,4.7087092,4.939069,5.169429,5.3997884,6.126007,6.8483214,7.57454,8.300759,9.023073,13.466284,17.909492,22.352703,26.795912,31.239122,29.20493,27.170734,25.140446,23.106253,21.075964,21.044727,21.013493,20.986162,20.954927,20.92369,19.490776,18.053955,16.62104,15.18422,13.751305,14.153459,14.555612,14.957765,15.359919,15.762072,14.801589,13.841106,12.880623,11.924045,10.963562,13.040704,15.12175,17.202797,19.283842,21.360985,23.879324,26.393759,28.908194,31.42263,33.937065,33.64814,33.359215,33.066383,32.77746,32.488533,30.13808,27.78763,25.437181,23.086731,20.73628,19.92026,19.10424,18.284315,17.468296,16.64837,15.445815,14.243259,13.040704,11.838148,10.6355915,9.655587,8.675582,7.6955767,6.715572,5.735567,5.0640097,4.388548,3.7130866,3.0376248,2.3621633,2.5495746,2.736986,2.9243972,3.1118085,3.2992198,4.2050414,5.1108627,6.016684,6.918601,7.824422,6.5554914,5.2865605,4.0137253,2.7447948,1.475864,1.3001659,1.1244678,0.94876975,0.77307165,0.60127795,0.8745861,1.1517987,1.4251068,1.698415,1.9756275,1.7062237,1.43682,1.1635119,0.8941081,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.113227665,0.1717937,0.23035973,0.28892577,0.3513962,0.41386664,0.47633708,0.5388075,0.60127795,0.61689556,0.63641757,0.6520352,0.6715572,0.6871748,0.75354964,0.8160201,0.8823949,0.94876975,1.0112402,0.8667773,0.71841,0.5700427,0.42167544,0.27330816,0.22645533,0.1756981,0.12494087,0.07418364,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.1639849,0.3318742,0.4958591,0.659844,0.8238289,1.620327,2.416825,3.2094188,4.0059166,4.7985106,4.220659,3.638903,3.0610514,2.4792955,1.901444,1.678893,1.456342,1.2337911,1.0112402,0.78868926,1.0190489,1.2494087,1.475864,1.7062237,1.9365835,2.1083772,2.2840753,2.455869,2.6276627,2.7994564,2.455869,2.1161861,1.7725986,1.4290112,1.0893283,1.0854238,1.0815194,1.0815194,1.077615,1.0737107,0.96048295,0.8433509,0.7301232,0.61689556,0.4997635,0.7106012,0.92143893,1.1283722,1.33921,1.5500476,1.4094892,1.2689307,1.1283722,0.9917182,0.8511597,0.80430686,0.75354964,0.7066968,0.659844,0.61299115,0.5466163,0.47633708,0.40996224,0.3435874,0.27330816,0.29673457,0.31625658,0.3357786,0.3553006,0.37482262,0.3513962,0.3240654,0.30063897,0.27330816,0.24988174,0.26159495,0.26940376,0.28111696,0.28892577,0.30063897,1.2259823,2.15523,3.084478,4.009821,4.939069,5.805846,6.676528,7.5472097,8.4178915,9.288573,9.194867,9.101162,9.01136,8.917655,8.823949,8.800523,8.773191,8.749765,8.726339,8.699008,10.561408,12.419904,14.278399,16.140799,17.999294,23.84809,29.696884,35.541775,41.390568,47.239365,64.24694,81.25452,98.26209,115.26576,132.27724,138.92644,145.57564,152.22484,158.87404,165.52713,160.30304,155.07895,149.85876,144.63467,139.41449,124.18342,108.95235,93.721275,78.4941,63.26303,58.187305,53.111584,48.035862,42.964043,37.88832,33.749653,29.610987,25.476225,21.337559,17.198893,16.378967,15.559043,14.739119,13.919194,13.09927,12.041177,10.979179,9.921086,8.859089,7.800996,7.238762,6.6804323,6.1181984,5.559869,5.001539,4.564246,4.1308575,3.6935644,3.260176,2.8267872,3.2836022,3.7443218,4.2050414,4.6657605,5.12648,1.2142692,1.3235924,1.43682,1.5500476,1.6632754,1.7765031,1.5969005,1.4212024,1.2415999,1.0659018,0.8862993,0.8902037,0.8941081,0.8941081,0.8980125,0.9019169,1.0815194,1.2650263,1.4485333,1.6281357,1.8116426,1.9756275,2.135708,2.2996929,2.463678,2.6237583,2.7994564,2.9751544,3.1508527,3.3265507,3.4983444,3.8692627,4.2362766,4.60329,4.970304,5.337318,5.1577153,4.9781127,4.7985106,4.618908,4.4393053,4.181615,3.9278288,3.6740425,3.416352,3.1625657,3.2055142,3.2484627,3.2914112,3.3343596,3.3734035,3.1781836,2.9868677,2.7916477,2.5964274,2.4012074,2.174752,1.9482968,1.7257458,1.4992905,1.2767396,1.1049459,0.93315214,0.76526284,0.59346914,0.42557985,0.71841,1.0112402,1.3040704,1.5969005,1.8858263,2.959537,4.0332475,5.1069584,6.1767645,7.250475,7.0201154,6.7897553,6.559396,6.329036,6.098676,6.211904,6.3251314,6.4383593,6.551587,6.66091,7.1060123,7.5472097,7.988407,8.433509,8.874706,8.995743,9.116779,9.2339115,9.354948,9.475985,11.193921,12.911859,14.625891,16.343828,18.061766,15.793307,13.528754,11.260296,8.991838,6.7233806,5.5247293,4.3260775,3.1235218,1.9248703,0.7262188,1.8663043,3.0063896,4.1464753,5.2865605,6.426646,6.3407493,6.2548523,6.168956,6.083059,6.001066,6.016684,6.036206,6.0518236,6.0713453,6.086963,5.9776397,5.8683167,5.758993,5.645766,5.5364423,6.461786,7.3832245,8.304664,9.226103,10.151445,9.636065,9.120684,8.605303,8.089922,7.57454,6.0596323,4.5447245,3.0298162,1.5149081,0.0,0.19131571,0.37872702,0.5700427,0.76135844,0.94876975,1.4407244,1.9365835,2.4285383,2.920493,3.4124475,2.8189783,2.2294137,1.6359446,1.0424755,0.44900626,0.3709182,0.28892577,0.21083772,0.12884527,0.05075723,0.046852827,0.046852827,0.042948425,0.039044023,0.039044023,1.2806439,2.522244,3.7638438,5.009348,6.250948,7.6135845,8.976221,10.338858,11.701493,13.06413,12.537036,12.013845,11.486752,10.963562,10.436467,10.84643,11.252487,11.6585455,12.068507,12.4745655,13.083652,13.696643,14.30573,14.914817,15.523903,15.695697,15.863586,16.03538,16.20327,16.375063,17.26917,18.159374,19.053482,19.943687,20.837795,22.85637,24.871042,26.889618,28.908194,30.926771,32.8165,34.710136,36.60377,38.493504,40.38714,42.46428,44.54142,46.618565,48.695705,50.776752,44.455524,38.134296,31.81307,25.495747,19.174519,20.21309,21.251661,22.286327,23.3249,24.36347,21.216522,18.073479,14.92653,11.783486,8.636538,7.773665,6.9068875,6.044015,5.1772375,4.3143644,4.716518,5.1186714,5.520825,5.9229784,6.3251314,7.387129,8.449126,9.511124,10.573121,11.639023,12.564366,13.4858055,14.411149,15.336493,16.261835,14.446288,12.626837,10.81129,8.991838,7.1762915,6.590631,6.0049706,5.4193106,4.83365,4.251894,5.45445,6.66091,7.8634663,9.069926,10.276386,12.240301,14.204215,16.168129,18.135948,20.099863,20.947119,21.794373,22.641628,23.488884,24.33614,22.844658,21.353176,19.861694,18.366308,16.874826,14.153459,11.428185,8.706817,5.985449,3.2640803,4.6930914,6.126007,7.558923,8.991838,10.424754,12.751778,15.078801,17.405825,19.736753,22.063778,22.809519,23.559164,24.304905,25.050644,25.80029,22.99693,20.189665,17.386303,14.579038,11.775677,11.623405,11.471134,11.318862,11.166591,11.014318,9.643873,8.273428,6.902983,5.532538,4.1620927,4.7672753,5.3724575,5.9776397,6.5828223,7.1880045,7.1099167,7.0318284,6.9537406,6.8756523,6.801469,10.128019,13.45457,16.78112,20.111576,23.438128,20.12329,16.808453,13.493614,10.178777,6.8639393,8.082112,9.304191,10.522364,11.744442,12.962616,17.749413,22.53621,27.326912,32.11371,36.900505,44.041656,51.178905,58.320057,65.461205,72.59846,60.241024,47.879684,35.51835,23.160913,10.799577,10.709775,10.619974,10.530173,10.4403715,10.350571,9.093353,7.8361354,6.578918,5.3217,4.0605783,4.0137253,3.9668727,3.9200199,3.873167,3.8263142,4.0605783,4.298747,4.5369153,4.775084,5.0132523,10.25296,15.492668,20.732376,25.972084,31.211792,28.728592,26.241488,23.758287,21.271183,18.787983,18.81141,18.830933,18.854359,18.877785,18.90121,17.655706,16.414106,15.172507,13.930907,12.689307,13.481901,14.278399,15.070992,15.867491,16.663988,15.656653,14.653222,13.645885,12.642454,11.639023,12.90405,14.169076,15.434102,16.69913,17.964155,19.73285,21.501543,23.274141,25.042835,26.811531,26.33129,25.847143,25.366901,24.882755,24.39861,23.910559,23.426414,22.938364,22.450314,21.962263,21.25947,20.556679,19.853886,19.151093,18.448301,16.605423,14.75864,12.915763,11.06898,9.226103,8.347612,7.4691215,6.590631,5.716045,4.8375545,4.337791,3.8380275,3.338264,2.8385005,2.338737,2.475391,2.612045,2.7486992,2.8892577,3.0259118,3.7521305,4.478349,5.2084727,5.9346914,6.66091,5.4895897,4.318269,3.1430438,1.9717231,0.80040246,0.7262188,0.6481308,0.57394713,0.4997635,0.42557985,0.77307165,1.1244678,1.475864,1.8233559,2.174752,1.8038338,1.4290112,1.0580931,0.6832704,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.0,0.0,0.0,0.0,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.21083772,0.24988174,0.28892577,0.3240654,0.3631094,0.42557985,0.49195468,0.5583295,0.62079996,0.6871748,0.80821127,0.92924774,1.0463798,1.1674163,1.2884527,1.0815194,0.8784905,0.6715572,0.46852827,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.19522011,0.39044023,0.58566034,0.78088045,0.97610056,1.4992905,2.018576,2.541766,3.0649557,3.5881457,3.174279,2.7565079,2.3426414,1.9287747,1.5110037,1.3079748,1.1010414,0.8980125,0.6910792,0.48805028,0.62860876,0.76916724,0.9058213,1.0463798,1.1869383,1.2415999,1.2962615,1.3509232,1.4055848,1.4641509,1.3118792,1.1557031,1.0034313,0.8511597,0.698888,0.71841,0.7340276,0.75354964,0.76916724,0.78868926,0.7066968,0.62079996,0.5388075,0.45681506,0.37482262,0.5036679,0.63641757,0.76526284,0.8941081,1.0268579,0.96829176,0.9097257,0.8511597,0.79649806,0.737932,0.7066968,0.679366,0.6481308,0.61689556,0.58566034,0.5231899,0.45681506,0.39434463,0.3279698,0.26159495,0.27330816,0.28111696,0.29283017,0.30063897,0.31235218,0.30063897,0.28892577,0.27330816,0.26159495,0.24988174,0.26940376,0.28502136,0.30063897,0.32016098,0.3357786,1.2572175,2.1786566,3.096191,4.01763,4.939069,5.860508,6.7819467,7.703386,8.628729,9.550168,9.308095,9.069926,8.831758,8.589685,8.351517,8.335898,8.324185,8.312472,8.300759,8.289046,10.342762,12.396477,14.454097,16.507812,18.56153,25.429373,32.297215,39.16506,46.0329,52.900745,74.37496,95.849174,117.31948,138.78978,160.26399,170.34908,180.43805,190.52702,200.61209,210.70107,204.64534,198.58961,192.53389,186.48206,180.42633,160.29523,140.16805,120.04085,99.91756,79.78646,72.836624,65.88679,58.93695,51.987118,45.03728,39.676537,34.311886,28.951143,23.586494,18.22575,17.27698,16.32821,15.383345,14.434575,13.4858055,12.380859,11.275913,10.170968,9.066022,7.9610763,7.4691215,6.9771667,6.4852123,5.9932575,5.5013027,4.958591,4.415879,3.873167,3.330455,2.787743,3.193801,3.5959544,4.0020123,4.40807,4.814128,1.1869383,1.3001659,1.4133936,1.5266213,1.6359446,1.7491722,1.5617609,1.3743496,1.1869383,0.999527,0.81211567,0.8238289,0.8394465,0.8511597,0.8628729,0.8745861,1.0112402,1.1517987,1.2884527,1.4251068,1.5617609,1.6867018,1.8116426,1.9365835,2.0615244,2.1864653,2.3855898,2.5886188,2.787743,2.9868677,3.1859922,3.6232853,4.0605783,4.5017757,4.939069,5.376362,5.298274,5.22409,5.1499066,5.0757227,5.001539,4.786797,4.575959,4.3612175,4.1503797,3.9356375,3.9239242,3.912211,3.900498,3.8887846,3.873167,3.5491016,3.2250361,2.900971,2.5769055,2.2489357,2.0498111,1.8506867,1.6515622,1.4485333,1.2494087,1.0893283,0.92534333,0.76135844,0.60127795,0.43729305,0.81211567,1.1869383,1.5617609,1.9365835,2.3114061,3.4514916,4.5876727,5.7238536,6.8639393,8.00012,7.648724,7.3012323,6.949836,6.5984397,6.250948,6.3134184,6.375889,6.4383593,6.5008297,6.5633,7.0747766,7.5862536,8.101635,8.6131115,9.124588,8.898132,8.675582,8.449126,8.226576,8.00012,10.174872,12.349625,14.524376,16.69913,18.87388,16.324306,13.774731,11.225157,8.675582,6.126007,4.9234514,3.7247996,2.5261483,1.3235924,0.12494087,1.5734742,3.0259118,4.474445,5.9268827,7.375416,7.262188,7.1489606,7.0357327,6.9264097,6.813182,6.910792,7.012306,7.113821,7.211431,7.3129454,7.137247,6.9615493,6.785851,6.6140575,6.4383593,7.336372,8.238289,9.136301,10.0382185,10.936231,10.249056,9.561881,8.874706,8.187531,7.5003567,6.001066,4.5017757,2.998581,1.4992905,0.0,0.22645533,0.44900626,0.6754616,0.9019169,1.1244678,1.737459,2.35045,2.9634414,3.5764325,4.1894236,3.4632049,2.736986,2.0107672,1.2884527,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.0,0.0,0.0,0.0,0.0,1.1635119,2.3231194,3.4866312,4.650143,5.813655,7.1762915,8.538928,9.901564,11.2642,12.626837,12.138786,11.650736,11.162686,10.674636,10.186585,10.6355915,11.088503,11.537509,11.986515,12.439425,13.263254,14.087084,14.9109125,15.738646,16.562475,16.738173,16.91387,17.085665,17.261362,17.437061,18.436588,19.436115,20.435642,21.439074,22.4386,24.511837,26.58898,28.662216,30.739359,32.812595,34.760895,36.713093,38.661392,40.613594,42.56189,44.236877,45.911865,47.586853,49.261845,50.936832,43.873768,36.81461,29.751545,22.688482,15.625418,16.999767,18.374117,19.748466,21.12672,22.50107,19.311174,16.125181,12.939189,9.749292,6.5633,6.036206,5.5130157,4.985922,4.462732,3.9356375,4.661856,5.388075,6.114294,6.8366084,7.562827,8.226576,8.886419,9.550168,10.213917,10.87376,11.736633,12.599506,13.462379,14.325252,15.188125,13.751305,12.314485,10.87376,9.43694,8.00012,6.785851,5.575486,4.3612175,3.1508527,1.9365835,3.7013733,5.462259,7.223144,8.987934,10.748819,12.825961,14.899199,16.976341,19.049578,21.12672,22.262901,23.399082,24.539167,25.67535,26.811531,25.437181,24.062832,22.688482,21.314133,19.935879,16.375063,12.814248,9.249529,5.688714,2.1239948,3.213323,4.298747,5.388075,6.473499,7.562827,10.073358,12.587793,15.098324,17.612759,20.12329,20.986162,21.849035,22.711908,23.574781,24.437654,21.501543,18.56153,15.625418,12.689307,9.749292,10.311526,10.87376,11.435994,11.998228,12.564366,10.799577,9.0386915,7.2739015,5.5130157,3.7482262,4.349504,4.950782,5.548156,6.1494336,6.7507114,6.7233806,6.699954,6.676528,6.649197,6.6257706,10.100689,13.575606,17.050524,20.525442,24.00036,20.138906,16.273548,12.412095,8.550641,4.689187,6.211904,7.7385254,9.261242,10.787864,12.31058,17.589333,22.86418,28.139027,33.413876,38.68872,47.73913,56.785625,65.83603,74.88644,83.93684,68.94784,53.96274,38.973743,23.988647,8.999647,9.187058,9.37447,9.561881,9.749292,9.936704,8.726339,7.5120697,6.3017054,5.087436,3.873167,3.5491016,3.2250361,2.900971,2.5769055,2.2489357,1.999054,1.7491722,1.4992905,1.2494087,0.999527,7.039637,13.075843,19.11205,25.148254,31.188366,28.24835,25.31224,22.37613,19.436115,16.500004,16.574188,16.64837,16.72646,16.800642,16.874826,15.824542,14.774258,13.723974,12.67369,11.623405,12.814248,14.001186,15.188125,16.375063,17.562002,16.511717,15.461433,14.411149,13.360865,12.31058,12.763491,13.212498,13.661504,14.114414,14.56342,15.586374,16.613232,17.636185,18.663042,19.685997,19.010534,18.338978,17.663515,16.988054,16.312593,17.686943,19.061293,20.435642,21.813896,23.188246,22.59868,22.01302,21.423454,20.837795,20.24823,17.761126,15.274021,12.786918,10.299813,7.812709,7.0357327,6.262661,5.4856853,4.7126136,3.9356375,3.611572,3.2875066,2.9634414,2.639376,2.3114061,2.4012074,2.4871042,2.5769055,2.6628022,2.7486992,3.2992198,3.8497405,4.4002614,4.950782,5.5013027,4.423688,3.349977,2.2762666,1.1986516,0.12494087,0.14836729,0.1756981,0.19912452,0.22645533,0.24988174,0.6754616,1.1010414,1.5266213,1.9482968,2.3738766,1.901444,1.4251068,0.94876975,0.47633708,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.23816854,0.3513962,0.46071947,0.57394713,0.6871748,0.8628729,1.038571,1.2142692,1.3860629,1.5617609,1.3001659,1.038571,0.77307165,0.5114767,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22645533,0.44900626,0.6754616,0.9019169,1.1244678,1.3743496,1.6242313,1.8741131,2.1239948,2.3738766,2.1239948,1.8741131,1.6242313,1.3743496,1.1244678,0.93705654,0.74964523,0.5622339,0.37482262,0.18741131,0.23816854,0.28892577,0.3357786,0.38653582,0.43729305,0.37482262,0.31235218,0.24988174,0.18741131,0.12494087,0.1639849,0.19912452,0.23816854,0.27330816,0.31235218,0.3513962,0.38653582,0.42557985,0.46071947,0.4997635,0.44900626,0.39824903,0.3513962,0.30063897,0.24988174,0.30063897,0.3513962,0.39824903,0.44900626,0.4997635,0.5231899,0.5505207,0.57394713,0.60127795,0.62470436,0.61299115,0.60127795,0.58566034,0.57394713,0.5622339,0.4997635,0.43729305,0.37482262,0.31235218,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.27330816,0.30063897,0.3240654,0.3513962,0.37482262,1.2884527,2.1981785,3.1118085,4.025439,4.939069,5.911265,6.8873653,7.8634663,8.835662,9.811763,9.425227,9.0386915,8.648251,8.261715,7.8751793,7.8751793,7.8751793,7.8751793,7.8751793,7.8751793,10.124115,12.373051,14.625891,16.874826,19.123762,27.014559,34.90145,42.788345,50.675236,58.56213,84.502975,110.43992,136.37686,162.3099,188.25075,201.7756,215.30046,228.8253,242.35016,65535.0,248.98764,242.10027,235.2129,228.32555,221.43817,196.41095,171.38374,146.36043,121.33711,96.3138,87.48594,78.661995,69.83804,61.014095,52.18624,45.599514,39.012787,32.42606,25.839334,19.248703,18.174992,17.101282,16.023666,14.949956,13.8762455,12.724447,11.576552,10.424754,9.276859,8.125061,7.699481,7.2739015,6.8483214,6.426646,6.001066,5.349031,4.7009,4.0488653,3.4007344,2.7486992,3.1000953,3.4514916,3.7989833,4.1503797,4.5017757,1.0737107,1.1674163,1.261122,1.3509232,1.4446288,1.5383345,1.397776,1.2572175,1.116659,0.97610056,0.8394465,0.8511597,0.8667773,0.8823949,0.8980125,0.9136301,1.0268579,1.1439898,1.2572175,1.3743496,1.4875772,1.6125181,1.737459,1.8623998,1.9873407,2.1122816,2.2918842,2.4675822,2.6432803,2.822883,2.998581,3.39683,3.795079,4.193328,4.591577,4.985922,4.950782,4.9156423,4.884407,4.8492675,4.814128,4.6384296,4.466636,4.2948427,4.123049,3.951255,3.9239242,3.8965936,3.8692627,3.8419318,3.8106966,3.7638438,3.716991,3.6701381,3.6232853,3.5764325,3.377308,3.1781836,2.9829633,2.7838387,2.5886188,2.3855898,2.1864653,1.9873407,1.7882162,1.5890918,1.9834363,2.377781,2.7721257,3.1664703,3.5608149,4.290938,5.017157,5.743376,6.473499,7.1997175,6.9537406,6.7116675,6.46569,6.2197127,5.9737353,5.9932575,6.016684,6.036206,6.055728,6.0752497,6.461786,6.8483214,7.238762,7.6252975,8.011833,7.882988,7.7541428,7.621393,7.492548,7.363703,9.331521,11.303245,13.271063,15.242786,17.210606,15.242786,13.271063,11.303245,9.331521,7.363703,6.196286,5.0327744,3.8692627,2.7018464,1.5383345,3.0805733,4.6228123,6.165051,7.70729,9.249529,8.952794,8.65606,8.359325,8.058686,7.7619514,7.605776,7.445695,7.289519,7.1333427,6.9732623,7.1880045,7.3988423,7.6135845,7.824422,8.039165,8.320281,8.601398,8.886419,9.167537,9.448653,8.991838,8.531119,8.070399,7.60968,7.1489606,6.133816,5.114767,4.095718,3.0805733,2.0615244,1.9482968,1.8389735,1.7257458,1.6125181,1.4992905,2.0068626,2.5105307,3.0141985,3.521771,4.025439,3.4436827,2.8658314,2.2840753,1.7062237,1.1244678,1.2767396,1.4290112,1.5812829,1.7335546,1.8858263,1.5188124,1.1478943,0.77697605,0.40605783,0.039044023,1.261122,2.4831998,3.7052777,4.927356,6.1494336,7.2582836,8.371038,9.479889,10.588739,11.701493,11.053363,10.409137,9.76491,9.120684,8.476458,8.8083315,9.14411,9.479889,9.815667,10.151445,11.221252,12.291059,13.360865,14.430671,15.500477,15.926057,16.351637,16.773312,17.198893,17.624472,18.87388,20.119385,21.368793,22.614298,23.863707,25.468416,27.073126,28.677835,30.282543,31.887253,33.85898,35.8307,37.806328,39.77805,41.749775,43.33496,44.920147,46.505337,48.090523,49.67571,43.026512,36.373413,29.724215,23.075018,16.42582,17.273075,18.124235,18.975395,19.826555,20.67381,18.061766,15.449719,12.837675,10.22563,7.6135845,6.735094,5.8566036,4.9781127,4.1035266,3.2250361,4.3455997,5.4700675,6.590631,7.715099,8.835662,8.831758,8.827853,8.823949,8.81614,8.812236,9.63216,10.452085,11.272009,12.091934,12.911859,11.998228,11.080693,10.167064,9.253433,8.335898,7.687768,7.0357327,6.387602,5.735567,5.087436,6.086963,7.08649,8.086017,9.089449,10.088976,11.85767,13.626364,15.398962,17.167656,18.936352,20.19357,21.450787,22.711908,23.969126,25.226343,24.792953,24.359566,23.926178,23.496693,23.063305,19.170614,15.277926,11.385237,7.492548,3.5998588,4.3026514,5.0054436,5.708236,6.4110284,7.113821,9.077735,11.04165,13.009468,14.973383,16.937298,17.796265,18.659138,19.518106,20.377075,21.236044,18.877785,16.515621,14.157363,11.799104,9.43694,10.046027,10.6590185,11.268105,11.877192,12.486279,10.889378,9.288573,7.687768,6.086963,4.4861584,5.1460023,5.805846,6.46569,7.1294384,7.7892823,7.47693,7.1606736,6.8483214,6.5359693,6.223617,9.499411,12.775204,16.050997,19.326792,22.59868,19.482967,16.36335,13.247637,10.128019,7.012306,7.8790836,8.745861,9.616543,10.48332,11.350098,16.87873,22.411268,27.939903,33.468536,39.001076,45.591705,52.18624,58.77687,65.37141,71.962036,59.514805,47.071472,34.628143,22.18091,9.737579,9.897659,10.05774,10.217821,10.377901,10.537982,9.780528,9.026978,8.273428,7.5159745,6.7624245,5.794133,4.8219366,3.853645,2.8814487,1.9131571,1.737459,1.5617609,1.3860629,1.2142692,1.038571,5.9737353,10.912805,15.851873,20.787037,25.726107,23.937891,22.149673,20.361458,18.573242,16.788929,16.191557,15.594183,14.996809,14.395531,13.798158,13.673217,13.548276,13.423335,13.298394,13.173453,14.184693,15.195933,16.20327,17.21451,18.22575,17.10909,15.996336,14.879677,13.766922,12.650263,12.455043,12.259823,12.064603,11.869383,11.674163,13.028991,14.379913,15.730837,17.085665,18.436588,17.519053,16.601519,15.683984,14.766449,13.848915,15.730837,17.608854,19.490776,21.368793,23.250715,22.21605,21.181383,20.146715,19.108145,18.073479,15.969006,13.864532,11.760059,9.655587,7.551114,6.9654536,6.379793,5.794133,5.2084727,4.6267166,4.2284675,3.8341231,3.4397783,3.0454338,2.6510892,2.639376,2.631567,2.619854,2.6081407,2.6003318,3.1039999,3.6037633,4.1074314,4.6110992,5.1108627,4.1191444,3.1274261,2.135708,1.1439898,0.14836729,0.23035973,0.30844778,0.39044023,0.46852827,0.5505207,0.8355421,1.1205635,1.4055848,1.6906061,1.9756275,1.5812829,1.1869383,0.78868926,0.39434463,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.10932326,0.14055848,0.1717937,0.20693332,0.23816854,0.30844778,0.38263142,0.45681506,0.5270943,0.60127795,0.7301232,0.8589685,0.9917182,1.1205635,1.2494087,1.1205635,0.9917182,0.8589685,0.7301232,0.60127795,0.48024148,0.359205,0.23816854,0.12103647,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.3318742,0.5270943,0.7223144,0.91753453,1.1127546,1.2767396,1.43682,1.6008049,1.7608855,1.9248703,1.7296503,1.53443,1.33921,1.1439898,0.94876975,0.80430686,0.6559396,0.5075723,0.359205,0.21083772,0.24597734,0.28111696,0.31625658,0.3513962,0.38653582,0.3357786,0.28111696,0.23035973,0.1756981,0.12494087,0.15227169,0.1796025,0.20693332,0.23426414,0.26159495,0.30063897,0.3435874,0.38263142,0.42167544,0.46071947,0.41386664,0.3670138,0.32016098,0.27330816,0.22645533,0.30844778,0.39044023,0.47243267,0.5544251,0.63641757,0.63641757,0.63641757,0.63641757,0.63641757,0.63641757,0.61299115,0.58566034,0.5622339,0.5388075,0.5114767,0.46071947,0.41386664,0.3631094,0.31235218,0.26159495,0.25769055,0.25378615,0.24597734,0.24207294,0.23816854,0.23426414,0.23426414,0.23035973,0.22645533,0.22645533,0.24207294,0.26159495,0.27721256,0.29673457,0.31235218,1.2494087,2.182561,3.1157131,4.0527697,4.985922,5.794133,6.602344,7.4105554,8.218767,9.023073,8.577971,8.128965,7.6838636,7.2348576,6.785851,6.9068875,7.0240197,7.141152,7.2582836,7.375416,10.108498,12.841579,15.570756,18.303837,21.036919,27.459661,33.882404,40.305145,46.727886,53.150627,74.29687,95.447014,116.59326,137.7395,158.88574,169.34564,179.80553,190.26152,200.71751,211.17351,209.28377,207.39404,205.5043,203.61458,201.72485,180.89876,160.07268,139.2505,118.42442,97.59834,93.22541,88.856384,84.48346,80.11053,75.737595,68.96736,62.19713,55.426895,48.656662,41.88643,37.263615,32.636898,28.014086,23.38737,18.760653,16.863113,14.96167,13.06413,11.162686,9.261242,8.65606,8.046973,7.4417906,6.832704,6.223617,5.579391,4.9351645,4.290938,3.6467118,2.998581,3.213323,3.4241607,3.638903,3.8497405,4.0605783,0.96438736,1.0346665,1.1088502,1.1791295,1.2533131,1.3235924,1.2337911,1.1400855,1.0463798,0.95657855,0.8628729,0.8784905,0.8980125,0.9136301,0.93315214,0.94876975,1.0424755,1.1361811,1.2259823,1.319688,1.4133936,1.5383345,1.6632754,1.7882162,1.9131571,2.0380979,2.194274,2.3465457,2.5027218,2.6588979,2.8111696,3.1703746,3.5256753,3.8848803,4.2440853,4.5993857,4.60329,4.6110992,4.6150036,4.618908,4.6267166,4.493967,4.3612175,4.2284675,4.095718,3.9629683,3.9200199,3.8770714,3.8341231,3.7911747,3.7482262,3.978586,4.2089458,4.4393053,4.6696653,4.900025,4.704805,4.5095844,4.3143644,4.1191444,3.9239242,3.6857557,3.4514916,3.213323,2.9751544,2.736986,3.1508527,3.5686235,3.9824903,4.396357,4.814128,5.1303844,5.446641,5.7668023,6.083059,6.3993154,6.2587566,6.1181984,5.9815445,5.840986,5.700427,5.677001,5.6535745,5.6340523,5.610626,5.5871997,5.8487945,6.114294,6.375889,6.6374836,6.899079,6.8639393,6.8287997,6.79366,6.75852,6.7233806,8.488171,10.256865,12.021654,13.786445,15.551234,14.161267,12.771299,11.381332,9.991365,8.601398,7.4691215,6.3407493,5.2084727,4.0801005,2.951728,4.5837684,6.2197127,7.8556576,9.491602,11.123642,10.6434,10.159255,9.679013,9.194867,8.710721,8.296855,7.882988,7.4691215,7.0513506,6.6374836,7.238762,7.8361354,8.437413,9.0386915,9.636065,9.304191,8.968412,8.632633,8.296855,7.9610763,7.7307167,7.4964523,7.266093,7.0318284,6.801469,6.266566,5.7316628,5.196759,4.661856,4.126953,3.6740425,3.2250361,2.77603,2.3231194,1.8741131,2.2723622,2.6706111,3.06886,3.4632049,3.8614538,3.4280653,2.9907722,2.5573835,2.1239948,1.6867018,2.1044729,2.522244,2.9400148,3.357786,3.775557,3.0337205,2.2957885,1.5539521,0.8160201,0.07418364,1.358732,2.639376,3.9239242,5.2045684,6.4891167,7.3441806,8.203149,9.058213,9.917182,10.77615,9.971844,9.171441,8.367134,7.5667315,6.7624245,6.9810715,7.2036223,7.422269,7.6409154,7.8634663,9.17925,10.491129,11.806912,13.122696,14.438479,15.113941,15.789403,16.46096,17.136421,17.811884,19.30727,20.802654,22.29804,23.793427,25.288813,26.42109,27.557272,28.693453,29.82573,30.96191,32.957058,34.95221,36.947357,38.94251,40.937656,42.433044,43.92843,45.423817,46.9192,48.410683,42.175354,35.93612,29.700788,23.461554,17.226223,17.550287,17.874353,18.19842,18.526388,18.850454,16.812357,14.774258,12.73616,10.698062,8.663869,7.433982,6.2040954,4.9742084,3.7443218,2.514435,4.0332475,5.55206,7.0708723,8.59359,10.112402,9.440845,8.769287,8.093826,7.422269,6.7507114,7.5276875,8.304664,9.081639,9.858616,10.6355915,10.2451515,9.850807,9.460366,9.066022,8.675582,8.58578,8.499884,8.413987,8.324185,8.238289,8.476458,8.710721,8.94889,9.187058,9.425227,10.889378,12.353529,13.821584,15.285735,16.749886,18.12814,19.506393,20.880743,22.258997,23.63725,24.148727,24.6563,25.167776,25.679255,26.186827,21.966167,17.741604,13.520945,9.296382,5.0757227,5.3919797,5.708236,6.028397,6.3446536,6.66091,8.078208,9.495506,10.916709,12.334006,13.751305,14.606369,15.465338,16.324306,17.17937,18.038338,16.254026,14.473619,12.689307,10.9089,9.124588,9.784432,10.4403715,11.096312,11.756155,12.412095,10.975275,9.538455,8.101635,6.66091,5.22409,5.9464045,6.6648145,7.3832245,8.105539,8.823949,8.226576,7.6252975,7.0240197,6.426646,5.825368,8.902037,11.974802,15.051471,18.124235,21.200905,18.827028,16.453152,14.0831785,11.709302,9.339331,9.546264,9.757101,9.967939,10.178777,10.38571,16.172033,21.958359,27.740778,33.527103,39.313427,43.44819,47.58295,51.717712,55.852474,59.987236,50.08567,40.18411,30.278639,20.377075,10.475512,10.608261,10.741011,10.87376,11.00651,11.139259,10.838621,10.541886,10.2451515,9.948417,9.651682,8.03526,6.4188375,4.806319,3.1898966,1.5734742,1.475864,1.3743496,1.2767396,1.175225,1.0737107,4.911738,8.749765,12.587793,16.42582,20.263847,19.623526,18.987108,18.35069,17.714273,17.073952,15.80502,14.53609,13.263254,11.994324,10.725393,11.525795,12.326198,13.1266,13.923099,14.723501,15.559043,16.39068,17.222319,18.053955,18.885593,17.706465,16.527334,15.348206,14.169076,12.986042,12.146595,11.307149,10.467703,9.628256,8.78881,10.467703,12.146595,13.829392,15.5082855,17.18718,16.02757,14.867964,13.708356,12.548749,11.389141,13.770826,16.156416,18.542006,20.927597,23.313187,21.829514,20.34584,18.866072,17.382399,15.8987255,14.176885,12.455043,10.733202,9.01136,7.2856145,6.89127,6.4969254,6.1025805,5.708236,5.3138914,4.8492675,4.380739,3.9161155,3.4514916,2.9868677,2.8814487,2.7721257,2.6667068,2.5573835,2.4480603,2.9048753,3.3616903,3.814601,4.271416,4.7243266,3.814601,2.9048753,1.9951496,1.0854238,0.1756981,0.30844778,0.44510186,0.58175594,0.7145056,0.8511597,0.9956226,1.1400855,1.2845483,1.4290112,1.5734742,1.261122,0.94486535,0.62860876,0.31625658,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.14055848,0.19131571,0.24597734,0.29673457,0.3513962,0.38263142,0.41386664,0.44900626,0.48024148,0.5114767,0.59737355,0.6832704,0.76916724,0.8511597,0.93705654,0.94096094,0.94096094,0.94486535,0.94876975,0.94876975,0.76135844,0.5700427,0.37872702,0.19131571,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05466163,0.10932326,0.1639849,0.21864653,0.27330816,0.44119745,0.60518235,0.76916724,0.93315214,1.1010414,1.175225,1.2494087,1.3235924,1.4016805,1.475864,1.3353056,1.1947471,1.0541886,0.9136301,0.77307165,0.6676528,0.5583295,0.45291066,0.3435874,0.23816854,0.25769055,0.27721256,0.29673457,0.31625658,0.3357786,0.29673457,0.25378615,0.21083772,0.1678893,0.12494087,0.14055848,0.16008049,0.1756981,0.19522011,0.21083772,0.25378615,0.29673457,0.339683,0.38263142,0.42557985,0.37872702,0.3357786,0.28892577,0.24597734,0.19912452,0.31625658,0.42948425,0.5466163,0.659844,0.77307165,0.74964523,0.7262188,0.698888,0.6754616,0.6481308,0.61299115,0.57394713,0.5388075,0.4997635,0.46071947,0.42557985,0.38653582,0.3513962,0.31235218,0.27330816,0.26549935,0.25378615,0.24597734,0.23426414,0.22645533,0.21864653,0.21474212,0.21083772,0.20693332,0.19912452,0.21083772,0.21864653,0.23035973,0.23816854,0.24988174,1.2064602,2.1630387,3.1235218,4.0801005,5.036679,5.677001,6.3173227,6.957645,7.5979667,8.238289,7.7307167,7.223144,6.715572,6.2079997,5.700427,5.9346914,6.168956,6.4032197,6.6413884,6.8756523,10.088976,13.306203,16.519526,19.736753,22.950077,27.908667,32.86726,37.821945,42.780537,47.73913,64.094666,80.45411,96.809654,113.16519,129.52464,136.91568,144.3067,151.69383,159.08487,166.4759,169.5838,172.69171,175.79572,178.90361,182.01152,165.38658,148.76163,132.13669,115.51174,98.886795,98.96879,99.046875,99.12887,99.206955,99.28895,92.33521,85.38147,78.43163,71.47789,64.524155,56.348335,48.172516,40.000603,31.824783,23.648964,21.00178,18.35069,15.699601,13.048512,10.401327,9.608734,8.8200445,8.031356,7.238762,6.4500723,5.8097506,5.169429,4.5291066,3.8887846,3.2484627,3.3265507,3.4007344,3.474918,3.5491016,3.6232853,0.8511597,0.9019169,0.95657855,1.0073358,1.0580931,1.1127546,1.0659018,1.0229534,0.97610056,0.93315214,0.8862993,0.9058213,0.92924774,0.94876975,0.96829176,0.9878138,1.0580931,1.1283722,1.1986516,1.2689307,1.33921,1.4641509,1.5890918,1.7140326,1.8389735,1.9639144,2.096664,2.2294137,2.358259,2.4910088,2.6237583,2.9439192,3.260176,3.5764325,3.8965936,4.21285,4.2557983,4.3026514,4.3455997,4.3924527,4.4393053,4.3455997,4.251894,4.1581883,4.068387,3.9746814,3.9161155,3.8614538,3.802888,3.7443218,3.6857557,4.193328,4.7009,5.2084727,5.716045,6.223617,6.0323014,5.840986,5.645766,5.45445,5.263134,4.985922,4.7126136,4.4393053,4.1620927,3.8887846,4.322173,4.755562,5.192855,5.6262436,6.0635366,5.969831,5.8761253,5.786324,5.6926184,5.5989127,5.563773,5.5286336,5.493494,5.4583545,5.423215,5.3607445,5.2943697,5.2318993,5.165524,5.099149,5.2358036,5.376362,5.5130157,5.64967,5.786324,5.8487945,5.9073606,5.9659266,6.028397,6.086963,7.648724,9.20658,10.768341,12.326198,13.887959,13.075843,12.267632,11.45942,10.647305,9.839094,8.741957,7.648724,6.551587,5.4583545,4.3612175,6.0908675,7.816613,9.546264,11.272009,13.001659,12.334006,11.666354,10.998701,10.331048,9.663396,8.991838,8.316377,7.6448197,6.9732623,6.3017054,7.2856145,8.273428,9.261242,10.249056,11.23687,10.284196,9.331521,8.378847,7.426173,6.473499,6.4695945,6.46569,6.461786,6.453977,6.4500723,6.3993154,6.3446536,6.2938967,6.239235,6.1884775,5.3997884,4.6110992,3.8263142,3.0376248,2.2489357,2.541766,2.8306916,3.1196175,3.408543,3.7013733,3.408543,3.1196175,2.8306916,2.541766,2.2489357,2.9322062,3.6154766,4.298747,4.9781127,5.661383,4.552533,3.4436827,2.330928,1.2220778,0.113227665,1.456342,2.795552,4.138666,5.481781,6.824895,7.4300776,8.03526,8.640442,9.245625,9.850807,8.890324,7.929841,6.969358,6.008875,5.0483923,5.153811,5.2592297,5.364649,5.4700675,5.575486,7.1333427,8.695104,10.256865,11.814721,13.376482,14.301826,15.223265,16.148607,17.073952,17.999294,19.740658,21.485926,23.22729,24.968653,26.71392,27.377668,28.041416,28.70907,29.372818,30.036566,32.05514,34.07372,36.08839,38.106964,40.12554,41.531128,42.93671,44.33839,45.743977,47.149563,41.324192,35.498825,29.673458,23.84809,18.026625,17.823597,17.624472,17.425346,17.226223,17.023193,15.562947,14.098797,12.63855,11.174399,9.714153,8.128965,6.547683,4.9663997,3.3812122,1.7999294,3.716991,5.6340523,7.551114,9.468176,11.389141,10.046027,8.706817,7.367607,6.028397,4.689187,5.423215,6.1572423,6.89127,7.629202,8.36323,8.492075,8.62092,8.75367,8.882515,9.01136,9.487698,9.964035,10.436467,10.912805,11.389141,10.862047,10.338858,9.811763,9.288573,8.761478,9.921086,11.080693,12.244205,13.403813,14.56342,16.058807,17.558098,19.053482,20.552773,22.048159,23.500597,24.953035,26.409376,27.861814,29.314253,24.761719,20.209187,15.656653,11.10412,6.551587,6.481308,6.4149327,6.348558,6.278279,6.211904,7.082586,7.9532676,8.823949,9.690726,10.561408,11.416472,12.271536,13.1266,13.981665,14.836729,13.634172,12.427712,11.221252,10.018696,8.812236,9.518932,10.221725,10.928422,11.631214,12.337912,11.061172,9.788337,8.511597,7.238762,5.9620223,6.7429028,7.523783,8.300759,9.081639,9.86252,8.976221,8.086017,7.1997175,6.3134184,5.423215,8.300759,11.174399,14.051944,16.925583,19.799223,18.171087,16.546856,14.918721,13.2905855,11.66245,11.213444,10.768341,10.319335,9.874233,9.425227,15.465338,21.505447,27.545557,33.585667,39.62578,41.300766,42.97966,44.658554,46.33354,48.012436,40.652637,33.29284,25.93304,18.573242,11.213444,11.318862,11.424281,11.525795,11.631214,11.736633,11.896713,12.056794,12.216875,12.376955,12.537036,10.276386,8.015738,5.758993,3.4983444,1.2376955,1.2142692,1.1869383,1.1635119,1.1361811,1.1127546,3.8497405,6.5867267,9.323712,12.0606985,14.801589,15.313066,15.824542,16.33602,16.8514,17.362877,15.418485,13.477997,11.533605,9.593117,7.648724,9.37447,11.100216,12.825961,14.551707,16.273548,16.92949,17.585428,18.241367,18.893402,19.549341,18.303837,17.058334,15.816733,14.571229,13.325725,11.838148,10.354475,8.870802,7.3832245,5.899552,7.9064145,9.913278,11.924045,13.930907,15.93777,14.53609,13.134409,11.728825,10.327144,8.925464,11.814721,14.703979,17.593237,20.486399,23.375656,21.442978,19.514202,17.585428,15.656653,13.723974,12.384764,11.045554,9.706344,8.36323,7.0240197,6.8209906,6.6140575,6.4110284,6.2040954,6.001066,5.466163,4.93126,4.396357,3.8614538,3.3265507,3.1196175,2.9165885,2.7096553,2.5066261,2.2996929,2.7057507,3.1157131,3.521771,3.9317331,4.337791,3.5100577,2.6823244,1.8545911,1.0268579,0.19912452,0.39044023,0.58175594,0.76916724,0.96048295,1.1517987,1.1557031,1.1596074,1.1635119,1.1713207,1.175225,0.94096094,0.7066968,0.46852827,0.23426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.1717937,0.24597734,0.31625658,0.39044023,0.46071947,0.45681506,0.44900626,0.44119745,0.43338865,0.42557985,0.46462387,0.5036679,0.5466163,0.58566034,0.62470436,0.76135844,0.8941081,1.0307622,1.1635119,1.3001659,1.038571,0.78088045,0.5192855,0.26159495,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08199245,0.1639849,0.24597734,0.3318742,0.41386664,0.5466163,0.6832704,0.8160201,0.95267415,1.0893283,1.0737107,1.0619974,1.0502841,1.038571,1.0268579,0.94096094,0.8550641,0.76916724,0.6832704,0.60127795,0.5309987,0.46462387,0.39824903,0.3318742,0.26159495,0.26940376,0.27330816,0.27721256,0.28111696,0.28892577,0.25378615,0.22255093,0.19131571,0.15617609,0.12494087,0.13274968,0.14055848,0.14836729,0.15617609,0.1639849,0.20693332,0.25378615,0.29673457,0.3435874,0.38653582,0.3435874,0.30063897,0.26159495,0.21864653,0.1756981,0.3240654,0.46852827,0.61689556,0.76526284,0.9136301,0.8628729,0.81211567,0.76135844,0.7106012,0.6637484,0.61299115,0.5622339,0.5114767,0.46071947,0.41386664,0.38653582,0.3631094,0.3357786,0.31235218,0.28892577,0.27330816,0.25769055,0.24207294,0.22645533,0.21083772,0.20693332,0.19912452,0.19131571,0.1835069,0.1756981,0.1756981,0.1796025,0.1835069,0.1835069,0.18741131,1.1674163,2.1474214,3.1274261,4.1074314,5.087436,5.559869,6.0323014,6.504734,6.9771667,7.4495993,6.883461,6.3134184,5.74728,5.181142,4.6110992,4.9663997,5.3177958,5.6691923,6.0205884,6.375889,10.073358,13.770826,17.468296,21.165764,24.863234,28.35377,31.84821,35.338745,38.833183,42.32372,53.892464,65.461205,77.02605,88.594795,100.163536,104.48571,108.807884,113.13006,117.45223,121.7744,129.87994,137.98547,146.09102,154.19266,162.29819,149.87439,137.44667,125.022865,112.59906,100.17525,104.70826,109.24127,113.774284,118.30339,122.8364,115.70306,108.56581,101.432465,94.299126,87.16187,75.43696,63.712036,51.987118,40.262196,28.537275,25.136541,21.735807,18.338978,14.938243,11.537509,10.565312,9.593117,8.62092,7.648724,6.676528,6.04011,5.4036927,4.7711797,4.134762,3.4983444,3.435874,3.3734035,3.310933,3.2484627,3.1859922,0.737932,0.76916724,0.80430686,0.8355421,0.8667773,0.9019169,0.9019169,0.9058213,0.9058213,0.9097257,0.9136301,0.93315214,0.95657855,0.98000497,1.0034313,1.0268579,1.0737107,1.1205635,1.1674163,1.2142692,1.261122,1.3860629,1.5110037,1.6359446,1.7608855,1.8858263,1.999054,2.1083772,2.2177005,2.3270237,2.436347,2.7135596,2.9907722,3.2718892,3.5491016,3.8263142,3.9083066,3.9942036,4.0801005,4.165997,4.251894,4.1972322,4.1464753,4.0918136,4.041056,3.9863946,3.9161155,3.8419318,3.7716527,3.697469,3.6232853,4.40807,5.196759,5.9815445,6.7663293,7.551114,7.3597984,7.168483,6.9810715,6.7897553,6.5984397,6.2860875,5.9737353,5.661383,5.349031,5.036679,5.493494,5.9464045,6.4032197,6.8561306,7.3129454,6.8092775,6.3056097,5.805846,5.3021784,4.7985106,4.8687897,4.939069,5.009348,5.0796275,5.1499066,5.040583,4.9351645,4.825841,4.7204223,4.6110992,4.6267166,4.6384296,4.650143,4.661856,4.6735697,4.829746,4.985922,5.138193,5.2943697,5.4505453,6.805373,8.160201,9.515028,10.869856,12.224684,11.994324,11.763964,11.533605,11.303245,11.076789,10.0147915,8.956698,7.8947015,6.8366084,5.774611,7.5940623,9.413514,11.23687,13.056321,14.875772,14.020708,13.169549,12.318389,11.4633255,10.612165,9.682918,8.75367,7.824422,6.89127,5.9620223,7.336372,8.710721,10.088976,11.4633255,12.837675,11.268105,9.698535,8.128965,6.559396,4.985922,5.2084727,5.4310236,5.6535745,5.8761253,6.098676,6.5281606,6.9615493,7.3910336,7.8205175,8.250002,7.125534,6.001066,4.8765984,3.7482262,2.6237583,2.8072653,2.9907722,3.174279,3.3538816,3.5373883,3.3929255,3.2484627,3.1039999,2.9556324,2.8111696,3.7599394,4.7087092,5.6535745,6.602344,7.551114,6.0713453,4.591577,3.1118085,1.6281357,0.14836729,1.5539521,2.9556324,4.357313,5.758993,7.1606736,7.5159745,7.8673706,8.218767,8.574067,8.925464,7.8088045,6.688241,5.571582,4.454923,3.338264,3.3265507,3.3187418,3.3070288,3.2992198,3.2875066,5.0913405,6.899079,8.702912,10.506746,12.31058,13.4858055,14.661031,15.836256,17.01148,18.186707,20.177952,22.169195,24.156536,26.147781,28.139027,28.334248,28.525562,28.720783,28.916002,29.111223,31.153225,33.191322,35.233326,37.271423,39.313427,40.62921,41.94109,43.256874,44.572655,45.88844,40.476936,35.06153,29.65003,24.23853,18.823124,18.10081,17.37459,16.64837,15.926057,15.199838,14.313539,13.423335,12.537036,11.650736,10.764437,8.827853,6.89127,4.958591,3.0220075,1.0893283,3.4007344,5.716045,8.031356,10.346666,12.661977,10.655114,8.648251,6.6413884,4.630621,2.6237583,3.3187418,4.009821,4.7009,5.395884,6.086963,6.7389984,7.3910336,8.046973,8.699008,9.351044,10.38571,11.424281,12.4628525,13.501423,14.53609,13.251541,11.963089,10.674636,9.386183,8.101635,8.956698,9.811763,10.666827,11.521891,12.376955,13.993378,15.6098,17.226223,18.84655,20.462973,22.85637,25.253674,27.647072,30.044374,32.437775,27.553368,22.672863,17.788456,12.907954,8.023546,7.570636,7.1216297,6.6687193,6.2158084,5.7628975,6.083059,6.407124,6.7311897,7.0513506,7.375416,8.226576,9.081639,9.932799,10.783959,11.639023,11.010414,10.381805,9.753197,9.128492,8.499884,9.253433,10.003078,10.756628,11.510178,12.263727,11.150972,10.0382185,8.925464,7.812709,6.699954,7.5394006,8.378847,9.218294,10.061645,10.901091,9.725866,8.550641,7.375416,6.2001905,5.024966,7.699481,10.373997,13.048512,15.726933,18.401447,17.519053,16.636658,15.754263,14.871868,13.985569,12.880623,11.775677,10.670732,9.565785,8.460839,14.75864,21.052536,27.346434,33.644234,39.93813,39.15725,38.37637,37.599392,36.818512,36.037632,31.2196,26.401567,21.583536,16.765503,11.951375,12.025558,12.103647,12.181735,12.259823,12.337912,12.954806,13.571702,14.188598,14.809398,15.426293,12.521418,9.616543,6.7116675,3.8067923,0.9019169,0.94876975,0.999527,1.0502841,1.1010414,1.1517987,2.787743,4.423688,6.0635366,7.699481,9.339331,10.998701,12.661977,14.325252,15.988527,17.651802,15.035853,12.419904,9.803954,7.191909,4.575959,7.2270484,9.874233,12.525322,15.176412,17.823597,18.303837,18.780174,19.256512,19.736753,20.21309,18.90121,17.593237,16.281357,14.973383,13.661504,11.533605,9.4018,7.2739015,5.142098,3.0141985,5.349031,7.6838636,10.018696,12.353529,14.688361,13.040704,11.39695,9.753197,8.105539,6.461786,9.858616,13.251541,16.64837,20.041296,23.438128,21.060347,18.682566,16.304783,13.927003,11.549222,10.592644,9.636065,8.675582,7.719003,6.7624245,6.746807,6.7311897,6.715572,6.703859,6.688241,6.083059,5.477876,4.872694,4.267512,3.6623292,3.3616903,3.057147,2.7565079,2.4519646,2.1513257,2.5105307,2.8697357,3.2289407,3.5881457,3.951255,3.2055142,2.4597735,1.7140326,0.96829176,0.22645533,0.46852827,0.7145056,0.96048295,1.2064602,1.4485333,1.3157835,1.1791295,1.0463798,0.9097257,0.77307165,0.62079996,0.46462387,0.30844778,0.15617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.20693332,0.29673457,0.39044023,0.48414588,0.57394713,0.5270943,0.48024148,0.43338865,0.38653582,0.3357786,0.3318742,0.3279698,0.3240654,0.31625658,0.31235218,0.58175594,0.8472553,1.116659,1.3821584,1.6515622,1.319688,0.9917182,0.659844,0.3318742,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10932326,0.21864653,0.3318742,0.44119745,0.5505207,0.6559396,0.76135844,0.8667773,0.96829176,1.0737107,0.97610056,0.8745861,0.77307165,0.6754616,0.57394713,0.5466163,0.5153811,0.48414588,0.45681506,0.42557985,0.39824903,0.3709182,0.3435874,0.31625658,0.28892577,0.27721256,0.26940376,0.25769055,0.24597734,0.23816854,0.21474212,0.19131571,0.1717937,0.14836729,0.12494087,0.12103647,0.12103647,0.11713207,0.113227665,0.113227665,0.16008049,0.20693332,0.25378615,0.30063897,0.3513962,0.30844778,0.26940376,0.23035973,0.19131571,0.14836729,0.3318742,0.5114767,0.6910792,0.8706817,1.0502841,0.97610056,0.9019169,0.8238289,0.74964523,0.6754616,0.61299115,0.5505207,0.48805028,0.42557985,0.3631094,0.3513962,0.3357786,0.3240654,0.31235218,0.30063897,0.28111696,0.26159495,0.23816854,0.21864653,0.19912452,0.19131571,0.1796025,0.1717937,0.16008049,0.14836729,0.14446288,0.14055848,0.13665408,0.12884527,0.12494087,1.1283722,2.1318035,3.1313305,4.134762,5.138193,5.4427366,5.74728,6.0518236,6.356367,6.66091,6.036206,5.407597,4.7789884,4.154284,3.5256753,3.9942036,4.466636,4.9351645,5.4036927,5.8761253,10.053836,14.235451,18.417065,22.594776,26.77639,28.802776,30.82916,32.85945,34.885834,36.91222,43.69026,50.468304,57.246346,64.020485,70.79852,72.05574,73.30906,74.56628,75.81959,77.076805,90.17998,103.28315,116.38242,129.4856,142.58878,134.3622,126.13562,117.91295,109.68637,101.4637,110.44773,119.43176,128.41579,137.40372,146.38776,139.0709,131.75015,124.4333,117.11645,109.7996,94.52558,79.24765,63.973633,48.699608,33.425587,29.275208,25.124828,20.97445,16.82407,12.67369,11.517986,10.366188,9.2104845,8.054782,6.899079,6.27047,5.6418614,5.009348,4.380739,3.7482262,3.5491016,3.349977,3.1508527,2.951728,2.7486992,0.62470436,0.63641757,0.6481308,0.6637484,0.6754616,0.6871748,0.737932,0.78868926,0.8394465,0.8862993,0.93705654,0.96438736,0.9878138,1.0112402,1.038571,1.0619974,1.0893283,1.1127546,1.1361811,1.1635119,1.1869383,1.3118792,1.43682,1.5617609,1.6867018,1.8116426,1.901444,1.9873407,2.0732377,2.1630387,2.2489357,2.4871042,2.7252727,2.9634414,3.2016098,3.435874,3.5608149,3.6857557,3.8106966,3.9356375,4.0605783,4.0488653,4.037152,4.025439,4.0137253,3.998108,3.912211,3.8263142,3.736513,3.6506162,3.5608149,4.6267166,5.688714,6.7507114,7.812709,8.874706,8.687295,8.499884,8.312472,8.125061,7.9376497,7.5862536,7.238762,6.8873653,6.5359693,6.1884775,6.66091,7.137247,7.6135845,8.086017,8.562354,7.648724,6.7389984,5.825368,4.911738,3.998108,4.173806,4.349504,4.5252023,4.7009,4.8765984,4.7243266,4.575959,4.423688,4.2753205,4.123049,4.0137253,3.900498,3.78727,3.6740425,3.5608149,3.8106966,4.0605783,4.3143644,4.564246,4.814128,5.9620223,7.113821,8.261715,9.413514,10.561408,10.912805,11.2642,11.611692,11.963089,12.31058,11.287627,10.260769,9.237816,8.210958,7.1880045,9.101162,11.014318,12.923572,14.836729,16.749886,15.711315,14.676648,13.638077,12.599506,11.560935,10.373997,9.187058,8.00012,6.813182,5.6262436,7.387129,9.148014,10.912805,12.67369,14.438479,12.24811,10.061645,7.8751793,5.688714,3.4983444,3.951255,4.4002614,4.8492675,5.298274,5.7511845,6.66091,7.57454,8.488171,9.4018,10.311526,8.85128,7.387129,5.9268827,4.462732,2.998581,3.076669,3.1508527,3.2250361,3.2992198,3.3734035,3.3734035,3.3734035,3.3734035,3.3734035,3.3734035,4.5876727,5.7980375,7.012306,8.226576,9.43694,7.5862536,5.7394714,3.8887846,2.0380979,0.18741131,1.6515622,3.1118085,4.575959,6.036206,7.5003567,7.601871,7.699481,7.800996,7.898606,8.00012,6.7233806,5.4505453,4.173806,2.900971,1.6242313,1.4992905,1.3743496,1.2494087,1.1244678,0.999527,3.049338,5.099149,7.1489606,9.198771,11.248583,12.67369,14.098797,15.523903,16.94901,18.374117,20.61134,22.848562,25.085785,27.326912,29.564135,29.28692,29.013613,28.7364,28.463093,28.18588,30.251308,32.31283,34.37436,36.435883,38.501312,39.72339,40.94937,42.175354,43.401337,44.623413,39.62578,34.62424,29.626604,24.625065,19.623526,18.374117,17.124708,15.875299,14.625891,13.376482,13.06413,12.751778,12.439425,12.123169,11.810817,9.526741,7.238762,4.950782,2.6628022,0.37482262,3.0883822,5.7980375,8.511597,11.225157,13.938716,11.2642,8.58578,5.911265,3.2367494,0.5622339,1.2142692,1.8623998,2.514435,3.1625657,3.8106966,4.985922,6.1611466,7.336372,8.511597,9.686822,11.287627,12.888432,14.489237,16.086138,17.686943,15.637131,13.58732,11.537509,9.487698,7.437886,7.988407,8.538928,9.089449,9.636065,10.186585,11.924045,13.661504,15.398962,17.136421,18.87388,22.212145,25.550407,28.888672,32.226936,35.561295,30.348919,25.136541,19.924164,14.711788,9.499411,8.663869,7.824422,6.98888,6.1494336,5.3138914,5.087436,4.860981,4.6384296,4.4119744,4.1894236,5.036679,5.8878384,6.7389984,7.5862536,8.437413,8.386656,8.335898,8.289046,8.238289,8.187531,8.987934,9.788337,10.588739,11.389141,12.185639,11.23687,10.2881,9.339331,8.386656,7.437886,8.335898,9.237816,10.135828,11.037745,11.935758,10.475512,9.01136,7.551114,6.086963,4.6267166,7.098203,9.573594,12.0489855,14.524376,16.999767,16.863113,16.72646,16.585901,16.449247,16.312593,14.551707,12.786918,11.0260315,9.261242,7.5003567,14.051944,20.599627,27.151213,33.698895,40.250484,37.013733,33.776985,30.53633,27.29958,24.062832,21.786564,19.514202,17.237936,14.96167,12.689307,12.73616,12.786918,12.837675,12.888432,12.939189,14.012899,15.086611,16.164225,17.237936,18.311647,14.762545,11.213444,7.6643414,4.1113358,0.5622339,0.6871748,0.81211567,0.93705654,1.0619974,1.1869383,1.7257458,2.260649,2.7994564,3.338264,3.873167,6.688241,9.499411,12.314485,15.125654,17.936825,14.649317,11.361811,8.074304,4.786797,1.4992905,5.0757227,8.648251,12.224684,15.801116,19.373644,19.674282,19.974922,20.27556,20.5762,20.876839,19.498585,18.124235,16.749886,15.375536,14.001186,11.225157,8.449126,5.6730967,2.900971,0.12494087,2.787743,5.4505453,8.113348,10.77615,13.438952,11.549222,9.663396,7.773665,5.8878384,3.998108,7.898606,11.799104,15.699601,19.6001,23.500597,20.67381,17.850927,15.024139,12.201257,9.37447,8.800523,8.226576,7.648724,7.0747766,6.5008297,6.676528,6.8483214,7.0240197,7.1997175,7.375416,6.699954,6.0244927,5.349031,4.6735697,3.998108,3.5998588,3.2016098,2.7994564,2.4012074,1.999054,2.3114061,2.6237583,2.9361105,3.2484627,3.5608149,2.900971,2.2372224,1.5734742,0.9136301,0.24988174,0.5505207,0.8511597,1.1517987,1.4485333,1.7491722,1.475864,1.1986516,0.92534333,0.6481308,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.23816854,0.3513962,0.46071947,0.57394713,0.6871748,0.60127795,0.5114767,0.42557985,0.3357786,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.39824903,0.80040246,1.1986516,1.6008049,1.999054,1.6008049,1.1986516,0.80040246,0.39824903,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13665408,0.27330816,0.41386664,0.5505207,0.6871748,0.76135844,0.8394465,0.9136301,0.9878138,1.0619974,0.8745861,0.6871748,0.4997635,0.31235218,0.12494087,0.14836729,0.1756981,0.19912452,0.22645533,0.24988174,0.26159495,0.27330816,0.28892577,0.30063897,0.31235218,0.28892577,0.26159495,0.23816854,0.21083772,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.113227665,0.1639849,0.21083772,0.26159495,0.31235218,0.27330816,0.23816854,0.19912452,0.1639849,0.12494087,0.3357786,0.5505207,0.76135844,0.97610056,1.1869383,1.0893283,0.9878138,0.8862993,0.78868926,0.6871748,0.61299115,0.5388075,0.46071947,0.38653582,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.28892577,0.26159495,0.23816854,0.21083772,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,1.0893283,2.1122816,3.1391394,4.1620927,5.1889505,5.3256044,5.462259,5.5989127,5.735567,5.8761253,5.1889505,4.5017757,3.8106966,3.1235218,2.436347,3.0259118,3.611572,4.2011366,4.786797,5.376362,10.0382185,14.700074,19.36193,24.023787,28.685644,29.251781,29.814016,30.37625,30.938484,31.500717,33.48806,35.4754,37.462738,39.45008,41.43742,39.62578,37.814137,35.99859,34.186947,32.375305,50.476112,68.57692,86.67383,104.774635,122.87544,118.850006,114.82457,110.799126,106.77369,102.74825,116.1872,129.62616,143.0612,156.50015,169.9391,162.43875,154.9384,147.43803,139.93768,132.43732,113.6103,94.78327,75.960144,57.137024,38.3139,33.413876,28.51385,23.613825,18.7138,13.813775,12.4745655,11.139259,9.80005,8.460839,7.125534,6.5008297,5.8761253,5.251421,4.6267166,3.998108,3.6623292,3.3265507,2.9868677,2.6510892,2.3114061,0.62470436,0.62860876,0.63641757,0.64032197,0.6442264,0.6481308,0.6910792,0.7340276,0.77697605,0.8199245,0.8628729,0.8862993,0.9136301,0.93705654,0.96438736,0.9878138,1.0268579,1.0619974,1.1010414,1.1361811,1.175225,1.2884527,1.4016805,1.5110037,1.6242313,1.737459,1.8350691,1.9326792,2.0302892,2.1278992,2.2255092,2.4831998,2.7408905,2.998581,3.2562714,3.513962,3.5842414,3.6506162,3.7208953,3.7911747,3.8614538,3.8575494,3.853645,3.8458362,3.8419318,3.8380275,3.8770714,3.9161155,3.959064,3.998108,4.037152,4.911738,5.786324,6.66091,7.5394006,8.413987,8.207053,8.0040245,7.7970915,7.5940623,7.387129,7.043542,6.703859,6.3602715,6.016684,5.6730967,6.184573,6.6960497,7.2036223,7.715099,8.226576,7.5003567,6.774138,6.0518236,5.3256044,4.5993857,4.950782,5.3060827,5.657479,6.008875,6.364176,5.9659266,5.5676775,5.169429,4.7711797,4.376835,4.138666,3.9044023,3.6701381,3.435874,3.2016098,3.4007344,3.6037633,3.8067923,4.009821,4.21285,5.376362,6.5437784,7.70729,8.870802,10.0382185,10.455989,10.87376,11.291532,11.709302,12.123169,10.963562,9.80005,8.636538,7.47693,6.3134184,7.8205175,9.327617,10.834716,12.341816,13.848915,13.228115,12.603411,11.982611,11.361811,10.737106,9.772718,8.8083315,7.843944,6.8756523,5.911265,7.3519893,8.792714,10.2334385,11.674163,13.110983,11.420377,9.725866,8.03526,6.3407493,4.650143,5.1108627,5.571582,6.028397,6.4891167,6.949836,7.531592,8.109444,8.691199,9.269051,9.850807,8.726339,7.605776,6.481308,5.3607445,4.2362766,4.0332475,3.8263142,3.6232853,3.416352,3.213323,3.6935644,4.173806,4.6540475,5.134289,5.610626,6.1299114,6.649197,7.164578,7.6838636,8.1992445,6.703859,5.2045684,3.7091823,2.2098918,0.7106012,2.05762,3.4007344,4.747753,6.0908675,7.437886,7.6643414,7.890797,8.121157,8.347612,8.574067,7.60968,6.6452928,5.6809053,4.716518,3.7482262,3.7287042,3.7091823,3.68966,3.6701381,3.6506162,5.3841705,7.1216297,8.855185,10.588739,12.326198,13.634172,14.938243,16.246218,17.554192,18.862167,21.450787,24.043308,26.631927,29.224451,31.81307,32.129326,32.441677,32.757935,33.074192,33.386543,34.530533,35.67062,36.81461,37.9586,39.098682,39.688248,40.28172,40.871284,41.460846,42.05041,37.396366,32.746223,28.092175,23.438128,18.787983,17.671324,16.55857,15.441911,14.329156,13.212498,12.888432,12.564366,12.236397,11.912332,11.588266,9.331521,7.0786815,4.8219366,2.5690966,0.31235218,3.1586614,6.001066,8.847376,11.693685,14.53609,11.818625,9.097258,6.375889,3.6584249,0.93705654,1.6242313,2.3114061,2.998581,3.6857557,4.376835,5.2318993,6.083059,6.9381227,7.793187,8.648251,9.917182,11.186112,12.4511385,13.72007,14.989,13.751305,12.517513,11.283723,10.046027,8.812236,9.456462,10.096785,10.741011,11.381332,12.025558,14.161267,16.300879,18.436588,20.5762,22.711908,24.976461,27.241014,29.509472,31.774025,34.038578,29.966288,25.893995,21.821705,17.745508,13.673217,12.130978,10.584834,9.0386915,7.4964523,5.950309,5.6965227,5.4388323,5.185046,4.93126,4.6735697,5.2006636,5.7316628,6.2587566,6.785851,7.3129454,7.2739015,7.230953,7.191909,7.152865,7.113821,7.6916723,8.265619,8.843472,9.421323,9.999174,9.4291315,8.859089,8.289046,7.719003,7.1489606,7.676055,8.203149,8.734148,9.261242,9.788337,9.694631,9.600925,9.511124,9.4174185,9.323712,10.951848,12.579984,14.208119,15.836256,17.464392,16.578093,15.695697,14.813302,13.930907,13.048512,12.560462,12.068507,11.580457,11.088503,10.600452,15.562947,20.525442,25.487938,30.450434,35.41293,33.058575,30.70422,28.34596,25.991606,23.63725,21.470308,19.303364,17.136421,14.965574,12.798631,12.86891,12.935285,13.001659,13.0719385,13.138313,14.258877,15.375536,16.4961,17.616663,18.737226,15.808925,12.8767185,9.948417,7.016211,4.087909,3.7404175,3.3929255,3.0454338,2.697942,2.35045,2.533957,2.7213683,2.9048753,3.0883822,3.2757936,6.055728,8.835662,11.615597,14.395531,17.175465,14.668839,12.158309,9.651682,7.1450562,4.6384296,7.168483,9.702439,12.236397,14.766449,17.300406,18.214037,19.13157,20.0452,20.958832,21.876366,20.259943,18.64352,17.031002,15.41458,13.798158,11.115833,8.429605,5.743376,3.0610514,0.37482262,2.7330816,5.0913405,7.445695,9.803954,12.162213,10.373997,8.581876,6.79366,5.001539,3.213323,6.617962,10.0226,13.427239,16.831879,20.236517,18.003199,15.773785,13.540467,11.307149,9.073831,8.359325,7.6448197,6.930314,6.2158084,5.5013027,5.758993,6.0205884,6.278279,6.5398736,6.801469,6.4891167,6.180669,5.8683167,5.559869,5.251421,4.93126,4.6150036,4.298747,3.978586,3.6623292,3.619381,3.5725281,3.5256753,3.4827268,3.435874,2.8463092,2.25284,1.6593709,1.0659018,0.47633708,0.6637484,0.8511597,1.038571,1.2259823,1.4133936,1.1908426,0.96829176,0.74574083,0.5231899,0.30063897,0.24597734,0.19131571,0.13665408,0.078088045,0.023426414,0.15227169,0.28111696,0.40605783,0.5349031,0.6637484,0.79259366,0.92143893,1.0541886,1.183034,1.3118792,1.717937,2.1239948,2.5261483,2.9322062,3.338264,3.533484,3.7326086,3.9317331,4.126953,4.3260775,3.5295796,2.7330816,1.9404879,1.1439898,0.3513962,0.28111696,0.21083772,0.14055848,0.07027924,0.0,0.37872702,0.76135844,1.1400855,1.5188124,1.901444,1.5227169,1.1439898,0.76916724,0.39044023,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.1756981,0.31235218,0.44900626,0.58566034,0.7262188,0.76526284,0.80430686,0.8433509,0.8862993,0.92534333,0.76916724,0.60908675,0.45291066,0.29673457,0.13665408,0.16008049,0.1835069,0.20693332,0.22645533,0.24988174,0.25769055,0.26549935,0.27330816,0.28111696,0.28892577,0.26159495,0.23816854,0.21083772,0.18741131,0.1639849,0.14836729,0.13665408,0.12494087,0.113227665,0.10151446,0.093705654,0.08980125,0.08589685,0.078088045,0.07418364,0.16008049,0.24597734,0.3318742,0.41386664,0.4997635,0.48805028,0.48024148,0.46852827,0.46071947,0.44900626,0.62079996,0.79649806,0.96829176,1.1400855,1.3118792,1.1713207,1.0268579,0.8862993,0.7418364,0.60127795,0.5388075,0.47633708,0.41386664,0.3513962,0.28892577,0.28892577,0.29283017,0.29673457,0.29673457,0.30063897,0.28111696,0.26159495,0.23816854,0.21864653,0.19912452,0.19131571,0.1835069,0.1756981,0.1717937,0.1639849,0.14836729,0.13274968,0.11713207,0.10151446,0.08589685,1.0619974,2.0341935,3.0063896,3.978586,4.950782,4.9663997,4.9781127,4.9937305,5.009348,5.024966,4.493967,3.959064,3.4280653,2.893162,2.3621633,3.049338,3.7326086,4.415879,5.1030536,5.786324,10.373997,14.96167,19.549341,24.137014,28.724688,28.947239,29.169788,29.39234,29.614891,29.837442,31.469482,33.09762,34.725754,36.357796,37.98593,36.916122,35.846317,34.776512,33.706703,32.636898,47.231556,61.82621,76.41696,91.00771,105.598465,102.54522,99.488075,96.43483,93.38159,90.32444,101.4598,112.59125,123.7227,134.85416,145.9895,146.84848,147.71135,148.57422,149.43709,150.29996,135.14697,119.993996,104.84101,89.691925,74.53504,64.020485,53.502026,42.983566,32.46901,21.95055,19.260416,16.574188,13.887959,11.20173,8.511597,7.6955767,6.8756523,6.0596323,5.2436123,4.423688,4.193328,3.9668727,3.736513,3.506153,3.2757936,0.62470436,0.62079996,0.62079996,0.61689556,0.61689556,0.61299115,0.6481308,0.6832704,0.71841,0.75354964,0.78868926,0.81211567,0.8394465,0.8628729,0.8862993,0.9136301,0.96438736,1.0112402,1.0619974,1.1127546,1.1635119,1.261122,1.3626363,1.4641509,1.5617609,1.6632754,1.7686942,1.8780174,1.9834363,2.0927596,2.1981785,2.4792955,2.7565079,3.0337205,3.310933,3.5881457,3.6037633,3.619381,3.631094,3.6467118,3.6623292,3.6662338,3.6662338,3.6701381,3.6740425,3.6740425,3.8419318,4.009821,4.1777105,4.3455997,4.513489,5.2006636,5.8878384,6.575013,7.262188,7.9493628,7.726812,7.504261,7.28171,7.0591593,6.8366084,6.5008297,6.168956,5.833177,5.4973984,5.1616197,5.708236,6.250948,6.7975645,7.3441806,7.8868923,7.348085,6.813182,6.2743745,5.735567,5.2006636,5.7316628,6.2587566,6.7897553,7.320754,7.8517528,7.2036223,6.559396,5.9151692,5.270943,4.6267166,4.267512,3.9083066,3.5530062,3.193801,2.8385005,2.9907722,3.1469483,3.3031244,3.4593005,3.611572,4.7907014,5.9737353,7.152865,8.331994,9.511124,9.999174,10.48332,10.967466,11.4516115,11.935758,10.6355915,9.339331,8.039165,6.7389984,5.4388323,6.5398736,7.6409154,8.745861,9.846903,10.951848,10.741011,10.534078,10.327144,10.120211,9.913278,9.171441,8.4257,7.6838636,6.942027,6.2001905,7.3168497,8.433509,9.554072,10.670732,11.787391,10.588739,9.393991,8.19534,6.996689,5.801942,6.27047,6.7389984,7.211431,7.6799593,8.148487,8.398369,8.644346,8.894228,9.140205,9.386183,8.605303,7.824422,7.039637,6.2587566,5.473972,4.989826,4.50568,4.0215344,3.533484,3.049338,4.009821,4.970304,5.930787,6.89127,7.8517528,7.6721506,7.4964523,7.3168497,7.141152,6.9615493,5.8175592,4.6735697,3.5256753,2.3816853,1.2376955,2.463678,3.6935644,4.919547,6.1494336,7.375416,7.7307167,8.086017,8.441318,8.796618,9.151918,8.495979,7.8400397,7.1841,6.5281606,5.8761253,5.958118,6.044015,6.1299114,6.2158084,6.3017054,7.719003,9.140205,10.561408,11.978706,13.399908,14.590752,15.781594,16.968533,18.159374,19.350218,22.294136,25.234152,28.178072,31.12199,34.062004,34.967827,35.87365,36.77947,37.681385,38.587208,38.809757,39.03231,39.25486,39.47741,39.699963,39.65311,39.61016,39.56331,39.52036,39.473507,35.170856,30.8643,26.56165,22.255093,17.948538,16.968533,15.988527,15.008522,14.028518,13.048512,12.712734,12.376955,12.037272,11.701493,11.361811,9.140205,6.918601,4.6930914,2.4714866,0.24988174,3.2289407,6.2040954,9.183154,12.158309,15.137367,12.373051,9.608734,6.8405128,4.0761957,1.3118792,2.0380979,2.7643168,3.4866312,4.21285,4.939069,5.473972,6.008875,6.5437784,7.0786815,7.6135845,8.546737,9.483793,10.416945,11.354002,12.287154,11.869383,11.447707,11.0260315,10.608261,10.186585,10.920613,11.6585455,12.392572,13.1266,13.860628,16.398489,18.936352,21.474213,24.012074,26.549934,27.740778,28.935526,30.126368,31.321115,32.51196,29.579752,26.647545,23.71534,20.783133,17.850927,15.598087,13.345247,11.092407,8.839567,6.5867267,6.3017054,6.016684,5.7316628,5.446641,5.1616197,5.368553,5.571582,5.7785153,5.9815445,6.1884775,6.1572423,6.126007,6.098676,6.067441,6.036206,6.3915067,6.746807,7.1021075,7.4574084,7.812709,7.621393,7.433982,7.2426662,7.0513506,6.8639393,7.016211,7.172387,7.328563,7.480835,7.6370106,8.913751,10.194394,11.471134,12.747873,14.024612,14.805493,15.586374,16.36335,17.14423,17.92511,16.296974,14.668839,13.040704,11.416472,9.788337,10.569217,11.354002,12.134882,12.915763,13.700547,17.073952,20.45126,23.824663,27.201971,30.575375,29.103415,27.631454,26.15559,24.683632,23.211672,21.15405,19.092527,17.031002,14.973383,12.911859,12.997755,13.083652,13.165645,13.251541,13.337439,14.50095,15.668366,16.831879,17.999294,19.162806,16.8514,14.543899,12.232492,9.921086,7.6135845,6.79366,5.9737353,5.153811,4.3338866,3.513962,3.3460727,3.1781836,3.0102942,2.8424048,2.6745155,5.423215,8.16801,10.916709,13.665408,16.414106,14.684457,12.958711,11.229061,9.503315,7.773665,9.265146,10.756628,12.244205,13.735687,15.223265,16.75379,18.284315,19.814842,21.345367,22.875893,21.021301,19.16671,17.308216,15.453624,13.599033,11.00651,8.410083,5.813655,3.2211318,0.62470436,2.67842,4.728231,6.7819467,8.835662,10.889378,9.194867,7.504261,5.8097506,4.1191444,2.4246337,5.3334136,8.246098,11.154878,14.063657,16.976341,15.336493,13.696643,12.056794,10.413041,8.773191,7.918128,7.066968,6.211904,5.35684,4.5017757,4.845363,5.1889505,5.5364423,5.8800297,6.223617,6.278279,6.336845,6.3915067,6.446168,6.5008297,6.266566,6.028397,5.794133,5.559869,5.3256044,4.9234514,4.521298,4.1191444,3.7130866,3.310933,2.7916477,2.2684577,1.7452679,1.2220778,0.698888,0.77307165,0.8511597,0.92534333,0.999527,1.0737107,0.9058213,0.7340276,0.5661383,0.39434463,0.22645533,0.19131571,0.15617609,0.12103647,0.08589685,0.05075723,0.30454338,0.5583295,0.8160201,1.0698062,1.3235924,1.5851873,1.8467822,2.1044729,2.366068,2.6237583,3.408543,4.193328,4.9781127,5.7668023,6.551587,6.832704,7.113821,7.3988423,7.6799593,7.9610763,6.461786,4.958591,3.455396,1.9522011,0.44900626,0.359205,0.26940376,0.1796025,0.08980125,0.0,0.359205,0.71841,1.0815194,1.4407244,1.7999294,1.4446288,1.0893283,0.7340276,0.37872702,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.21083772,0.3513962,0.48805028,0.62470436,0.76135844,0.76916724,0.77307165,0.77697605,0.78088045,0.78868926,0.659844,0.5309987,0.40605783,0.27721256,0.14836729,0.1717937,0.19131571,0.21083772,0.23035973,0.24988174,0.25378615,0.25378615,0.25769055,0.26159495,0.26159495,0.23816854,0.21083772,0.18741131,0.1639849,0.13665408,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.078088045,0.078088045,0.08199245,0.08589685,0.08589685,0.20693332,0.3279698,0.44900626,0.5661383,0.6871748,0.7066968,0.7223144,0.7418364,0.75745404,0.77307165,0.9058213,1.038571,1.1713207,1.3040704,1.43682,1.2533131,1.0659018,0.8823949,0.698888,0.5114767,0.46071947,0.41386664,0.3631094,0.31235218,0.26159495,0.26940376,0.27330816,0.27721256,0.28111696,0.28892577,0.27330816,0.25769055,0.24207294,0.22645533,0.21083772,0.21083772,0.20693332,0.20693332,0.20302892,0.19912452,0.1835069,0.1639849,0.14836729,0.12884527,0.113227665,1.0307622,1.9522011,2.87364,3.7911747,4.7126136,4.60329,4.4978714,4.388548,4.283129,4.173806,3.7989833,3.4202564,3.0415294,2.6667068,2.2879796,3.06886,3.853645,4.6345253,5.4193106,6.2001905,10.71368,15.223265,19.736753,24.250242,28.763731,28.646599,28.525562,28.40843,28.291298,28.174168,29.447002,30.719837,31.992672,33.265507,34.53834,34.210373,33.882404,33.554432,33.226463,32.898495,43.986996,55.071594,66.15619,77.24079,88.325386,86.24044,84.15549,82.07053,79.98559,77.900635,86.728485,95.55634,104.38419,113.208145,122.035995,131.2621,140.4882,149.71431,158.93651,168.1626,156.68367,145.20082,133.72188,122.24293,110.763985,94.62709,78.4902,62.35721,46.224216,30.087324,26.05017,22.01302,17.975868,13.938716,9.901564,8.890324,7.8790836,6.871748,5.860508,4.8492675,4.728231,4.60329,4.482254,4.3612175,4.2362766,0.62470436,0.61689556,0.60518235,0.59346914,0.58566034,0.57394713,0.60127795,0.62860876,0.6559396,0.6832704,0.7106012,0.737932,0.76135844,0.78868926,0.81211567,0.8394465,0.9019169,0.96438736,1.0268579,1.0893283,1.1517987,1.2376955,1.3235924,1.4133936,1.4992905,1.5890918,1.7062237,1.8233559,1.9404879,2.05762,2.174752,2.4714866,2.7682211,3.06886,3.3655949,3.6623292,3.6232853,3.5842414,3.541293,3.5022488,3.4632049,3.4710135,3.4827268,3.49444,3.5022488,3.513962,3.8067923,4.1035266,4.396357,4.6930914,4.985922,5.4856853,5.989353,6.4891167,6.98888,7.4886436,7.2465706,7.008402,6.7663293,6.5281606,6.2860875,5.958118,5.6340523,5.3060827,4.9781127,4.650143,5.2318993,5.8097506,6.3915067,6.969358,7.551114,7.1997175,6.8483214,6.5008297,6.1494336,5.801942,6.5086384,7.2153354,7.9220324,8.628729,9.339331,8.445222,7.551114,6.66091,5.7668023,4.8765984,4.396357,3.9161155,3.435874,2.9556324,2.475391,2.5808098,2.690133,2.795552,2.9048753,3.0141985,4.2089458,5.4036927,6.5984397,7.793187,8.987934,9.538455,10.09288,10.6434,11.197825,11.748346,10.311526,8.874706,7.437886,6.001066,4.564246,5.2592297,5.958118,6.6531014,7.3519893,8.050878,8.257811,8.464745,8.671678,8.878611,9.085544,8.566258,8.046973,7.5276875,7.008402,6.4891167,7.28171,8.078208,8.870802,9.6673,10.4637985,9.761005,9.058213,8.355421,7.6526284,6.949836,7.4300776,7.910319,8.39056,8.870802,9.351044,9.265146,9.17925,9.093353,9.01136,8.925464,8.484266,8.039165,7.5979667,7.1567693,6.7116675,5.9464045,5.181142,4.415879,3.6506162,2.8892577,4.3260775,5.7668023,7.2075267,8.648251,10.088976,9.21439,8.343708,7.4691215,6.5984397,5.7238536,4.93126,4.138666,3.3460727,2.5534792,1.7608855,2.87364,3.9824903,5.0913405,6.2040954,7.3129454,7.793187,8.277332,8.761478,9.24172,9.725866,9.378374,9.034787,8.691199,8.343708,8.00012,8.191436,8.378847,8.570163,8.761478,8.94889,10.053836,11.158782,12.263727,13.368673,14.473619,15.54733,16.62104,17.690847,18.764557,19.838268,23.133583,26.4289,29.724215,33.01953,36.31094,37.806328,39.301712,40.7971,42.292484,43.787872,43.08898,42.394,41.69511,40.996223,40.30124,39.621876,38.938602,38.25924,37.579872,36.900505,32.94144,28.986282,25.027218,21.068155,17.112995,16.26574,15.422389,14.579038,13.731783,12.888432,12.537036,12.185639,11.838148,11.486752,11.139259,8.94889,6.75852,4.5681505,2.377781,0.18741131,3.2992198,6.407124,9.518932,12.626837,15.738646,12.927476,10.116306,7.309041,4.4978714,1.6867018,2.4480603,3.213323,3.9746814,4.73604,5.5013027,5.716045,5.930787,6.1455293,6.3602715,6.575013,7.1762915,7.7814736,8.382751,8.98403,9.589212,9.983557,10.377901,10.772245,11.166591,11.560935,12.388668,13.216402,14.044135,14.871868,15.699601,18.635712,21.575727,24.511837,27.451853,30.387962,30.508999,30.626131,30.747168,30.868204,30.98924,29.193216,27.401094,25.608974,23.816854,22.024733,19.065197,16.10566,13.146122,10.186585,7.223144,6.910792,6.5945354,6.278279,5.9659266,5.64967,5.532538,5.4154058,5.298274,5.181142,5.0640097,5.040583,5.0210614,5.001539,4.9820175,4.9624953,5.095245,5.2279944,5.3607445,5.493494,5.6262436,5.813655,6.0049706,6.196286,6.3836975,6.575013,6.356367,6.141625,5.9229784,5.704332,5.4856853,8.136774,10.783959,13.431144,16.07833,18.725513,18.659138,18.58886,18.522484,18.45611,18.38583,16.015858,13.641981,11.268105,8.898132,6.524256,8.581876,10.6355915,12.689307,14.746927,16.800642,18.58886,20.37317,22.161386,23.949604,25.73782,25.148254,24.558691,23.969126,23.375656,22.78609,20.83389,18.88169,16.92949,14.977287,13.025085,13.1266,13.228115,13.333533,13.435048,13.536563,14.746927,15.957292,17.167656,18.378021,19.588387,17.89778,16.207174,14.516567,12.825961,11.139259,9.846903,8.554545,7.2582836,5.9659266,4.6735697,4.154284,3.6349986,3.1157131,2.5964274,2.0732377,4.7907014,7.504261,10.221725,12.935285,15.648844,14.703979,13.755209,12.806439,11.861574,10.912805,11.361811,11.806912,12.2559185,12.70102,13.150026,15.293544,17.440966,19.584482,21.731903,23.87542,21.778755,19.685997,17.589333,15.4965725,13.399908,10.893282,8.39056,5.883934,3.3812122,0.8745861,2.6237583,4.369026,6.1181984,7.8634663,9.612638,8.015738,6.422742,4.825841,3.232845,1.6359446,4.0527697,6.46569,8.882515,11.29934,13.712261,12.665881,11.615597,10.569217,9.522837,8.476458,7.480835,6.4852123,5.4895897,4.493967,3.4983444,3.9317331,4.3612175,4.7907014,5.2201858,5.64967,6.0713453,6.4891167,6.910792,7.328563,7.7502384,7.5979667,7.445695,7.2934237,7.141152,6.98888,6.2275214,5.466163,4.7087092,3.9473507,3.1859922,2.7330816,2.2840753,1.8311646,1.3782539,0.92534333,0.8862993,0.8511597,0.81211567,0.77307165,0.737932,0.62079996,0.5036679,0.38653582,0.26940376,0.14836729,0.13665408,0.12103647,0.10541886,0.08980125,0.07418364,0.45681506,0.8394465,1.2220778,1.6047094,1.9873407,2.377781,2.7682211,3.1586614,3.5491016,3.9356375,5.1030536,6.266566,7.433982,8.597494,9.761005,10.131924,10.498938,10.865952,11.232965,11.599979,9.390087,7.180196,4.970304,2.7604125,0.5505207,0.44119745,0.3318742,0.21864653,0.10932326,0.0,0.339683,0.679366,1.0190489,1.358732,1.698415,1.3665408,1.0346665,0.7027924,0.3709182,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.24988174,0.38653582,0.5231899,0.6637484,0.80040246,0.76916724,0.7418364,0.7106012,0.679366,0.6481308,0.5544251,0.45681506,0.359205,0.26159495,0.1639849,0.1796025,0.19912452,0.21474212,0.23426414,0.24988174,0.24597734,0.24597734,0.24207294,0.23816854,0.23816854,0.21083772,0.18741131,0.1639849,0.13665408,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.058566034,0.07027924,0.078088045,0.08980125,0.10151446,0.25378615,0.40996224,0.5661383,0.71841,0.8745861,0.92143893,0.96438736,1.0112402,1.0541886,1.1010414,1.1908426,1.2845483,1.3782539,1.4680552,1.5617609,1.3353056,1.1088502,0.8784905,0.6520352,0.42557985,0.38653582,0.3513962,0.31235218,0.27330816,0.23816854,0.24597734,0.25378615,0.26159495,0.26940376,0.27330816,0.26549935,0.25378615,0.24597734,0.23426414,0.22645533,0.22645533,0.23035973,0.23426414,0.23426414,0.23816854,0.21864653,0.19912452,0.1756981,0.15617609,0.13665408,1.0034313,1.8741131,2.7408905,3.6076677,4.474445,4.2440853,4.0137253,3.7833657,3.5569105,3.3265507,3.1039999,2.8814487,2.6588979,2.436347,2.2137961,3.0922866,3.970777,4.853172,5.7316628,6.6140575,11.0494585,15.488764,19.924164,24.36347,28.79887,28.342056,27.88524,27.428427,26.971611,26.510891,27.428427,28.342056,29.255686,30.173222,31.086851,31.500717,31.918488,32.332355,32.746223,33.163994,40.738533,48.31698,55.895424,63.469963,71.04841,69.93565,68.81899,67.70624,66.58958,65.47292,71.99718,78.52143,85.04179,91.56213,98.086395,115.67573,133.26506,150.85048,168.43591,186.02524,178.21645,170.41154,162.60274,154.79784,146.98903,125.2337,103.48228,81.73085,59.979427,38.2241,32.83602,27.447948,22.063778,16.675701,11.287627,10.085071,8.882515,7.6799593,6.477403,5.2748475,5.2592297,5.2436123,5.2318993,5.2162814,5.2006636,0.62470436,0.60908675,0.58956474,0.57394713,0.5544251,0.5388075,0.5583295,0.57785153,0.59737355,0.61689556,0.63641757,0.6637484,0.6871748,0.7106012,0.737932,0.76135844,0.8394465,0.9136301,0.9878138,1.0619974,1.1361811,1.2142692,1.2884527,1.3626363,1.43682,1.5110037,1.639849,1.7686942,1.893635,2.0224805,2.1513257,2.4675822,2.7838387,3.1039999,3.4202564,3.736513,3.6428072,3.5491016,3.4514916,3.357786,3.2640803,3.279698,3.2992198,3.3148375,3.3343596,3.349977,3.7716527,4.193328,4.618908,5.040583,5.462259,5.774611,6.086963,6.3993154,6.7116675,7.0240197,6.7663293,6.5086384,6.250948,5.9932575,5.735567,5.4193106,5.099149,4.7789884,4.4588275,4.138666,4.7516575,5.368553,5.9815445,6.5984397,7.211431,7.0513506,6.8873653,6.7233806,6.5633,6.3993154,7.2856145,8.171914,9.054309,9.940608,10.826907,9.686822,8.546737,7.406651,6.266566,5.12648,4.521298,3.9200199,3.3187418,2.7135596,2.1122816,2.1708477,2.233318,2.2918842,2.3543546,2.4129205,3.6232853,4.83365,6.044015,7.2543793,8.460839,9.081639,9.702439,10.323239,10.944039,11.560935,9.987461,8.413987,6.8366084,5.263134,3.6857557,3.978586,4.271416,4.564246,4.8570766,5.1499066,5.7707067,6.395411,7.016211,7.6409154,8.261715,7.9649806,7.6682463,7.3715115,7.0708723,6.774138,7.2465706,7.719003,8.191436,8.663869,9.136301,8.929368,8.722435,8.515501,8.308568,8.101635,8.589685,9.081639,9.56969,10.061645,10.549695,10.131924,9.714153,9.296382,8.878611,8.460839,8.359325,8.257811,8.156297,8.050878,7.9493628,6.9068875,5.860508,4.814128,3.7716527,2.7252727,4.646239,6.5633,8.484266,10.405232,12.326198,10.756628,9.190963,7.621393,6.055728,4.4861584,4.0488653,3.6076677,3.1664703,2.7291772,2.2879796,3.279698,4.271416,5.263134,6.2587566,7.250475,7.859562,8.468649,9.081639,9.690726,10.299813,10.264673,10.229534,10.194394,10.159255,10.124115,10.42085,10.71368,11.010414,11.303245,11.599979,12.388668,13.181262,13.969952,14.75864,15.551234,16.503908,17.460487,18.41316,19.36974,20.326319,23.97303,27.619741,31.266453,34.913166,38.56378,40.64873,42.733685,44.818634,46.903584,48.988537,47.36821,45.751785,44.135365,42.51894,40.898613,39.586735,38.27095,36.955166,35.639385,34.3236,30.715933,27.10436,23.496693,19.88512,16.273548,15.566852,14.856251,14.145649,13.435048,12.724447,12.361338,11.998228,11.639023,11.275913,10.912805,8.75367,6.5984397,4.4393053,2.2840753,0.12494087,3.3655949,6.610153,9.850807,13.095366,16.33602,13.481901,10.627783,7.773665,4.9156423,2.0615244,2.8619268,3.6623292,4.462732,5.263134,6.0635366,5.958118,5.852699,5.74728,5.6418614,5.5364423,5.805846,6.0791545,6.348558,6.617962,6.8873653,8.097731,9.308095,10.518459,11.728825,12.939189,13.856724,14.778163,15.695697,16.617136,17.538574,20.876839,24.211199,27.549461,30.887726,34.22599,33.273315,32.32064,31.367968,30.415293,29.46262,28.810585,28.158548,27.506514,26.854479,26.19854,22.532305,18.866072,15.195933,11.5297,7.8634663,7.5159745,7.172387,6.8287997,6.481308,6.13772,5.6965227,5.2592297,4.8180323,4.376835,3.9356375,3.9278288,3.9161155,3.9083066,3.8965936,3.8887846,3.7989833,3.7091823,3.619381,3.5256753,3.435874,4.0059166,4.575959,5.1460023,5.716045,6.2860875,5.6965227,5.1069584,4.5173936,3.9278288,3.338264,7.355894,11.373524,15.391153,19.408783,23.426414,22.508879,21.59525,20.68162,19.764084,18.850454,15.730837,12.615124,9.495506,6.379793,3.2640803,6.590631,9.917182,13.243732,16.574188,19.900738,20.099863,20.298986,20.498112,20.701141,20.900265,21.193096,21.485926,21.778755,22.071587,22.364416,20.517633,18.67085,16.827974,14.981192,13.138313,13.25935,13.376482,13.497519,13.618555,13.735687,14.992905,16.246218,17.503435,18.756748,20.013966,18.94416,17.874353,16.800642,15.730837,14.661031,12.89624,11.131451,9.366661,7.601871,5.8370814,4.9663997,4.0918136,3.2211318,2.3465457,1.475864,4.1581883,6.8405128,9.522837,12.205161,14.8874855,14.719597,14.551707,14.383818,14.215929,14.051944,13.45457,12.861101,12.263727,11.6702585,11.076789,13.833297,16.59371,19.354122,22.114534,24.874947,22.540113,20.205282,17.87045,15.535617,13.200784,10.783959,8.371038,5.9542136,3.541293,1.1244678,2.5690966,4.009821,5.45445,6.8951745,8.335898,6.8405128,5.3412223,3.8458362,2.3465457,0.8511597,2.7682211,4.689187,6.610153,8.531119,10.44818,9.99527,9.538455,9.085544,8.628729,8.175818,7.039637,5.903456,4.7711797,3.6349986,2.4988174,3.0141985,3.5295796,4.044961,4.560342,5.0757227,5.860508,6.6452928,7.4300776,8.214863,8.999647,8.929368,8.859089,8.78881,8.718531,8.648251,7.531592,6.4149327,5.298274,4.181615,3.0610514,2.67842,2.2957885,1.9131571,1.53443,1.1517987,0.999527,0.8511597,0.698888,0.5505207,0.39824903,0.3357786,0.26940376,0.20693332,0.14055848,0.07418364,0.078088045,0.08589685,0.08980125,0.093705654,0.10151446,0.60908675,1.1205635,1.6281357,2.1396124,2.6510892,3.1703746,3.68966,4.2089458,4.728231,5.251421,6.79366,8.339804,9.885946,11.428185,12.974329,13.427239,13.88015,14.33306,14.785972,15.238882,12.318389,9.4018,6.4852123,3.5686235,0.6481308,0.5192855,0.39044023,0.26159495,0.12884527,0.0,0.32016098,0.64032197,0.96048295,1.2806439,1.6008049,1.2884527,0.98000497,0.6715572,0.359205,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.28892577,0.42557985,0.5622339,0.698888,0.8394465,0.77307165,0.7066968,0.6442264,0.57785153,0.5114767,0.44510186,0.37872702,0.30844778,0.24207294,0.1756981,0.19131571,0.20693332,0.21864653,0.23426414,0.24988174,0.24207294,0.23426414,0.22645533,0.21864653,0.21083772,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.042948425,0.058566034,0.078088045,0.093705654,0.113227665,0.30063897,0.49195468,0.6832704,0.8706817,1.0619974,1.1361811,1.2064602,1.2806439,1.3509232,1.4251068,1.475864,1.5305257,1.5812829,1.6359446,1.6867018,1.4172981,1.1478943,0.8784905,0.60908675,0.3357786,0.31235218,0.28892577,0.26159495,0.23816854,0.21083772,0.22255093,0.23426414,0.24207294,0.25378615,0.26159495,0.25769055,0.25378615,0.24597734,0.24207294,0.23816854,0.24597734,0.25378615,0.26159495,0.26940376,0.27330816,0.25378615,0.23035973,0.20693332,0.1835069,0.1639849,0.97610056,1.7921207,2.6081407,3.4241607,4.2362766,3.8848803,3.533484,3.1781836,2.8267872,2.475391,2.4090161,2.338737,2.2723622,2.2059872,2.135708,3.1157131,4.0918136,5.0718184,6.0479193,7.0240197,11.389141,15.750359,20.111576,24.472794,28.837915,28.041416,27.241014,26.444517,25.648018,24.85152,25.405945,25.964275,26.522604,27.080935,27.639263,28.794966,29.95067,31.110277,32.26598,33.425587,37.493977,41.566265,45.634655,49.70304,53.775333,53.63087,53.48641,53.33804,53.193577,53.049114,57.26587,61.486526,65.70328,69.92004,74.13679,100.089355,126.041916,151.98666,177.93532,203.88788,199.75313,195.61836,191.4836,187.34883,183.21408,155.84032,128.47046,101.10059,73.734634,46.360874,39.62578,32.88678,26.151686,19.412687,12.67369,11.279819,9.885946,8.488171,7.094299,5.700427,5.794133,5.883934,5.9776397,6.0713453,6.1611466,0.62470436,0.60127795,0.57394713,0.5505207,0.5231899,0.4997635,0.5114767,0.5231899,0.5388075,0.5505207,0.5622339,0.58566034,0.61299115,0.63641757,0.6637484,0.6871748,0.77307165,0.8628729,0.94876975,1.038571,1.1244678,1.1869383,1.2494087,1.3118792,1.3743496,1.43682,1.5734742,1.7140326,1.8506867,1.9873407,2.1239948,2.463678,2.7994564,3.1391394,3.474918,3.8106966,3.6623292,3.513962,3.3616903,3.213323,3.0610514,3.0883822,3.1118085,3.1391394,3.1625657,3.1859922,3.736513,4.2870336,4.8375545,5.388075,5.938596,6.0635366,6.1884775,6.3134184,6.4383593,6.5633,6.2860875,6.012779,5.735567,5.462259,5.1889505,4.8765984,4.564246,4.251894,3.9356375,3.6232853,4.2753205,4.9234514,5.575486,6.223617,6.8756523,6.899079,6.9264097,6.949836,6.9732623,7.000593,8.062591,9.124588,10.186585,11.248583,12.31058,10.924518,9.538455,8.148487,6.7624245,5.376362,4.650143,3.9239242,3.2016098,2.475391,1.7491722,1.7608855,1.7765031,1.7882162,1.7999294,1.8116426,3.0376248,4.263607,5.4856853,6.7116675,7.9376497,8.624825,9.311999,9.999174,10.686349,11.373524,9.663396,7.9493628,6.239235,4.5252023,2.8111696,2.7018464,2.5886188,2.475391,2.3621633,2.2489357,3.2875066,4.3260775,5.3607445,6.3993154,7.437886,7.363703,7.2856145,7.211431,7.137247,7.0630636,7.211431,7.363703,7.5120697,7.6643414,7.812709,8.101635,8.386656,8.675582,8.960603,9.249529,9.749292,10.249056,10.748819,11.248583,11.748346,10.998701,10.249056,9.499411,8.749765,8.00012,8.238289,8.476458,8.710721,8.94889,9.187058,7.8634663,6.5359693,5.212377,3.8887846,2.5612879,4.9624953,7.363703,9.761005,12.162213,14.56342,12.298867,10.0382185,7.773665,5.5130157,3.2484627,3.1625657,3.076669,2.9868677,2.900971,2.8111696,3.6857557,4.564246,5.4388323,6.3134184,7.1880045,7.9259367,8.663869,9.4018,10.135828,10.87376,11.150972,11.424281,11.701493,11.974802,12.24811,12.650263,13.048512,13.450665,13.848915,14.251068,14.723501,15.199838,15.676175,16.148607,16.624945,17.464392,18.299932,19.13938,19.974922,20.81437,24.812477,28.810585,32.812595,36.810703,40.812717,43.487232,46.161747,48.83626,51.51078,54.189198,51.651337,49.113476,46.575615,44.037754,41.499893,39.551594,37.599392,35.651096,33.698895,31.750599,28.486519,25.226343,21.962263,18.698183,15.438006,14.864059,14.286208,13.712261,13.138313,12.564366,12.185639,11.810817,11.435994,11.061172,10.686349,8.562354,6.4383593,4.3143644,2.1864653,0.062470436,3.435874,6.813182,10.186585,13.563893,16.937298,14.036326,11.139259,8.238289,5.337318,2.436347,3.2757936,4.1113358,4.950782,5.786324,6.6257706,6.2001905,5.774611,5.349031,4.9234514,4.5017757,4.4393053,4.376835,4.3143644,4.251894,4.1894236,6.211904,8.238289,10.260769,12.287154,14.313539,15.324779,16.33602,17.351164,18.362404,19.373644,23.114061,26.850574,30.587088,34.3236,38.06402,36.037632,34.01125,31.988768,29.962383,27.935999,28.42405,28.912098,29.400148,29.888199,30.37625,25.999414,21.626484,17.24965,12.8767185,8.499884,8.125061,7.7502384,7.375416,7.000593,6.6257706,5.8644123,5.099149,4.337791,3.5764325,2.8111696,2.8111696,2.8111696,2.8111696,2.8111696,2.8111696,2.4988174,2.1864653,1.8741131,1.5617609,1.2494087,2.1981785,3.1508527,4.0996222,5.0483923,6.001066,5.036679,4.0761957,3.1118085,2.1513257,1.1869383,6.575013,11.963089,17.351164,22.739239,28.12341,26.362524,24.601639,22.83685,21.075964,19.311174,15.449719,11.588266,7.726812,3.8614538,0.0,4.5993857,9.198771,13.802062,18.401447,23.000834,21.610867,20.224804,18.838741,17.448774,16.062712,17.237936,18.41316,19.588387,20.76361,21.938837,20.201378,18.463919,16.72646,14.989,13.251541,13.388195,13.524849,13.661504,13.798158,13.938716,15.238882,16.539047,17.839214,19.13938,20.435642,19.986635,19.537628,19.088623,18.635712,18.186707,15.949483,13.712261,11.475039,9.237816,7.000593,5.774611,4.548629,3.3265507,2.1005683,0.8745861,3.5256753,6.1767645,8.823949,11.475039,14.126127,14.739119,15.348206,15.961197,16.574188,17.18718,15.551234,13.911386,12.27544,10.6355915,8.999647,12.376955,15.750359,19.123762,22.50107,25.874474,23.301472,20.724567,18.151566,15.57466,13.001659,10.674636,8.351517,6.0244927,3.7013733,1.3743496,2.514435,3.6506162,4.786797,5.9268827,7.0630636,5.661383,4.263607,2.8619268,1.4641509,0.062470436,1.4875772,2.912684,4.337791,5.7628975,7.1880045,7.3246584,7.461313,7.601871,7.7385254,7.8751793,6.5984397,5.3256044,4.0488653,2.77603,1.4992905,2.1005683,2.7018464,3.2992198,3.900498,4.5017757,5.64967,6.801469,7.9493628,9.101162,10.249056,10.260769,10.276386,10.2881,10.299813,10.311526,8.835662,7.363703,5.8878384,4.4119744,2.9361105,2.6237583,2.3114061,1.999054,1.6867018,1.3743496,1.1127546,0.8511597,0.58566034,0.3240654,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.76135844,1.4016805,2.0380979,2.6745155,3.310933,3.9629683,4.6110992,5.263134,5.911265,6.5633,8.488171,10.413041,12.337912,14.262781,16.187653,16.72646,17.261362,17.800169,18.338978,18.87388,15.250595,11.623405,8.00012,4.376835,0.74964523,0.60127795,0.44900626,0.30063897,0.14836729,0.0,0.30063897,0.60127795,0.9019169,1.1986516,1.4992905,1.2142692,0.92534333,0.63641757,0.3513962,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.3240654,0.46071947,0.60127795,0.737932,0.8745861,0.77307165,0.6754616,0.57394713,0.47633708,0.37482262,0.3357786,0.30063897,0.26159495,0.22645533,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,0.23816854,0.22645533,0.21083772,0.19912452,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.3513962,0.57394713,0.80040246,1.0268579,1.2494087,1.3509232,1.4485333,1.5500476,1.6515622,1.7491722,1.7608855,1.7765031,1.7882162,1.7999294,1.8116426,1.4992905,1.1869383,0.8745861,0.5622339,0.24988174,0.23816854,0.22645533,0.21083772,0.19912452,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.26159495,0.27330816,0.28892577,0.30063897,0.31235218,0.28892577,0.26159495,0.23816854,0.21083772,0.18741131,0.94876975,1.7140326,2.475391,3.2367494,3.998108,3.5256753,3.049338,2.5769055,2.1005683,1.6242313,1.7140326,1.7999294,1.8858263,1.9756275,2.0615244,3.1391394,4.21285,5.2865605,6.364176,7.437886,11.72492,16.011953,20.298986,24.586021,28.873055,27.736874,26.600693,25.460608,24.324427,23.188246,23.38737,23.586494,23.785618,23.988647,24.187773,26.089216,27.986755,29.888199,31.785738,33.687183,34.249416,34.81165,35.373886,35.93612,36.498352,37.326084,38.149914,38.973743,39.801476,40.625305,42.538464,44.45162,46.360874,48.27403,50.187187,84.502975,118.814865,153.12675,187.43474,221.75052,221.2859,220.82518,220.36057,219.89984,219.43912,186.44691,153.45863,120.474236,87.489845,54.501553,46.41163,38.32561,30.235691,22.149673,14.063657,12.4745655,10.885473,9.300286,7.7111945,6.126007,6.3251314,6.524256,6.7233806,6.9264097,7.125534,0.58566034,0.58566034,0.58175594,0.58175594,0.57785153,0.57394713,0.58566034,0.60127795,0.61299115,0.62470436,0.63641757,0.6481308,0.6637484,0.6754616,0.6871748,0.698888,0.78088045,0.8589685,0.94096094,1.0190489,1.1010414,1.1713207,1.2455044,1.3157835,1.3899672,1.4641509,1.6008049,1.737459,1.8741131,2.0107672,2.1513257,2.436347,2.7213683,3.0063896,3.2914112,3.5764325,3.5451972,3.513962,3.4866312,3.455396,3.4241607,3.4514916,3.4788225,3.506153,3.533484,3.5608149,3.9942036,4.423688,4.853172,5.282656,5.7121406,5.7668023,5.8175592,5.8683167,5.9229784,5.9737353,5.7316628,5.4895897,5.2475166,5.0054436,4.7633705,4.5369153,4.3143644,4.087909,3.8614538,3.638903,4.40807,5.181142,5.9542136,6.727285,7.5003567,7.621393,7.7385254,7.859562,7.9805984,8.101635,8.921559,9.745388,10.569217,11.389141,12.212971,11.096312,9.983557,8.866898,7.7541428,6.6374836,5.6691923,4.7009,3.736513,2.7682211,1.7999294,1.7686942,1.7335546,1.7023194,1.6710842,1.6359446,2.8111696,3.9863946,5.1616197,6.336845,7.5120697,8.316377,9.120684,9.928895,10.733202,11.537509,9.768814,7.996216,6.2275214,4.4588275,2.6862288,2.6354716,2.5808098,2.5300527,2.4792955,2.4246337,3.4593005,4.493967,5.5286336,6.5633,7.601871,7.4300776,7.2582836,7.0903945,6.918601,6.7507114,6.8951745,7.039637,7.1841,7.328563,7.47693,7.687768,7.898606,8.113348,8.324185,8.538928,8.976221,9.413514,9.850807,10.2881,10.725393,10.272482,9.8195715,9.366661,8.913751,8.460839,8.550641,8.636538,8.726339,8.812236,8.898132,7.996216,7.0903945,6.184573,5.278752,4.376835,6.329036,8.285142,10.241247,12.193448,14.149553,11.935758,9.725866,7.5120697,5.298274,3.0883822,2.9634414,2.8385005,2.7135596,2.5886188,2.463678,3.1391394,3.8185053,4.493967,5.173333,5.8487945,6.5398736,7.230953,7.918128,8.609207,9.300286,9.643873,9.991365,10.334952,10.67854,11.0260315,11.771772,12.513609,13.25935,14.005091,14.750832,15.258404,15.76988,16.281357,16.788929,17.300406,18.432684,19.56496,20.697237,21.829514,22.96179,26.245392,29.528994,32.808693,36.092293,39.375896,42.921093,46.46629,50.01149,53.556686,57.101883,54.32195,51.545918,48.765984,45.989956,43.213924,40.890804,38.567684,36.244568,33.921448,31.598328,28.119505,24.636778,21.15405,17.671324,14.188598,13.743496,13.298394,12.853292,12.408191,11.963089,11.557031,11.150972,10.748819,10.342762,9.936704,8.109444,6.282183,4.454923,2.6276627,0.80040246,3.4280653,6.055728,8.683391,11.311053,13.938716,11.947471,9.956225,7.968885,5.9776397,3.9863946,4.6540475,5.3217,5.989353,6.657006,7.3246584,6.7311897,6.133816,5.5403466,4.9468775,4.349504,4.7087092,5.0640097,5.423215,5.7785153,6.13772,8.039165,9.936704,11.838148,13.735687,15.637131,16.113468,16.585901,17.062239,17.538574,18.011007,22.1731,26.339098,30.50119,34.663284,38.825375,36.677956,34.530533,32.383114,30.235691,28.08827,28.529467,28.970665,29.415766,29.856964,30.29816,26.179018,22.05597,17.93292,13.809871,9.686822,9.20658,8.726339,8.246098,7.7658563,7.2856145,6.590631,5.891743,5.196759,4.4978714,3.7989833,3.8419318,3.8809757,3.9200199,3.959064,3.998108,3.638903,3.279698,2.920493,2.5612879,2.1981785,2.9243972,3.6506162,4.376835,5.099149,5.825368,5.165524,4.50568,3.8458362,3.1859922,2.5261483,7.1060123,11.685876,16.26574,20.845604,25.425468,23.438128,21.45469,19.471254,17.483913,15.500477,13.048512,10.600452,8.148487,5.700427,3.2484627,6.7429028,10.2334385,13.727879,17.218414,20.712854,19.615717,18.51858,17.421442,16.324306,15.223265,16.152512,17.08176,18.007103,18.936352,19.861694,18.436588,17.01148,15.586374,14.161267,12.73616,12.771299,12.806439,12.841579,12.8767185,12.911859,14.294017,15.672271,17.054428,18.432684,19.810938,19.07691,18.342882,17.608854,16.870922,16.136894,14.512663,12.888432,11.2642,9.636065,8.011833,7.336372,6.66091,5.989353,5.3138914,4.6384296,6.153338,7.6721506,9.190963,10.705871,12.224684,12.857197,13.48971,14.122223,14.754736,15.387249,14.301826,13.212498,12.123169,11.037745,9.948417,13.06413,16.175938,19.287746,22.399555,25.511364,23.820759,22.134056,20.44345,18.752844,17.062239,15.180316,13.298394,11.416472,9.530646,7.648724,7.8400397,8.031356,8.218767,8.410083,8.601398,6.942027,5.2865605,3.6271896,1.9717231,0.31235218,1.4407244,2.5730011,3.7013733,4.83365,5.9620223,6.055728,6.153338,6.2470436,6.3407493,6.4383593,5.704332,4.9663997,4.2323723,3.4983444,2.7643168,2.9439192,3.1235218,3.3031244,3.4827268,3.6623292,4.7087092,5.7511845,6.7975645,7.843944,8.886419,8.769287,8.652155,8.535024,8.4178915,8.300759,7.1177254,5.9346914,4.7516575,3.5686235,2.3855898,2.1591344,1.9326792,1.7062237,1.475864,1.2494087,1.0112402,0.76916724,0.5309987,0.28892577,0.05075723,0.31625658,0.58175594,0.8433509,1.1088502,1.3743496,1.3314011,1.2845483,1.2415999,1.1947471,1.1517987,1.8506867,2.5495746,3.2484627,3.951255,4.650143,5.040583,5.434928,5.8292727,6.2197127,6.6140575,8.13287,9.651682,11.174399,12.693212,14.212025,15.141272,16.074425,17.003672,17.93292,18.862167,15.543426,12.228588,8.909846,5.591104,2.2762666,1.8858263,1.4953861,1.1049459,0.7145056,0.3240654,0.5036679,0.679366,0.8589685,1.0346665,1.2142692,1.0112402,0.81211567,0.61299115,0.41386664,0.21083772,0.1717937,0.12884527,0.08589685,0.042948425,0.0,0.031235218,0.06637484,0.09761006,0.12884527,0.1639849,0.28502136,0.40605783,0.5309987,0.6520352,0.77307165,0.6832704,0.59346914,0.5036679,0.41386664,0.3240654,0.29283017,0.26159495,0.22645533,0.19522011,0.1639849,0.1756981,0.19131571,0.20693332,0.22255093,0.23816854,0.23035973,0.22255093,0.21474212,0.20693332,0.19912452,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.14446288,0.15227169,0.16008049,0.1678893,0.1756981,0.1796025,0.1835069,0.19131571,0.19522011,0.19912452,0.40605783,0.60908675,0.8160201,1.0190489,1.2259823,1.3431144,1.4641509,1.5851873,1.7062237,1.8233559,1.7804074,1.7335546,1.6906061,1.6437533,1.6008049,1.3353056,1.0698062,0.80430686,0.5388075,0.27330816,0.26159495,0.24597734,0.23035973,0.21474212,0.19912452,0.20693332,0.21474212,0.22255093,0.23035973,0.23816854,0.23426414,0.22645533,0.22255093,0.21864653,0.21083772,0.23426414,0.25378615,0.27330816,0.29283017,0.31235218,0.30063897,0.29283017,0.28111696,0.27330816,0.26159495,0.9058213,1.5539521,2.1981785,2.8424048,3.4866312,3.06886,2.6471848,2.2294137,1.8077383,1.3860629,1.6164225,1.8467822,2.077142,2.3075018,2.5378613,3.4436827,4.3534083,5.2592297,6.168956,7.0747766,10.897186,14.719597,18.542006,22.364416,26.186827,25.417658,24.64849,23.879324,23.106253,22.337086,22.383938,22.430792,22.481548,22.5284,22.575254,25.484034,28.388908,31.297688,34.206467,37.111343,36.951263,36.791183,36.631104,36.47102,36.31094,36.271896,36.228947,36.186,36.14305,36.1001,37.583775,39.071354,40.555027,42.0387,43.526276,71.54817,99.57397,127.591965,155.61386,183.63965,184.22531,184.81488,185.40054,185.9862,186.57576,161.03317,135.49057,109.95578,84.41708,58.87448,50.12081,41.36714,32.61738,23.863707,15.113941,13.407718,11.701493,9.999174,8.292951,6.5867267,6.5672045,6.547683,6.5281606,6.5086384,6.4891167,0.5505207,0.5700427,0.58956474,0.60908675,0.62860876,0.6481308,0.6637484,0.6754616,0.6871748,0.698888,0.7106012,0.7106012,0.7106012,0.7106012,0.7106012,0.7106012,0.78478485,0.8589685,0.92924774,1.0034313,1.0737107,1.1557031,1.2415999,1.3235924,1.4055848,1.4875772,1.6242313,1.7608855,1.901444,2.0380979,2.174752,2.4090161,2.639376,2.87364,3.1039999,3.338264,3.4280653,3.5178664,3.6076677,3.697469,3.78727,3.8185053,3.8458362,3.8770714,3.9083066,3.9356375,4.2479897,4.5564375,4.8687897,5.1772375,5.4856853,5.466163,5.446641,5.4271193,5.407597,5.388075,5.1772375,4.9663997,4.755562,4.548629,4.337791,4.2011366,4.0605783,3.9239242,3.78727,3.6506162,4.5447245,5.4388323,6.336845,7.230953,8.125061,8.339804,8.554545,8.769287,8.98403,9.198771,9.784432,10.366188,10.947944,11.5297,12.111456,11.268105,10.4286585,9.585307,8.741957,7.898606,6.688241,5.481781,4.271416,3.0610514,1.8506867,1.7725986,1.6945106,1.6164225,1.5383345,1.4641509,2.5886188,3.7130866,4.8375545,5.9620223,7.08649,8.011833,8.933272,9.854712,10.77615,11.701493,9.874233,8.046973,6.2158084,4.388548,2.5612879,2.5690966,2.5769055,2.5847144,2.592523,2.6003318,3.631094,4.6657605,5.6965227,6.7311897,7.7619514,7.4964523,7.230953,6.969358,6.703859,6.4383593,6.578918,6.715572,6.8561306,6.996689,7.137247,7.2739015,7.4105554,7.551114,7.687768,7.824422,8.1992445,8.574067,8.94889,9.323712,9.698535,9.546264,9.390087,9.2339115,9.081639,8.925464,8.862993,8.800523,8.738052,8.675582,8.6131115,8.128965,7.6409154,7.1567693,6.6726236,6.1884775,7.6955767,9.20658,10.717585,12.228588,13.735687,11.576552,9.413514,7.250475,5.087436,2.9243972,2.7643168,2.6003318,2.436347,2.2762666,2.1122816,2.592523,3.0727646,3.5530062,4.0332475,4.513489,5.153811,5.7980375,6.4383593,7.082586,7.726812,8.140678,8.554545,8.968412,9.386183,9.80005,10.889378,11.978706,13.0719385,14.161267,15.250595,15.793307,16.339924,16.88654,17.429253,17.975868,19.400974,20.829987,22.258997,23.684105,25.113115,27.678308,30.2435,32.808693,35.373886,37.939075,42.35105,46.76693,51.182808,55.598686,60.010662,56.996464,53.978363,50.96026,47.942154,44.924053,42.230015,39.535976,36.838036,34.143997,31.44996,27.748587,24.043308,20.341936,16.640562,12.939189,12.622932,12.306676,11.994324,11.678067,11.361811,10.928422,10.491129,10.05774,9.6243515,9.187058,7.656533,6.126007,4.5993857,3.06886,1.5383345,3.416352,5.298274,7.1762915,9.058213,10.936231,9.858616,8.777096,7.6955767,6.617962,5.5364423,6.036206,6.532065,7.0318284,7.5276875,8.023546,7.2582836,6.4969254,5.7316628,4.9663997,4.2011366,4.9781127,5.755089,6.532065,7.309041,8.086017,9.86252,11.639023,13.411622,15.188125,16.960724,16.898252,16.835783,16.773312,16.710842,16.64837,21.236044,25.823717,30.411388,34.99906,39.586735,37.318275,35.045914,32.77746,30.508999,28.236637,28.634886,29.033134,29.431385,29.82573,30.223978,26.354715,22.485453,18.61619,14.743023,10.87376,10.2881,9.706344,9.120684,8.535024,7.9493628,7.3168497,6.6843367,6.0518236,5.4193106,4.786797,4.8687897,4.9468775,5.02887,5.1069584,5.1889505,4.7789884,4.3729305,3.9668727,3.5569105,3.1508527,3.6506162,4.1503797,4.650143,5.1499066,5.64967,5.2943697,4.9351645,4.575959,4.220659,3.8614538,7.6370106,11.408664,15.180316,18.95197,22.723621,20.517633,18.311647,16.101755,13.895767,11.685876,10.651209,9.612638,8.574067,7.5394006,6.5008297,8.886419,11.268105,13.653695,16.039284,18.424873,17.616663,16.808453,16.004145,15.195933,14.387722,15.067088,15.746454,16.42582,17.10909,17.788456,16.675701,15.562947,14.450192,13.337439,12.224684,12.158309,12.091934,12.021654,11.955279,11.888905,13.349152,14.809398,16.26574,17.725986,19.186234,18.167183,17.148134,16.129086,15.1061325,14.087084,13.075843,12.0606985,11.0494585,10.0382185,9.023073,8.898132,8.773191,8.648251,8.52331,8.398369,8.784905,9.171441,9.554072,9.940608,10.323239,10.979179,11.631214,12.28325,12.935285,13.58732,13.048512,12.513609,11.974802,11.435994,10.901091,13.751305,16.601519,19.451733,22.301945,25.148254,24.343948,23.53964,22.735334,21.931028,21.12672,19.685997,18.245272,16.804546,15.363823,13.923099,13.165645,12.408191,11.650736,10.893282,10.135828,8.2226715,6.309514,4.3924527,2.4792955,0.5622339,1.397776,2.233318,3.06886,3.9044023,4.73604,4.7907014,4.841459,4.8961205,4.9468775,5.001539,4.806319,4.6110992,4.415879,4.220659,4.025439,3.7833657,3.5451972,3.3031244,3.0649557,2.8267872,3.7638438,4.704805,5.645766,6.5867267,7.523783,7.277806,7.0318284,6.7819467,6.5359693,6.2860875,5.395884,4.50568,3.619381,2.7291772,1.8389735,1.6945106,1.5539521,1.4094892,1.2689307,1.1244678,0.9058213,0.6910792,0.47243267,0.25378615,0.039044023,0.58175594,1.1205635,1.6632754,2.2059872,2.7486992,2.6354716,2.5183394,2.4051118,2.2918842,2.174752,2.9361105,3.7013733,4.462732,5.22409,5.989353,6.1221027,6.2587566,6.3915067,6.5281606,6.66091,7.7775693,8.894228,10.006983,11.123642,12.236397,13.559989,14.883581,16.20327,17.526861,18.850454,15.84016,12.829865,9.8195715,6.8092775,3.7989833,3.1703746,2.541766,1.9092526,1.2806439,0.6481308,0.7066968,0.76135844,0.8160201,0.8706817,0.92534333,0.81211567,0.698888,0.58566034,0.47633708,0.3631094,0.28892577,0.21864653,0.14446288,0.07418364,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.24597734,0.3513962,0.46071947,0.5661383,0.6754616,0.59346914,0.5153811,0.43338865,0.3553006,0.27330816,0.24597734,0.21864653,0.19131571,0.1639849,0.13665408,0.15617609,0.1717937,0.19131571,0.20693332,0.22645533,0.22255093,0.21864653,0.21864653,0.21474212,0.21083772,0.21083772,0.21083772,0.21083772,0.21083772,0.21083772,0.23816854,0.26940376,0.29673457,0.3240654,0.3513962,0.3357786,0.32016098,0.30454338,0.28892577,0.27330816,0.46071947,0.6442264,0.8316377,1.0151446,1.1986516,1.33921,1.4797685,1.620327,1.7608855,1.901444,1.796025,1.6945106,1.5929961,1.4914817,1.3860629,1.1713207,0.95267415,0.7340276,0.5192855,0.30063897,0.28111696,0.26549935,0.24597734,0.23035973,0.21083772,0.21474212,0.21864653,0.21864653,0.22255093,0.22645533,0.21474212,0.20693332,0.19522011,0.1835069,0.1756981,0.20302892,0.23035973,0.25769055,0.28502136,0.31235218,0.31625658,0.3240654,0.3279698,0.3318742,0.3357786,0.8667773,1.3938715,1.9209659,2.4480603,2.9751544,2.6081407,2.2450314,1.8819219,1.5149081,1.1517987,1.5227169,1.893635,2.2684577,2.639376,3.0141985,3.7521305,4.493967,5.2318993,5.9737353,6.7116675,10.069453,13.427239,16.785025,20.14281,23.500597,23.098444,22.696291,22.294136,21.888079,21.485926,21.38441,21.278992,21.173573,21.068155,20.962736,24.87885,28.791061,32.707176,36.623295,40.53941,39.65311,38.770714,37.88832,37.005924,36.12353,35.213802,34.304077,33.394352,32.484627,31.574902,32.632996,33.691086,34.74918,35.803368,36.86146,58.597267,80.32917,102.06107,123.78907,145.52489,147.16083,148.80067,150.43661,152.07646,153.71242,135.61942,117.52641,99.43341,81.344315,63.251316,53.833897,44.412575,34.99906,25.581644,16.164225,14.34087,12.517513,10.694158,8.870802,7.0513506,6.8092775,6.571109,6.329036,6.0908675,5.8487945,0.5114767,0.5544251,0.59737355,0.64032197,0.6832704,0.7262188,0.737932,0.74964523,0.76135844,0.77307165,0.78868926,0.77307165,0.76135844,0.74964523,0.737932,0.7262188,0.78868926,0.8550641,0.92143893,0.98390937,1.0502841,1.1439898,1.2337911,1.3274968,1.4212024,1.5110037,1.6515622,1.7882162,1.9248703,2.0615244,2.1981785,2.3816853,2.5612879,2.7408905,2.920493,3.1000953,3.310933,3.521771,3.7287042,3.9395418,4.1503797,4.181615,4.2167544,4.2479897,4.279225,4.3143644,4.5017757,4.6930914,4.884407,5.0718184,5.263134,5.169429,5.0757227,4.985922,4.892216,4.7985106,4.6228123,4.4432096,4.267512,4.0918136,3.912211,3.8614538,3.8106966,3.7638438,3.7130866,3.6623292,4.6813784,5.6965227,6.715572,7.7307167,8.749765,9.058213,9.370565,9.679013,9.991365,10.299813,10.6434,10.983084,11.326671,11.6702585,12.013845,11.443803,10.87376,10.303718,9.733675,9.163632,7.7111945,6.2587566,4.806319,3.3538816,1.901444,1.7765031,1.6554666,1.53443,1.4094892,1.2884527,2.3621633,3.435874,4.513489,5.5871997,6.66091,7.703386,8.741957,9.784432,10.823003,11.861574,9.975748,8.093826,6.2079997,4.322173,2.436347,2.5066261,2.5730011,2.639376,2.7057507,2.77603,3.8067923,4.83365,5.8644123,6.8951745,7.9259367,7.5667315,7.2036223,6.844417,6.4852123,6.126007,6.2587566,6.395411,6.5281606,6.6648145,6.801469,6.8639393,6.9264097,6.98888,7.0513506,7.113821,7.426173,7.7385254,8.050878,8.36323,8.675582,8.81614,8.960603,9.101162,9.245625,9.386183,9.175345,8.960603,8.749765,8.538928,8.324185,8.261715,8.19534,8.128965,8.066495,8.00012,9.066022,10.131924,11.193921,12.259823,13.325725,11.213444,9.101162,6.98888,4.8765984,2.7643168,2.5612879,2.3621633,2.1630387,1.9639144,1.7608855,2.0459068,2.3270237,2.6081407,2.893162,3.174279,3.7716527,4.365122,4.958591,5.5559645,6.1494336,6.6335793,7.1216297,7.605776,8.089922,8.574067,10.010887,11.443803,12.880623,14.313539,15.750359,16.32821,16.909966,17.491722,18.069574,18.651329,20.37317,22.095013,23.816854,25.538694,27.26444,29.111223,30.958006,32.804787,34.65157,36.498352,41.784912,47.071472,52.35413,57.64069,62.923347,59.667076,56.410805,53.150627,49.894356,46.638084,43.569225,40.50427,37.43541,34.36655,31.301594,27.377668,23.453745,19.533724,15.6098,11.685876,11.502369,11.318862,11.131451,10.947944,10.760532,10.295909,9.8312845,9.366661,8.902037,8.437413,7.2036223,5.9737353,4.7399445,3.506153,2.2762666,3.408543,4.5408196,5.6730967,6.805373,7.9376497,7.7658563,7.5979667,7.426173,7.2582836,7.08649,7.4144597,7.7424297,8.070399,8.398369,8.726339,7.7892823,6.8561306,5.919074,4.985922,4.0488653,5.2475166,6.446168,7.6409154,8.839567,10.0382185,11.685876,13.337439,14.989,16.636658,18.28822,17.686943,17.085665,16.48829,15.8870125,15.285735,20.298986,25.31224,30.325493,35.338745,40.34809,37.9586,35.5652,33.171803,30.778402,28.388908,28.740305,29.091702,29.443098,29.798397,30.149794,26.534317,22.914936,19.295555,15.680079,12.0606985,11.373524,10.682445,9.991365,9.304191,8.6131115,8.046973,7.47693,6.910792,6.3407493,5.774611,5.8956475,6.016684,6.133816,6.2548523,6.375889,5.919074,5.466163,5.009348,4.5564375,4.0996222,4.376835,4.650143,4.9234514,5.2006636,5.473972,5.4193106,5.364649,5.309987,5.2553253,5.2006636,8.164105,11.131451,14.0948925,17.058334,20.025679,17.593237,15.164699,12.73616,10.303718,7.8751793,8.250002,8.624825,8.999647,9.37447,9.749292,11.0260315,12.306676,13.583415,14.860155,16.136894,15.621513,15.102228,14.586847,14.067561,13.548276,13.981665,14.415053,14.848442,15.281831,15.711315,14.9109125,14.114414,13.314012,12.513609,11.713207,11.541413,11.373524,11.20173,11.033841,10.862047,12.404286,13.94262,15.480955,17.023193,18.56153,17.257458,15.953387,14.649317,13.341343,12.037272,11.639023,11.23687,10.838621,10.436467,10.0382185,10.4637985,10.889378,11.311053,11.736633,12.162213,11.416472,10.666827,9.921086,9.171441,8.4257,9.097258,9.768814,10.444276,11.115833,11.787391,11.799104,11.810817,11.826434,11.838148,11.849861,14.438479,17.023193,19.611813,22.200432,24.78905,24.867138,24.949131,25.027218,25.109211,25.1873,24.191677,23.19215,22.196527,21.197,20.201378,18.495153,16.788929,15.086611,13.380386,11.674163,9.503315,7.328563,5.1577153,2.9868677,0.81211567,1.3509232,1.893635,2.4324427,2.97125,3.513962,3.521771,3.533484,3.541293,3.5530062,3.5608149,3.9083066,4.251894,4.5993857,4.942973,5.2865605,4.6267166,3.9668727,3.3070288,2.6471848,1.9873407,2.822883,3.6584249,4.493967,5.3256044,6.1611466,5.786324,5.407597,5.02887,4.6540475,4.2753205,3.677947,3.0805733,2.4831998,1.8858263,1.2884527,1.2298868,1.1713207,1.116659,1.0580931,0.999527,0.80430686,0.60908675,0.41386664,0.21864653,0.023426414,0.8433509,1.6632754,2.4831998,3.3031244,4.126953,3.9395418,3.7560349,3.5686235,3.3851168,3.2016098,4.025439,4.8492675,5.677001,6.5008297,7.3246584,7.2036223,7.0786815,6.957645,6.8366084,6.7116675,7.422269,8.13287,8.843472,9.554072,10.260769,11.978706,13.692739,15.406772,17.120804,18.838741,16.13299,13.431144,10.729298,8.027451,5.3256044,4.454923,3.5842414,2.7135596,1.8467822,0.97610056,0.9058213,0.8394465,0.77307165,0.7066968,0.63641757,0.61299115,0.58566034,0.5622339,0.5388075,0.5114767,0.40996224,0.30844778,0.20693332,0.10151446,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.20693332,0.29673457,0.39044023,0.48414588,0.57394713,0.5036679,0.43338865,0.3631094,0.29673457,0.22645533,0.20302892,0.1796025,0.15617609,0.13665408,0.113227665,0.13274968,0.15227169,0.1717937,0.19131571,0.21083772,0.21474212,0.21864653,0.21864653,0.22255093,0.22645533,0.23816854,0.24988174,0.26159495,0.27330816,0.28892577,0.3357786,0.38263142,0.42948425,0.47633708,0.5231899,0.49195468,0.45681506,0.42167544,0.38653582,0.3513962,0.5153811,0.679366,0.8433509,1.0112402,1.175225,1.3353056,1.4953861,1.6554666,1.815547,1.9756275,1.815547,1.6554666,1.4953861,1.3353056,1.175225,1.0034313,0.8355421,0.6637484,0.4958591,0.3240654,0.30454338,0.28502136,0.26549935,0.24597734,0.22645533,0.22255093,0.21864653,0.21864653,0.21474212,0.21083772,0.19912452,0.1835069,0.1678893,0.15227169,0.13665408,0.1717937,0.20693332,0.24207294,0.27721256,0.31235218,0.3318742,0.3513962,0.3709182,0.39434463,0.41386664,0.8238289,1.2337911,1.6437533,2.0537157,2.463678,2.1513257,1.8428779,1.53443,1.2220778,0.9136301,1.4290112,1.9443923,2.455869,2.97125,3.4866312,4.0605783,4.630621,5.2045684,5.7785153,6.348558,9.24172,12.134882,15.028045,17.921206,20.81437,20.779228,20.74409,20.70895,20.67381,20.63867,20.38098,20.12329,19.865599,19.607908,19.350218,24.273668,29.19712,34.11667,39.04012,43.96357,42.35886,40.75415,39.14944,37.54083,35.93612,34.159615,32.383114,30.60661,28.826202,27.049698,27.678308,28.310822,28.93943,29.568039,30.200552,45.642464,61.084373,76.52628,91.96819,107.4101,110.10024,112.78647,115.472694,118.16283,120.84906,110.20175,99.55835,88.914955,78.27155,67.624245,57.54308,47.458008,37.376842,27.295675,17.210606,15.274021,13.333533,11.393045,9.452558,7.5120697,7.0513506,6.590631,6.133816,5.6730967,5.212377,0.47633708,0.5388075,0.60518235,0.6715572,0.7340276,0.80040246,0.81211567,0.8238289,0.8394465,0.8511597,0.8628729,0.8394465,0.81211567,0.78868926,0.76135844,0.737932,0.79649806,0.8511597,0.9097257,0.96829176,1.0268579,1.1283722,1.2298868,1.3314011,1.43682,1.5383345,1.6749885,1.8116426,1.9482968,2.0888553,2.2255092,2.3543546,2.4792955,2.6081407,2.7330816,2.8619268,3.193801,3.521771,3.853645,4.181615,4.513489,4.548629,4.5837684,4.618908,4.6540475,4.689187,4.755562,4.825841,4.8961205,4.9663997,5.036679,4.872694,4.7087092,4.5408196,4.376835,4.21285,4.068387,3.9239242,3.775557,3.631094,3.4866312,3.5256753,3.5608149,3.5998588,3.638903,3.6740425,4.814128,5.9542136,7.094299,8.234385,9.37447,9.780528,10.186585,10.588739,10.994797,11.400854,11.502369,11.603884,11.709302,11.810817,11.912332,11.615597,11.318862,11.018223,10.721489,10.424754,8.730244,7.0357327,5.3412223,3.6467118,1.9482968,1.7843118,1.6164225,1.4485333,1.2806439,1.1127546,2.135708,3.1625657,4.1894236,5.212377,6.239235,7.394938,8.550641,9.710248,10.865952,12.025558,10.081166,8.140678,6.196286,4.2557983,2.3114061,2.4402514,2.5690966,2.6940374,2.822883,2.951728,3.978586,5.0054436,6.0323014,7.0591593,8.086017,7.633106,7.1762915,6.7233806,6.266566,5.813655,5.9425,6.0713453,6.2040954,6.3329406,6.461786,6.4500723,6.4383593,6.426646,6.4110284,6.3993154,6.649197,6.899079,7.1489606,7.3988423,7.648724,8.089922,8.531119,8.968412,9.40961,9.850807,9.487698,9.124588,8.761478,8.398369,8.039165,8.39056,8.745861,9.101162,9.456462,9.811763,10.432563,11.053363,11.674163,12.291059,12.911859,10.850334,8.78881,6.7233806,4.661856,2.6003318,2.3621633,2.1239948,1.8858263,1.6515622,1.4133936,1.4992905,1.5812829,1.6671798,1.7530766,1.8389735,2.3855898,2.9322062,3.4788225,4.029343,4.575959,5.1303844,5.6848097,6.239235,6.79366,7.348085,9.128492,10.9089,12.689307,14.469715,16.250122,16.863113,17.48001,18.096905,18.709896,19.326792,21.341463,23.360039,25.378614,27.393286,29.411861,30.544138,31.672512,32.800884,33.93316,35.06153,41.218773,47.372112,53.529354,59.682693,65.83603,62.34159,58.843246,55.344902,51.846558,48.348213,44.908436,41.468655,38.028877,34.5891,31.14932,27.00675,22.86418,18.72161,14.579038,10.436467,10.381805,10.327144,10.272482,10.217821,10.163159,9.6673,9.171441,8.675582,8.183627,7.687768,6.7507114,5.8175592,4.884407,3.9473507,3.0141985,3.39683,3.7833657,4.165997,4.552533,4.939069,5.677001,6.4188375,7.1567693,7.898606,8.636538,8.796618,8.952794,9.108971,9.269051,9.425227,8.320281,7.2153354,6.1103897,5.0054436,3.900498,5.5169206,7.1333427,8.75367,10.370092,11.986515,13.513136,15.035853,16.562475,18.089096,19.611813,18.475632,17.33945,16.199366,15.063184,13.923099,19.36193,24.800762,30.239595,35.674522,41.113358,38.59892,36.084484,33.566147,31.051712,28.537275,28.845724,29.154171,29.458715,29.767162,30.075611,26.710016,23.344421,19.978827,16.613232,13.251541,12.455043,11.6585455,10.865952,10.069453,9.276859,8.773191,8.269524,7.7658563,7.266093,6.7624245,6.9225054,7.082586,7.2426662,7.4027467,7.562827,7.0591593,6.559396,6.055728,5.55206,5.0483923,5.099149,5.1499066,5.2006636,5.251421,5.298274,5.548156,5.794133,6.044015,6.289992,6.5359693,8.695104,10.8542385,13.009468,15.168603,17.323833,14.672744,12.021654,9.366661,6.715572,4.0605783,5.8487945,7.6370106,9.425227,11.213444,13.001659,13.169549,13.341343,13.509232,13.6810255,13.848915,13.622459,13.396004,13.165645,12.939189,12.712734,12.89624,13.083652,13.2671585,13.450665,13.638077,13.150026,12.661977,12.173926,11.685876,11.20173,10.928422,10.655114,10.381805,10.108498,9.839094,11.45942,13.075843,14.69617,16.316498,17.936825,16.347733,14.75864,13.165645,11.576552,9.987461,10.198298,10.413041,10.6238785,10.838621,11.0494585,12.025558,13.001659,13.973856,14.949956,15.926057,14.044135,12.166118,10.284196,8.406178,6.524256,7.2192397,7.910319,8.601398,9.296382,9.987461,10.549695,11.111929,11.674163,12.236397,12.798631,15.125654,17.448774,19.775797,22.098917,24.425941,25.390327,26.354715,27.319103,28.28349,29.251781,28.693453,28.139027,27.584602,27.030176,26.475752,23.820759,21.169668,18.51858,15.863586,13.212498,10.783959,8.351517,5.9229784,3.4905357,1.0619974,1.3079748,1.5539521,1.796025,2.0420024,2.2879796,2.2567444,2.2216048,2.1903696,2.1591344,2.1239948,3.0102942,3.8965936,4.7789884,5.6652875,6.551587,5.4700675,4.388548,3.310933,2.2294137,1.1517987,1.8819219,2.6081407,3.338264,4.068387,4.7985106,4.290938,3.7833657,3.2757936,2.7682211,2.260649,1.9561055,1.6515622,1.3470187,1.0424755,0.737932,0.76526284,0.79259366,0.8199245,0.8472553,0.8745861,0.7027924,0.5309987,0.359205,0.1835069,0.011713207,1.1088502,2.2059872,3.3031244,4.4041657,5.5013027,5.2436123,4.989826,4.73604,4.478349,4.224563,5.1108627,6.001066,6.8873653,7.773665,8.663869,8.281238,7.90251,7.523783,7.141152,6.7624245,7.066968,7.3715115,7.676055,7.9805984,8.289046,10.393518,12.501896,14.610273,16.71865,18.823124,16.429726,14.036326,11.639023,9.245625,6.8483214,5.7394714,4.630621,3.521771,2.4090161,1.3001659,1.1088502,0.92143893,0.7301232,0.5388075,0.3513962,0.41386664,0.47633708,0.5388075,0.60127795,0.6637484,0.5309987,0.39824903,0.26549935,0.13274968,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.1639849,0.24207294,0.32016098,0.39824903,0.47633708,0.41386664,0.3553006,0.29673457,0.23426414,0.1756981,0.15617609,0.14055848,0.12103647,0.10541886,0.08589685,0.10932326,0.13274968,0.15617609,0.1756981,0.19912452,0.20693332,0.21474212,0.22255093,0.23035973,0.23816854,0.26159495,0.28892577,0.31235218,0.3357786,0.3631094,0.42948425,0.4958591,0.5661383,0.63251317,0.698888,0.6442264,0.58956474,0.5349031,0.48024148,0.42557985,0.5700427,0.7145056,0.8589685,1.0034313,1.1517987,1.3314011,1.5110037,1.6906061,1.8702087,2.0498111,1.8311646,1.6164225,1.397776,1.1791295,0.96438736,0.8394465,0.71841,0.59346914,0.47243267,0.3513962,0.3279698,0.30454338,0.28111696,0.26159495,0.23816854,0.23035973,0.22255093,0.21474212,0.20693332,0.19912452,0.1796025,0.16008049,0.14055848,0.12103647,0.10151446,0.14055848,0.1835069,0.22645533,0.26940376,0.31235218,0.3474918,0.38263142,0.41777104,0.45291066,0.48805028,0.78088045,1.0737107,1.3665408,1.6593709,1.9482968,1.6945106,1.4407244,1.1869383,0.92924774,0.6754616,1.3314011,1.9912452,2.6471848,3.3031244,3.9629683,4.369026,4.7711797,5.1772375,5.5832953,5.989353,8.413987,10.8425255,13.271063,15.695697,18.124235,18.45611,18.791887,19.123762,19.455637,19.78751,19.377548,18.967587,18.557625,18.147661,17.7377,23.668486,29.599274,35.526157,41.456944,47.38773,45.060707,42.733685,40.40666,38.07573,35.748707,33.105427,30.458242,27.814962,25.17168,22.524496,22.727526,22.930555,23.133583,23.336613,23.535736,32.69156,41.84348,50.9954,60.147316,69.29923,73.03575,76.77617,80.51268,84.24919,87.9857,84.788,81.590294,78.39649,75.198784,72.00108,61.252262,50.503445,39.75853,29.009708,18.26089,16.20327,14.145649,12.08803,10.034314,7.9766936,7.2934237,6.6140575,5.9346914,5.2553253,4.575959,0.43729305,0.5231899,0.61299115,0.698888,0.78868926,0.8745861,0.8862993,0.9019169,0.9136301,0.92534333,0.93705654,0.9019169,0.8628729,0.8238289,0.78868926,0.74964523,0.80040246,0.8511597,0.9019169,0.94876975,0.999527,1.1127546,1.2259823,1.33921,1.4485333,1.5617609,1.698415,1.8389735,1.9756275,2.1122816,2.2489357,2.3231194,2.4012074,2.475391,2.5495746,2.6237583,3.076669,3.5256753,3.9746814,4.423688,4.8765984,4.911738,4.950782,4.985922,5.024966,5.0640097,5.0132523,4.9624953,4.911738,4.860981,4.814128,4.575959,4.337791,4.0996222,3.8614538,3.6232853,3.513962,3.4007344,3.2875066,3.174279,3.0610514,3.1859922,3.310933,3.435874,3.5608149,3.6857557,4.950782,6.211904,7.47693,8.738052,9.999174,10.498938,10.998701,11.498465,11.998228,12.501896,12.361338,12.224684,12.08803,11.951375,11.810817,11.787391,11.763964,11.736633,11.713207,11.685876,9.749292,7.812709,5.8761253,3.9356375,1.999054,1.7882162,1.5734742,1.3626363,1.1517987,0.93705654,1.9131571,2.8892577,3.8614538,4.8375545,5.813655,7.08649,8.36323,9.636065,10.912805,12.185639,10.186585,8.187531,6.1884775,4.185519,2.1864653,2.3738766,2.5612879,2.7486992,2.9361105,3.1235218,4.1503797,5.173333,6.2001905,7.223144,8.250002,7.699481,7.1489606,6.5984397,6.0518236,5.5013027,5.6262436,5.7511845,5.8761253,6.001066,6.126007,6.036206,5.950309,5.8644123,5.774611,5.688714,5.8761253,6.0635366,6.250948,6.4383593,6.6257706,7.363703,8.101635,8.835662,9.573594,10.311526,9.80005,9.288573,8.773191,8.261715,7.7502384,8.52331,9.300286,10.073358,10.850334,11.623405,11.799104,11.974802,12.150499,12.326198,12.501896,10.487225,8.476458,6.461786,4.4510183,2.436347,2.1630387,1.8858263,1.6125181,1.33921,1.0619974,0.94876975,0.8394465,0.7262188,0.61299115,0.4997635,0.999527,1.4992905,1.999054,2.4988174,2.998581,3.6232853,4.251894,4.8765984,5.5013027,6.126007,8.250002,10.373997,12.501896,14.625891,16.749886,17.40192,18.05005,18.698183,19.350218,19.998348,22.31366,24.625065,26.936472,29.251781,31.563189,31.97315,32.387016,32.800884,33.210846,33.624714,40.64873,47.676655,54.700676,61.724697,68.74872,65.0122,61.27569,57.539177,53.79876,50.062244,46.25155,42.436947,38.62625,34.81165,31.000954,26.635832,22.274614,17.913397,13.548276,9.187058,9.261242,9.339331,9.413514,9.487698,9.561881,9.0386915,8.511597,7.988407,7.461313,6.9381227,6.3017054,5.661383,5.024966,4.388548,3.7482262,3.3890212,3.0259118,2.6628022,2.2996929,1.9365835,3.5881457,5.2358036,6.8873653,8.538928,10.186585,10.174872,10.163159,10.151445,10.135828,10.124115,8.85128,7.57454,6.3017054,5.024966,3.7482262,5.786324,7.824422,9.86252,11.900618,13.938716,15.336493,16.738173,18.135948,19.537628,20.93931,19.26432,17.589333,15.914344,14.239355,12.564366,18.424873,24.285381,30.149794,36.014206,41.874714,39.239243,36.599865,33.96049,31.32502,28.685644,28.951143,29.212738,29.474333,29.735928,30.001427,26.885714,23.773905,20.662096,17.550287,14.438479,13.536563,12.63855,11.736633,10.838621,9.936704,9.499411,9.062118,8.624825,8.187531,7.7502384,7.9493628,8.148487,8.351517,8.550641,8.749765,8.1992445,7.648724,7.098203,6.551587,6.001066,5.825368,5.64967,5.473972,5.298274,5.12648,5.6730967,6.223617,6.774138,7.3246584,7.8751793,9.226103,10.573121,11.924045,13.274967,14.625891,11.748346,8.874706,6.001066,3.1235218,0.24988174,3.4514916,6.649197,9.850807,13.048512,16.250122,15.313066,14.376009,13.438952,12.501896,11.560935,11.623405,11.685876,11.748346,11.810817,11.873287,11.810817,11.748346,11.685876,11.623405,11.560935,11.389141,11.213444,11.037745,10.862047,10.686349,10.311526,9.936704,9.561881,9.187058,8.812236,10.514555,12.212971,13.911386,15.613705,17.31212,15.438006,13.563893,11.685876,9.811763,7.9376497,8.761478,9.589212,10.413041,11.23687,12.0606985,13.58732,15.113941,16.636658,18.163279,19.685997,16.675701,13.661504,10.651209,7.6370106,4.6267166,5.337318,6.0518236,6.7624245,7.47693,8.187531,9.300286,10.413041,11.525795,12.63855,13.751305,15.812829,17.874353,19.935879,22.001307,24.062832,25.913517,27.764204,29.610987,31.461674,33.31236,33.19913,33.085903,32.97658,32.863354,32.750126,29.150267,25.550407,21.95055,18.35069,14.750832,12.0606985,9.37447,6.688241,3.998108,1.3118792,1.261122,1.2142692,1.1635119,1.1127546,1.0619974,0.9878138,0.9136301,0.8394465,0.76135844,0.6871748,2.1122816,3.5373883,4.9624953,6.387602,7.812709,6.3134184,4.814128,3.310933,1.8116426,0.31235218,0.93705654,1.5617609,2.1864653,2.8111696,3.435874,2.7994564,2.1630387,1.5266213,0.8862993,0.24988174,0.23816854,0.22645533,0.21083772,0.19912452,0.18741131,0.30063897,0.41386664,0.5231899,0.63641757,0.74964523,0.60127795,0.44900626,0.30063897,0.14836729,0.0,1.3743496,2.7486992,4.126953,5.5013027,6.8756523,6.551587,6.223617,5.899552,5.575486,5.251421,6.2001905,7.1489606,8.101635,9.050405,9.999174,9.362757,8.726339,8.086017,7.4495993,6.813182,6.7116675,6.6140575,6.5125427,6.4110284,6.3134184,8.812236,11.311053,13.813775,16.312593,18.81141,16.72646,14.637604,12.548749,10.4637985,8.374943,7.0240197,5.6730967,4.3260775,2.9751544,1.6242313,1.3118792,0.999527,0.6871748,0.37482262,0.062470436,0.21083772,0.3631094,0.5114767,0.6637484,0.81211567,0.6481308,0.48805028,0.3240654,0.1639849,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.37482262,0.3240654,0.27330816,0.22645533,0.1756981,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,0.28892577,0.3240654,0.3631094,0.39824903,0.43729305,0.5231899,0.61299115,0.698888,0.78868926,0.8745861,0.80040246,0.7262188,0.6481308,0.57394713,0.4997635,0.62470436,0.74964523,0.8745861,0.999527,1.1244678,1.3235924,1.5266213,1.7257458,1.9248703,2.1239948,1.8506867,1.5734742,1.3001659,1.0268579,0.74964523,0.6754616,0.60127795,0.5231899,0.44900626,0.37482262,0.3513962,0.3240654,0.30063897,0.27330816,0.24988174,0.23816854,0.22645533,0.21083772,0.19912452,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.113227665,0.1639849,0.21083772,0.26159495,0.31235218,0.3631094,0.41386664,0.46071947,0.5114767,0.5622339,0.737932,0.9136301,1.0893283,1.261122,1.43682,1.2376955,1.038571,0.8355421,0.63641757,0.43729305,1.2376955,2.0380979,2.8385005,3.638903,4.4393053,4.6735697,4.911738,5.1499066,5.388075,5.6262436,7.5862536,9.550168,11.514082,13.4740925,15.438006,16.136894,16.835783,17.538574,18.237463,18.936352,18.374117,17.811884,17.24965,16.687416,16.125181,23.063305,30.001427,36.93955,43.873768,50.81189,47.762554,44.713215,41.663876,38.61454,35.561295,32.05124,28.537275,25.023314,21.513256,17.999294,17.776743,17.550287,17.323833,17.101282,16.874826,19.736753,22.59868,25.464512,28.326439,31.188366,35.975163,40.76196,45.548756,50.335552,55.126255,59.374245,63.62614,67.87413,72.12602,76.374016,64.96144,53.548878,42.13631,30.727646,19.311174,17.136421,14.96167,12.786918,10.612165,8.437413,7.535496,6.6374836,5.735567,4.8375545,3.9356375,0.3631094,0.45681506,0.5466163,0.64032197,0.7340276,0.8238289,0.8355421,0.8433509,0.8550641,0.8667773,0.8745861,0.8941081,0.9136301,0.93315214,0.95657855,0.97610056,1.0268579,1.0815194,1.1322767,1.1869383,1.2376955,1.3235924,1.4055848,1.4914817,1.5773785,1.6632754,1.7882162,1.9170616,2.0459068,2.1708477,2.2996929,2.3933985,2.4910088,2.5847144,2.67842,2.77603,3.1157131,3.4593005,3.802888,4.1464753,4.4861584,4.607195,4.728231,4.8492675,4.9663997,5.087436,5.1108627,5.134289,5.153811,5.1772375,5.2006636,4.93126,4.661856,4.388548,4.1191444,3.8497405,3.6935644,3.541293,3.3851168,3.2289407,3.076669,3.240654,3.408543,3.5764325,3.7443218,3.912211,4.9663997,6.0205884,7.0786815,8.13287,9.187058,9.581403,9.971844,10.366188,10.756628,11.150972,11.400854,11.650736,11.900618,12.150499,12.400381,12.322293,12.244205,12.166118,12.091934,12.013845,10.2334385,8.456935,6.6804323,4.903929,3.1235218,2.9634414,2.803361,2.6432803,2.4831998,2.3231194,3.096191,3.8692627,4.6423345,5.4154058,6.1884775,7.238762,8.292951,9.343235,10.397423,11.4516115,9.714153,7.9805984,6.2431393,4.5095844,2.77603,3.0532427,3.3343596,3.6154766,3.8965936,4.173806,4.93126,5.688714,6.446168,7.2036223,7.9610763,7.6721506,7.3832245,7.094299,6.801469,6.5125427,6.6531014,6.7975645,6.9381227,7.082586,7.223144,6.9264097,6.6257706,6.3251314,6.0244927,5.7238536,6.001066,6.278279,6.559396,6.8366084,7.113821,7.918128,8.726339,9.534551,10.342762,11.150972,10.577025,10.003078,9.433036,8.859089,8.289046,9.0035515,9.718058,10.432563,11.147068,11.861574,12.068507,12.2793455,12.486279,12.693212,12.900145,10.862047,8.823949,6.785851,4.7516575,2.7135596,2.4090161,2.1005683,1.796025,1.4914817,1.1869383,1.2415999,1.2962615,1.3509232,1.4055848,1.4641509,1.9131571,2.3621633,2.8111696,3.2640803,3.7130866,4.3026514,4.892216,5.481781,6.0713453,6.66091,8.976221,11.287627,13.599033,15.914344,18.22575,18.72161,19.221373,19.717232,20.21309,20.712854,23.801235,26.885714,29.974096,33.062477,36.15086,35.87365,35.596436,35.31922,35.038105,34.760895,40.801003,46.841114,52.881226,58.921333,64.96144,60.54166,56.12188,51.702095,47.28231,42.86253,39.434464,36.002495,32.57443,29.142458,25.714394,22.36832,19.026152,15.683984,12.341816,8.999647,9.140205,9.280765,9.421323,9.561881,9.698535,9.136301,8.574067,8.011833,7.4495993,6.8873653,6.196286,5.5091114,4.8180323,4.126953,3.435874,3.135235,2.8306916,2.5300527,2.2294137,1.9248703,3.4671092,5.009348,6.551587,8.093826,9.636065,9.593117,9.554072,9.511124,9.468176,9.425227,8.164105,6.899079,5.6379566,4.376835,3.1118085,4.8687897,6.6257706,8.386656,10.143637,11.900618,13.1266,14.356487,15.582469,16.808453,18.038338,17.72989,17.421442,17.1169,16.808453,16.500004,22.770473,29.040943,35.311413,41.581882,47.84845,44.70931,41.566265,38.42322,35.280178,32.137135,30.708124,29.279112,27.846197,26.417185,24.988174,22.844658,20.701141,18.56153,16.41801,14.274494,13.610746,12.950902,12.287154,11.623405,10.963562,10.459893,9.956225,9.456462,8.952794,8.449126,8.433509,8.413987,8.398369,8.378847,8.36323,8.121157,7.882988,7.6409154,7.4027467,7.1606736,6.7663293,6.3719845,5.9776397,5.5832953,5.1889505,6.0791545,6.969358,7.8556576,8.745861,9.636065,11.072885,12.5058,13.94262,15.37944,16.812357,14.192502,11.572648,8.952794,6.3329406,3.7130866,5.8487945,7.9805984,10.116306,12.252014,14.387722,13.743496,13.09927,12.4511385,11.806912,11.162686,11.037745,10.912805,10.787864,10.662923,10.537982,10.471607,10.409137,10.342762,10.276386,10.213917,10.241247,10.272482,10.303718,10.331048,10.362284,10.167064,9.971844,9.776623,9.581403,9.386183,10.467703,11.549222,12.626837,13.708356,14.785972,13.349152,11.912332,10.475512,9.0386915,7.601871,8.265619,8.929368,9.593117,10.260769,10.924518,13.938716,16.94901,19.96321,22.973503,25.987701,22.75876,19.525915,16.296974,13.068034,9.839094,9.675109,9.511124,9.351044,9.187058,9.023073,9.671205,10.315431,10.959657,11.603884,12.24811,14.621986,16.995863,19.365835,21.739712,24.113588,25.866665,27.623646,29.376722,31.133703,32.88678,32.262077,31.637371,31.012667,30.387962,29.763258,28.021894,26.284435,24.543072,22.801708,21.06425,17.421442,13.778636,10.135828,6.493021,2.8502135,2.803361,2.7565079,2.7057507,2.6588979,2.612045,2.5495746,2.4871042,2.4246337,2.3621633,2.2996929,3.1703746,4.041056,4.911738,5.7785153,6.649197,5.493494,4.3338866,3.1781836,2.018576,0.8628729,1.3665408,1.8663043,2.3699722,2.87364,3.3734035,2.9751544,2.5769055,2.174752,1.7765031,1.3743496,1.2142692,1.0502841,0.8862993,0.7262188,0.5622339,0.57785153,0.59346914,0.60908675,0.62079996,0.63641757,0.5349031,0.43338865,0.3318742,0.22645533,0.12494087,1.261122,2.3933985,3.5295796,4.6657605,5.801942,5.6145306,5.4310236,5.2436123,5.0601053,4.8765984,5.571582,6.27047,6.969358,7.6643414,8.36323,7.7814736,7.2036223,6.621866,6.044015,5.462259,5.3841705,5.3021784,5.22409,5.142098,5.0640097,7.0591593,9.058213,11.053363,13.052417,15.051471,13.614651,12.181735,10.744915,9.308095,7.8751793,6.715572,5.559869,4.4041657,3.2445583,2.0888553,1.678893,1.2728351,0.8667773,0.45681506,0.05075723,0.19522011,0.339683,0.48414588,0.62860876,0.77307165,0.62079996,0.46462387,0.30844778,0.15617609,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.10151446,0.15617609,0.20693332,0.26159495,0.31235218,0.27330816,0.23426414,0.19131571,0.15227169,0.113227665,0.10932326,0.10151446,0.09761006,0.093705654,0.08589685,0.10932326,0.12884527,0.14836729,0.1678893,0.18741131,0.21083772,0.23816854,0.26159495,0.28892577,0.31235218,0.3474918,0.38263142,0.41777104,0.45291066,0.48805028,0.5544251,0.61689556,0.6832704,0.74574083,0.81211567,0.7418364,0.6676528,0.59346914,0.5231899,0.44900626,0.5388075,0.62860876,0.71841,0.80821127,0.9019169,1.0815194,1.261122,1.4407244,1.620327,1.7999294,1.5969005,1.3899672,1.1869383,0.98000497,0.77307165,0.7027924,0.62860876,0.5583295,0.48414588,0.41386664,0.38653582,0.359205,0.3318742,0.30063897,0.27330816,0.26940376,0.26159495,0.25378615,0.24597734,0.23816854,0.20693332,0.1717937,0.14055848,0.10932326,0.07418364,0.11713207,0.16008049,0.20302892,0.24597734,0.28892577,0.3279698,0.3670138,0.40605783,0.44900626,0.48805028,0.6481308,0.80821127,0.96829176,1.1283722,1.2884527,1.1517987,1.0112402,0.8745861,0.737932,0.60127795,1.261122,1.9248703,2.5886188,3.2484627,3.912211,4.2557983,4.5993857,4.939069,5.282656,5.6262436,7.0903945,8.554545,10.018696,11.486752,12.950902,14.008995,15.067088,16.121277,17.17937,18.237463,17.909492,17.581524,17.253553,16.925583,16.601519,23.047686,29.493855,35.943928,42.390095,48.83626,46.08366,43.331055,40.578453,37.825848,35.073246,32.437775,29.798397,27.162926,24.52355,21.888079,20.76361,19.643047,18.51858,17.398016,16.273548,18.573242,20.86903,23.168722,25.464512,27.764204,32.289406,36.818512,41.343716,45.87282,50.401928,53.748,57.094074,60.44405,63.790123,67.1362,57.36348,47.59076,37.81804,28.049225,18.276506,16.367254,14.458001,12.552653,10.6434,8.738052,8.234385,7.7307167,7.230953,6.727285,6.223617,0.28892577,0.38653582,0.48414588,0.58175594,0.679366,0.77307165,0.78088045,0.78868926,0.79649806,0.80430686,0.81211567,0.8902037,0.96829176,1.0463798,1.1205635,1.1986516,1.2533131,1.3118792,1.3665408,1.4212024,1.475864,1.53443,1.5890918,1.6476578,1.7062237,1.7608855,1.8819219,1.999054,2.1161861,2.233318,2.35045,2.463678,2.5808098,2.6940374,2.8111696,2.9243972,3.1586614,3.39683,3.631094,3.8653584,4.0996222,4.3026514,4.50568,4.7087092,4.911738,5.1108627,5.2084727,5.3021784,5.395884,5.493494,5.5871997,5.2865605,4.9820175,4.6813784,4.376835,4.0761957,3.8770714,3.6818514,3.4827268,3.2836022,3.0883822,3.2992198,3.506153,3.716991,3.9278288,4.138666,4.985922,5.833177,6.6804323,7.5276875,8.374943,8.659965,8.944985,9.230007,9.515028,9.80005,10.436467,11.076789,11.713207,12.349625,12.986042,12.857197,12.728352,12.595602,12.466757,12.337912,10.721489,9.101162,7.4847393,5.8683167,4.251894,4.142571,4.0332475,3.9278288,3.8185053,3.7130866,4.283129,4.853172,5.423215,5.9932575,6.5633,7.3910336,8.2226715,9.054309,9.882042,10.71368,9.24172,7.773665,6.3017054,4.83365,3.3616903,3.736513,4.1074314,4.478349,4.853172,5.22409,5.716045,6.2040954,6.6960497,7.1841,7.676055,7.6448197,7.6135845,7.5862536,7.5550184,7.523783,7.6838636,7.843944,8.0040245,8.164105,8.324185,7.812709,7.3012323,6.785851,6.2743745,5.7628975,6.1299114,6.4969254,6.8639393,7.230953,7.601871,8.476458,9.354948,10.2334385,11.111929,11.986515,11.354002,10.721489,10.088976,9.456462,8.823949,9.479889,10.135828,10.791768,11.443803,12.099743,12.341816,12.579984,12.818152,13.0602255,13.298394,11.23687,9.175345,7.113821,5.0483923,2.9868677,2.6510892,2.3192148,1.9834363,1.6476578,1.3118792,1.53443,1.756981,1.979532,2.2020829,2.4246337,2.8267872,3.2250361,3.6232853,4.025439,4.423688,4.9781127,5.5364423,6.0908675,6.6452928,7.1997175,9.698535,12.201257,14.700074,17.198893,19.701614,20.0452,20.388788,20.73628,21.079868,21.423454,25.288813,29.150267,33.011723,36.873177,40.738533,39.77024,38.80195,37.833656,36.86927,35.900978,40.953274,46.009476,51.065678,56.12188,61.174175,56.07112,50.97197,45.86892,40.765865,35.66281,32.613472,29.568039,26.5187,23.473267,20.423927,18.10081,15.781594,13.458474,11.135355,8.812236,9.019169,9.2221985,9.4291315,9.63216,9.839094,9.237816,8.636538,8.039165,7.437886,6.8366084,6.094772,5.3529353,4.6110992,3.8692627,3.1235218,2.8814487,2.639376,2.397303,2.15523,1.9131571,3.3460727,4.7828927,6.2158084,7.6526284,9.089449,9.0152645,8.941081,8.870802,8.796618,8.726339,7.47693,6.223617,4.9742084,3.7247996,2.475391,3.951255,5.4310236,6.9068875,8.386656,9.86252,10.916709,11.970898,13.028991,14.0831785,15.137367,16.199366,17.257458,18.319456,19.377548,20.435642,27.116074,33.792603,40.469128,47.149563,53.826088,50.17938,46.528763,42.88205,39.23534,35.588627,32.465103,29.341583,26.218061,23.098444,19.974922,18.8036,17.628376,16.457056,15.285735,14.114414,13.688834,13.263254,12.837675,12.412095,11.986515,11.420377,10.8542385,10.284196,9.718058,9.151918,8.913751,8.679486,8.445222,8.210958,7.9766936,8.043069,8.113348,8.183627,8.253906,8.324185,7.7111945,7.094299,6.481308,5.8644123,5.251421,6.481308,7.7111945,8.941081,10.170968,11.400854,12.919667,14.438479,15.961197,17.48001,18.998821,16.636658,14.27059,11.904523,9.538455,7.1762915,8.246098,9.315904,10.38571,11.455516,12.525322,12.173926,11.818625,11.46723,11.115833,10.764437,10.44818,10.135828,9.823476,9.511124,9.198771,9.132397,9.066022,8.995743,8.929368,8.862993,9.097258,9.331521,9.565785,9.803954,10.0382185,10.0226,10.006983,9.991365,9.975748,9.964035,10.42085,10.881569,11.342289,11.803008,12.263727,11.2642,10.260769,9.261242,8.261715,7.262188,7.7658563,8.273428,8.777096,9.280765,9.788337,14.286208,18.787983,23.285854,27.78763,32.289406,28.837915,25.394232,21.946646,18.499058,15.051471,14.012899,12.974329,11.935758,10.901091,9.86252,10.0382185,10.217821,10.393518,10.573121,10.748819,13.431144,16.113468,18.795792,21.478117,24.164345,25.823717,27.483088,29.142458,30.80183,32.4612,31.32502,30.188839,29.048752,27.91257,26.77639,26.893522,27.014559,27.135595,27.256632,27.373764,22.778282,18.178898,13.583415,8.98403,4.388548,4.3416953,4.298747,4.251894,4.2089458,4.1620927,4.1113358,4.0605783,4.0137253,3.9629683,3.912211,4.2284675,4.5408196,4.8570766,5.173333,5.4856853,4.6735697,3.8575494,3.0415294,2.2294137,1.4133936,1.7921207,2.1708477,2.5534792,2.9322062,3.310933,3.1508527,2.9868677,2.8267872,2.6628022,2.4988174,2.1864653,1.8741131,1.5617609,1.2494087,0.93705654,0.8550641,0.77307165,0.6910792,0.60908675,0.5231899,0.46852827,0.41386664,0.359205,0.30454338,0.24988174,1.1439898,2.0380979,2.9361105,3.8302186,4.7243266,4.6813784,4.6345253,4.591577,4.5447245,4.5017757,4.9468775,5.388075,5.833177,6.278279,6.7233806,6.2040954,5.6809053,5.1577153,4.6345253,4.1113358,4.0527697,3.9942036,3.9317331,3.873167,3.8106966,5.3060827,6.801469,8.296855,9.792241,11.287627,10.506746,9.721962,8.941081,8.156297,7.375416,6.4110284,5.446641,4.478349,3.513962,2.5495746,2.0459068,1.5461433,1.0424755,0.5388075,0.039044023,0.1756981,0.31625658,0.45681506,0.59737355,0.737932,0.58956474,0.44119745,0.29673457,0.14836729,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.078088045,0.12103647,0.1639849,0.20693332,0.24988174,0.21864653,0.19131571,0.16008049,0.12884527,0.10151446,0.10151446,0.10541886,0.10932326,0.10932326,0.113227665,0.12884527,0.14055848,0.15617609,0.1717937,0.18741131,0.22645533,0.26159495,0.30063897,0.3357786,0.37482262,0.40605783,0.44119745,0.47243267,0.5036679,0.5388075,0.58175594,0.62079996,0.6637484,0.7066968,0.74964523,0.679366,0.60908675,0.5388075,0.46852827,0.39824903,0.45681506,0.5114767,0.5661383,0.62079996,0.6754616,0.8355421,0.9956226,1.1557031,1.3157835,1.475864,1.33921,1.2064602,1.0698062,0.93315214,0.80040246,0.7301232,0.659844,0.58956474,0.5192855,0.44900626,0.42167544,0.39044023,0.359205,0.3318742,0.30063897,0.29673457,0.29673457,0.29283017,0.28892577,0.28892577,0.24597734,0.20693332,0.1678893,0.12884527,0.08589685,0.12103647,0.15617609,0.19131571,0.22645533,0.26159495,0.29283017,0.3240654,0.3513962,0.38263142,0.41386664,0.5583295,0.7027924,0.8472553,0.9917182,1.1361811,1.0619974,0.9878138,0.9136301,0.8394465,0.76135844,1.2884527,1.8116426,2.338737,2.8619268,3.3890212,3.8341231,4.283129,4.728231,5.1772375,5.6262436,6.590631,7.558923,8.527214,9.495506,10.4637985,11.877192,13.29449,14.707883,16.121277,17.538574,17.44487,17.351164,17.261362,17.167656,17.073952,23.032068,28.990187,34.948303,40.90642,46.860638,44.408672,41.9528,39.496933,37.041065,34.5891,32.82431,31.063425,29.298634,27.537748,25.776863,23.754383,21.735807,19.713327,17.694752,15.676175,17.405825,19.13938,20.872934,22.60649,24.33614,28.603651,32.871162,37.138676,41.406185,45.6737,48.121758,50.565914,53.01007,55.454224,57.89838,49.76551,41.63264,33.503677,25.370806,17.237936,15.598087,13.958238,12.318389,10.67854,9.0386915,8.933272,8.827853,8.722435,8.617016,8.511597,0.21083772,0.31625658,0.41777104,0.5192855,0.62079996,0.7262188,0.7301232,0.7340276,0.7418364,0.74574083,0.74964523,0.8862993,1.0190489,1.1557031,1.2884527,1.4251068,1.4836729,1.5383345,1.5969005,1.6554666,1.7140326,1.7413634,1.7725986,1.8038338,1.8311646,1.8623998,1.9717231,2.077142,2.1864653,2.2918842,2.4012074,2.533957,2.6706111,2.803361,2.9400148,3.076669,3.2016098,3.330455,3.4593005,3.5842414,3.7130866,3.998108,4.283129,4.5681505,4.853172,5.138193,5.3060827,5.473972,5.6418614,5.805846,5.9737353,5.6418614,5.3060827,4.970304,4.6345253,4.298747,4.0605783,3.8185053,3.5803368,3.338264,3.1000953,3.3538816,3.6037633,3.8575494,4.1113358,4.3612175,5.001539,5.6418614,6.282183,6.9225054,7.562827,7.7385254,7.918128,8.093826,8.273428,8.449126,9.475985,10.498938,11.525795,12.548749,13.575606,13.392099,13.208592,13.028991,12.845484,12.661977,11.205634,9.749292,8.289046,6.832704,5.376362,5.3217,5.263134,5.2084727,5.153811,5.099149,5.466163,5.833177,6.2040954,6.571109,6.9381227,7.5433054,8.152391,8.761478,9.366661,9.975748,8.769287,7.5667315,6.3602715,5.153811,3.951255,4.415879,4.8805027,5.3451266,5.8097506,6.2743745,6.4969254,6.719476,6.942027,7.164578,7.387129,7.617489,7.8478484,8.078208,8.308568,8.538928,8.714626,8.894228,9.069926,9.245625,9.425227,8.699008,7.9766936,7.250475,6.524256,5.801942,6.2587566,6.715572,7.172387,7.629202,8.086017,9.034787,9.983557,10.928422,11.877192,12.825961,12.130978,11.4398985,10.748819,10.053836,9.362757,9.956225,10.553599,11.147068,11.744442,12.337912,12.611219,12.880623,13.153932,13.427239,13.700547,11.611692,9.526741,7.437886,5.349031,3.2640803,2.8970666,2.533957,2.1669433,1.8038338,1.43682,1.8272603,2.2177005,2.6081407,2.998581,3.3890212,3.736513,4.087909,4.4393053,4.786797,5.138193,5.657479,6.1767645,6.6960497,7.2192397,7.7385254,10.424754,13.110983,15.801116,18.487345,21.173573,21.368793,21.56011,21.751425,21.946646,22.13796,26.77639,31.410915,36.049347,40.687775,45.326206,43.666836,42.011368,40.351997,38.69653,37.03716,41.105545,45.177837,49.246227,53.318516,57.386906,51.60058,45.81816,40.031837,34.245514,28.463093,25.796385,23.133583,20.466877,17.804073,15.137367,13.833297,12.533132,11.229061,9.928895,8.624825,8.894228,9.163632,9.43694,9.706344,9.975748,9.339331,8.699008,8.062591,7.426173,6.785851,5.9932575,5.196759,4.4041657,3.6076677,2.8111696,2.631567,2.4480603,2.2645533,2.0810463,1.901444,3.2289407,4.5564375,5.883934,7.211431,8.538928,8.433509,8.331994,8.23048,8.128965,8.023546,6.785851,5.548156,4.3143644,3.076669,1.8389735,3.0337205,4.2323723,5.4310236,6.6257706,7.824422,8.706817,9.589212,10.471607,11.354002,12.236397,14.664935,17.093473,19.52201,21.946646,24.375183,31.461674,38.54426,45.63075,52.713333,59.799824,55.649445,51.495163,47.340878,43.1905,39.036213,34.222084,29.407957,24.59383,19.775797,14.96167,14.75864,14.555612,14.356487,14.153459,13.950429,13.763018,13.575606,13.388195,13.200784,13.013372,12.380859,11.748346,11.115833,10.48332,9.850807,9.397896,8.944985,8.492075,8.039165,7.5862536,7.968885,8.347612,8.726339,9.108971,9.487698,8.652155,7.816613,6.9810715,6.1494336,5.3138914,6.883461,8.453031,10.0226,11.592171,13.16174,14.766449,16.371159,17.975868,19.584482,21.189192,19.07691,16.968533,14.856251,12.747873,10.639496,10.6434,10.647305,10.651209,10.6590185,10.662923,10.604357,10.541886,10.48332,10.42085,10.362284,9.86252,9.362757,8.862993,8.36323,7.8634663,7.793187,7.7229075,7.6526284,7.5823493,7.5120697,7.9532676,8.39056,8.831758,9.272955,9.714153,9.878138,10.042123,10.206107,10.373997,10.537982,10.377901,10.217821,10.05774,9.897659,9.737579,9.175345,8.6131115,8.050878,7.4886436,6.9264097,7.269997,7.6135845,7.9610763,8.304664,8.648251,14.637604,20.623053,26.612406,32.601757,38.587208,34.920975,31.258644,27.592411,23.926178,20.263847,18.35069,16.437534,14.524376,12.611219,10.701966,10.409137,10.120211,9.8312845,9.538455,9.249529,12.244205,15.234978,18.22575,21.220427,24.211199,25.776863,27.34253,28.908194,30.47386,32.03562,30.387962,28.7364,27.088743,25.437181,23.785618,25.769054,27.748587,29.728119,31.707651,33.687183,28.135122,22.583063,17.031002,11.478943,5.9268827,5.883934,5.840986,5.7980375,5.755089,5.7121406,5.6730967,5.6379566,5.5989127,5.563773,5.5247293,5.2865605,5.044488,4.806319,4.564246,4.3260775,3.853645,3.3812122,2.9087796,2.436347,1.9639144,2.2216048,2.4792955,2.7330816,2.9907722,3.2484627,3.3265507,3.4007344,3.474918,3.5491016,3.6232853,3.1625657,2.7018464,2.2372224,1.7765031,1.3118792,1.1322767,0.95267415,0.77307165,0.59346914,0.41386664,0.40605783,0.39824903,0.39044023,0.38263142,0.37482262,1.0307622,1.6867018,2.338737,2.9946766,3.6506162,3.7443218,3.8380275,3.9356375,4.029343,4.123049,4.318269,4.5095844,4.7009,4.8961205,5.087436,4.6228123,4.1581883,3.6935644,3.2289407,2.7643168,2.7213683,2.6823244,2.6432803,2.6042364,2.5612879,3.5569105,4.548629,5.5403466,6.532065,7.523783,7.394938,7.266093,7.1333427,7.0044975,6.8756523,6.1025805,5.3295093,4.5564375,3.7833657,3.0141985,2.416825,1.8194515,1.2181735,0.62079996,0.023426414,0.16008049,0.29673457,0.42948425,0.5661383,0.698888,0.5583295,0.42167544,0.28111696,0.14055848,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.058566034,0.08980125,0.12103647,0.15617609,0.18741131,0.1678893,0.14836729,0.12884527,0.10932326,0.08589685,0.09761006,0.10932326,0.11713207,0.12884527,0.13665408,0.14836729,0.15617609,0.1678893,0.1756981,0.18741131,0.23816854,0.28892577,0.3357786,0.38653582,0.43729305,0.46852827,0.4958591,0.5270943,0.5583295,0.58566034,0.60908675,0.62860876,0.6481308,0.6676528,0.6871748,0.62079996,0.5544251,0.48414588,0.41777104,0.3513962,0.3709182,0.39044023,0.40996224,0.42948425,0.44900626,0.58956474,0.7301232,0.8706817,1.0112402,1.1517987,1.0854238,1.0190489,0.95657855,0.8902037,0.8238289,0.75745404,0.6910792,0.62079996,0.5544251,0.48805028,0.45681506,0.42167544,0.39044023,0.359205,0.3240654,0.3279698,0.3318742,0.3318742,0.3357786,0.3357786,0.28892577,0.24207294,0.19522011,0.14836729,0.10151446,0.12884527,0.15617609,0.1835069,0.21083772,0.23816854,0.25769055,0.27721256,0.29673457,0.31625658,0.3357786,0.46852827,0.59737355,0.7262188,0.8589685,0.9878138,0.97610056,0.96438736,0.94876975,0.93705654,0.92534333,1.3118792,1.698415,2.0888553,2.475391,2.8619268,3.416352,3.9668727,4.521298,5.0718184,5.6262436,6.094772,6.5633,7.0357327,7.504261,7.9766936,9.749292,11.521891,13.2905855,15.063184,16.835783,16.980246,17.120804,17.265266,17.405825,17.550287,23.01645,28.486519,33.952682,39.418846,44.888912,42.72978,40.570644,38.415413,36.25628,34.101048,33.210846,32.324547,31.438248,30.551949,29.661743,26.745155,23.828568,20.908073,17.991486,15.074897,16.242313,17.409729,18.577147,19.744562,20.911978,24.921799,28.927717,32.93363,36.943455,40.94937,42.49161,44.033848,45.576088,47.11833,48.660564,42.167545,35.67843,29.185408,22.692387,16.199366,14.828919,13.45457,12.084125,10.709775,9.339331,9.628256,9.921086,10.213917,10.506746,10.799577,0.13665408,0.24597734,0.3513962,0.46071947,0.5661383,0.6754616,0.679366,0.679366,0.6832704,0.6832704,0.6871748,0.8784905,1.0737107,1.2650263,1.456342,1.6515622,1.7101282,1.7686942,1.8311646,1.8897307,1.9482968,1.9522011,1.9561055,1.9561055,1.9600099,1.9639144,2.0615244,2.1591344,2.2567444,2.3543546,2.4480603,2.6042364,2.7604125,2.9165885,3.06886,3.2250361,3.2445583,3.2640803,3.2836022,3.3031244,3.3265507,3.6935644,4.0605783,4.4275923,4.794606,5.1616197,5.4036927,5.6418614,5.883934,6.1221027,6.364176,5.9932575,5.6262436,5.2592297,4.892216,4.5252023,4.2440853,3.959064,3.677947,3.39683,3.1118085,3.408543,3.7013733,3.998108,4.290938,4.5876727,5.0210614,5.4505453,5.883934,6.3173227,6.7507114,6.8209906,6.89127,6.9615493,7.0318284,7.098203,8.511597,9.924991,11.338385,12.751778,14.161267,13.927003,13.692739,13.458474,13.224211,12.986042,11.68978,10.393518,9.093353,7.7970915,6.5008297,6.4969254,6.4969254,6.493021,6.4891167,6.4891167,6.6531014,6.817086,6.9810715,7.1489606,7.3129454,7.6955767,8.082112,8.468649,8.85128,9.237816,8.296855,7.355894,6.4188375,5.477876,4.5369153,5.095245,5.6535745,6.211904,6.7663293,7.3246584,7.28171,7.2348576,7.191909,7.1450562,7.098203,7.590158,8.078208,8.570163,9.058213,9.550168,9.745388,9.940608,10.135828,10.331048,10.526268,9.589212,8.648251,7.7111945,6.774138,5.8370814,6.3836975,6.9342184,7.480835,8.027451,8.574067,9.593117,10.608261,11.62731,12.6463585,13.661504,12.911859,12.158309,11.404759,10.651209,9.901564,10.436467,10.971371,11.506273,12.041177,12.576079,12.880623,13.185166,13.48971,13.794253,14.098797,11.986515,9.874233,7.7619514,5.64967,3.5373883,3.1430438,2.7486992,2.3543546,1.9561055,1.5617609,2.1200905,2.67842,3.2367494,3.7911747,4.349504,4.650143,4.950782,5.251421,5.548156,5.8487945,6.336845,6.8209906,7.3051367,7.7892823,8.273428,11.150972,14.024612,16.898252,19.775797,22.649437,22.688482,22.73143,22.770473,22.809519,22.848562,28.263968,33.67547,39.08697,44.498474,49.91388,47.563427,45.21688,42.87034,40.523792,38.17334,41.261723,44.3462,47.43068,50.515156,53.599632,47.133945,40.66435,34.198658,27.729065,21.263374,18.9793,16.69913,14.415053,12.130978,9.850807,9.565785,9.284669,9.0035515,8.718531,8.437413,8.773191,9.108971,9.440845,9.776623,10.112402,9.43694,8.761478,8.086017,7.4105554,6.7389984,5.891743,5.040583,4.193328,3.3460727,2.4988174,2.377781,2.2567444,2.1318035,2.0107672,1.8858263,3.1079042,4.3260775,5.548156,6.7663293,7.988407,7.8556576,7.7229075,7.590158,7.4574084,7.3246584,6.098676,4.8765984,3.6506162,2.4246337,1.1986516,2.1161861,3.0337205,3.951255,4.8687897,5.786324,6.4969254,7.2075267,7.918128,8.628729,9.339331,13.130505,16.925583,20.724567,24.515741,28.310822,35.803368,43.295918,50.788464,58.281013,65.77356,61.119514,56.46156,51.803608,47.145657,42.487705,35.979065,29.474333,22.965694,16.457056,9.948417,10.717585,11.486752,12.252014,13.021181,13.786445,13.837202,13.887959,13.938716,13.985569,14.036326,13.341343,12.642454,11.943566,11.248583,10.549695,9.878138,9.2104845,8.538928,7.871275,7.1997175,7.890797,8.581876,9.269051,9.96013,10.651209,9.593117,8.538928,7.4847393,6.4305506,5.376362,7.2856145,9.194867,11.10412,13.013372,14.92653,16.613232,18.303837,19.994444,21.685051,23.375656,21.521065,19.666473,17.811884,15.953387,14.098797,13.040704,11.978706,10.920613,9.858616,8.800523,9.030883,9.265146,9.499411,9.729771,9.964035,9.276859,8.58578,7.898606,7.211431,6.524256,6.453977,6.379793,6.3056097,6.2353306,6.1611466,6.8092775,7.453504,8.097731,8.741957,9.386183,9.733675,10.077262,10.42085,10.768341,11.111929,10.331048,9.554072,8.773191,7.9923115,7.211431,7.08649,6.9615493,6.8366084,6.7116675,6.5867267,6.774138,6.957645,7.141152,7.328563,7.5120697,14.989,22.462027,29.938957,37.411983,44.888912,41.004032,37.12306,33.23818,29.3572,25.476225,22.688482,19.900738,17.112995,14.325252,11.537509,10.780055,10.0226,9.265146,8.507692,7.7502384,11.053363,14.356487,17.655706,20.958832,24.261955,25.733915,27.201971,28.673931,30.141985,31.613945,29.450907,27.287867,25.124828,22.96179,20.79875,24.640682,28.47871,32.32064,36.15867,40.000603,33.491962,26.983324,20.47859,13.969952,7.461313,7.422269,7.3832245,7.3441806,7.3012323,7.262188,7.238762,7.211431,7.1880045,7.1606736,7.137247,6.3407493,5.548156,4.7516575,3.959064,3.1625657,3.0337205,2.900971,2.7721257,2.6432803,2.514435,2.6471848,2.7838387,2.9165885,3.0532427,3.1859922,3.4983444,3.8106966,4.126953,4.4393053,4.7516575,4.138666,3.5256753,2.912684,2.2996929,1.6867018,1.4094892,1.1322767,0.8550641,0.57785153,0.30063897,0.339683,0.37872702,0.42167544,0.46071947,0.4997635,0.9136301,1.3314011,1.7452679,2.1591344,2.5769055,2.8111696,3.0454338,3.279698,3.513962,3.7482262,3.68966,3.631094,3.5686235,3.5100577,3.4514916,3.0415294,2.6354716,2.2294137,1.8194515,1.4133936,1.3938715,1.3743496,1.3509232,1.3314011,1.3118792,1.8038338,2.2918842,2.7838387,3.2718892,3.7638438,4.283129,4.806319,5.3295093,5.852699,6.375889,5.794133,5.2162814,4.6345253,4.056674,3.474918,2.7838387,2.0888553,1.397776,0.7066968,0.011713207,0.14055848,0.27330816,0.40215343,0.5309987,0.6637484,0.5309987,0.39824903,0.26549935,0.13274968,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.03513962,0.058566034,0.078088045,0.10151446,0.12494087,0.113227665,0.10541886,0.093705654,0.08589685,0.07418364,0.093705654,0.10932326,0.12884527,0.14446288,0.1639849,0.1678893,0.1717937,0.1756981,0.1835069,0.18741131,0.24988174,0.31235218,0.37482262,0.43729305,0.4997635,0.5270943,0.5544251,0.58175594,0.60908675,0.63641757,0.63641757,0.63251317,0.62860876,0.62860876,0.62470436,0.5583295,0.4958591,0.42948425,0.3631094,0.30063897,0.28502136,0.26940376,0.25378615,0.23816854,0.22645533,0.3435874,0.46462387,0.58566034,0.7066968,0.8238289,0.8316377,0.8355421,0.8394465,0.8433509,0.8511597,0.78478485,0.71841,0.6559396,0.58956474,0.5231899,0.48805028,0.45681506,0.42167544,0.38653582,0.3513962,0.359205,0.3631094,0.3709182,0.37872702,0.38653582,0.3318742,0.27721256,0.22255093,0.1678893,0.113227665,0.13274968,0.15227169,0.1717937,0.19131571,0.21083772,0.22255093,0.23426414,0.24207294,0.25378615,0.26159495,0.37872702,0.49195468,0.60908675,0.7223144,0.8394465,0.8862993,0.93705654,0.9878138,1.038571,1.0893283,1.33921,1.5890918,1.8389735,2.0888553,2.338737,2.9946766,3.6506162,4.31046,4.9663997,5.6262436,5.5989127,5.571582,5.5442514,5.5169206,5.4856853,7.617489,9.749292,11.877192,14.008995,16.136894,16.515621,16.894348,17.26917,17.647898,18.026625,23.004738,27.978947,32.957058,37.935173,42.913284,41.050884,39.19239,37.333893,35.471493,33.613,33.601284,33.585667,33.573956,33.56224,33.55053,29.735928,25.921326,22.106726,18.292124,14.473619,15.078801,15.680079,16.281357,16.88654,17.487818,21.236044,24.98427,28.728592,32.476818,36.225044,36.865368,37.505688,38.14601,38.78633,39.426655,34.573483,29.72031,24.867138,20.013966,15.160794,14.055848,12.950902,11.845957,10.741011,9.636065,10.327144,11.018223,11.709302,12.396477,13.087557,0.062470436,0.1756981,0.28892577,0.39824903,0.5114767,0.62470436,0.62470436,0.62470436,0.62470436,0.62470436,0.62470436,0.8745861,1.1244678,1.3743496,1.6242313,1.8741131,1.9365835,1.999054,2.0615244,2.1239948,2.1864653,2.1630387,2.135708,2.1122816,2.0888553,2.0615244,2.1513257,2.2372224,2.3231194,2.4129205,2.4988174,2.6745155,2.8502135,3.0259118,3.2016098,3.3734035,3.2875066,3.2016098,3.1118085,3.0259118,2.9361105,3.3890212,3.8380275,4.2870336,4.73604,5.1889505,5.5013027,5.813655,6.126007,6.4383593,6.7507114,6.348558,5.950309,5.548156,5.1499066,4.7516575,4.423688,4.0996222,3.775557,3.4514916,3.1235218,3.4632049,3.7989833,4.138666,4.474445,4.814128,5.036679,5.263134,5.4856853,5.7121406,5.938596,5.899552,5.8644123,5.825368,5.786324,5.7511845,7.551114,9.351044,11.150972,12.950902,14.750832,14.461906,14.176885,13.887959,13.599033,13.314012,12.173926,11.037745,9.901564,8.761478,7.6252975,7.676055,7.726812,7.773665,7.824422,7.8751793,7.8361354,7.800996,7.7619514,7.726812,7.687768,7.8517528,8.011833,8.175818,8.335898,8.499884,7.824422,7.1489606,6.473499,5.801942,5.12648,5.774611,6.426646,7.0747766,7.726812,8.374943,8.062591,7.7502384,7.437886,7.125534,6.813182,7.562827,8.312472,9.062118,9.811763,10.561408,10.77615,10.986988,11.20173,11.412568,11.623405,10.475512,9.323712,8.175818,7.0240197,5.8761253,6.5125427,7.1489606,7.7892823,8.4257,9.062118,10.151445,11.23687,12.326198,13.411622,14.50095,13.688834,12.8767185,12.0606985,11.248583,10.436467,10.912805,11.389141,11.861574,12.337912,12.814248,13.150026,13.4858055,13.825488,14.161267,14.50095,12.361338,10.22563,8.086017,5.950309,3.8106966,3.3890212,2.9634414,2.5378613,2.1122816,1.6867018,2.4129205,3.1391394,3.8614538,4.5876727,5.3138914,5.563773,5.813655,6.0635366,6.3134184,6.5633,7.012306,7.461313,7.914223,8.36323,8.812236,11.873287,14.938243,17.999294,21.06425,24.125301,24.012074,23.898846,23.785618,23.676296,23.563068,29.751545,35.93612,42.124596,48.313072,54.501553,51.463924,48.4263,45.388676,42.35105,39.313427,41.413994,43.51066,45.61123,47.711796,49.812363,42.663403,35.514442,28.361578,21.212618,14.063657,12.162213,10.260769,8.36323,6.461786,4.564246,5.298274,6.036206,6.774138,7.5120697,8.250002,8.648251,9.050405,9.448653,9.850807,10.249056,9.538455,8.823949,8.113348,7.3988423,6.688241,5.786324,4.8883114,3.9863946,3.0883822,2.1864653,2.1239948,2.0615244,1.999054,1.9365835,1.8741131,2.9868677,4.0996222,5.212377,6.3251314,7.437886,7.2739015,7.113821,6.949836,6.785851,6.6257706,5.4115014,4.2011366,2.9868677,1.7765031,0.5622339,1.1986516,1.8389735,2.475391,3.1118085,3.7482262,4.2870336,4.825841,5.3607445,5.899552,6.4383593,11.599979,16.761599,21.923218,27.088743,32.250362,40.148968,48.05148,55.950085,63.84869,71.7512,66.58568,61.424057,56.262436,51.100815,45.939198,37.73605,29.536802,21.337559,13.138313,4.939069,6.676528,8.413987,10.151445,11.888905,13.626364,13.911386,14.200311,14.489237,14.774258,15.063184,14.301826,13.536563,12.775204,12.013845,11.248583,10.362284,9.475985,8.58578,7.699481,6.813182,7.812709,8.812236,9.811763,10.81129,11.810817,10.537982,9.261242,7.988407,6.7116675,5.4388323,7.687768,9.936704,12.185639,14.438479,16.687416,18.463919,20.236517,22.01302,23.785618,25.562122,23.961317,22.364416,20.76361,19.162806,17.562002,15.438006,13.314012,11.186112,9.062118,6.9381227,7.461313,7.988407,8.511597,9.0386915,9.561881,8.687295,7.812709,6.9381227,6.0635366,5.1889505,5.1108627,5.036679,4.9624953,4.8883114,4.814128,5.661383,6.5125427,7.363703,8.210958,9.062118,9.589212,10.112402,10.6355915,11.162686,11.685876,10.2881,8.886419,7.4886436,6.086963,4.689187,5.001539,5.3138914,5.6262436,5.938596,6.250948,6.2743745,6.3017054,6.3251314,6.348558,6.375889,15.336493,24.300999,33.261604,42.22611,51.186714,47.08709,42.98747,38.887848,34.788223,30.688602,27.026272,23.363943,19.701614,16.039284,12.373051,11.150972,9.924991,8.699008,7.47693,6.250948,9.86252,13.4740925,17.085665,20.701141,24.312714,25.687063,27.061413,28.435762,29.814016,31.188366,28.51385,25.839334,23.160913,20.486399,17.811884,23.51231,29.212738,34.913166,40.613594,46.31402,38.8488,31.38749,23.926178,16.46096,8.999647,8.960603,8.925464,8.886419,8.85128,8.812236,8.800523,8.78881,8.773191,8.761478,8.749765,7.3988423,6.0518236,4.7009,3.349977,1.999054,2.2137961,2.4246337,2.639376,2.8502135,3.0610514,3.076669,3.0883822,3.1000953,3.1118085,3.1235218,3.6740425,4.224563,4.775084,5.3256044,5.8761253,5.1108627,4.349504,3.5881457,2.8267872,2.0615244,1.6867018,1.3118792,0.93705654,0.5622339,0.18741131,0.27330816,0.3631094,0.44900626,0.5388075,0.62470436,0.80040246,0.97610056,1.1517987,1.3235924,1.4992905,1.8741131,2.2489357,2.6237583,2.998581,3.3734035,3.0610514,2.7486992,2.436347,2.1239948,1.8116426,1.4641509,1.1127546,0.76135844,0.41386664,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,1.175225,2.35045,3.5256753,4.7009,5.8761253,5.4856853,5.099149,4.7126136,4.3260775,3.9356375,3.1508527,2.3621633,1.5734742,0.78868926,0.0,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.26159495,0.3357786,0.41386664,0.48805028,0.5622339,0.58566034,0.61299115,0.63641757,0.6637484,0.6871748,0.6637484,0.63641757,0.61299115,0.58566034,0.5622339,0.4997635,0.43729305,0.37482262,0.31235218,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.57394713,0.6481308,0.7262188,0.80040246,0.8745861,0.81211567,0.74964523,0.6871748,0.62470436,0.5622339,0.5231899,0.48805028,0.44900626,0.41386664,0.37482262,0.38653582,0.39824903,0.41386664,0.42557985,0.43729305,0.37482262,0.31235218,0.24988174,0.18741131,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.28892577,0.38653582,0.48805028,0.58566034,0.6871748,0.80040246,0.9136301,1.0268579,1.1361811,1.2494087,1.3626363,1.475864,1.5890918,1.698415,1.8116426,2.5769055,3.338264,4.0996222,4.860981,5.6262436,5.099149,4.575959,4.0488653,3.5256753,2.998581,5.4895897,7.9766936,10.4637985,12.950902,15.438006,16.050997,16.663988,17.273075,17.886066,18.499058,22.98912,27.475279,31.961437,36.4515,40.937656,39.375896,37.814137,36.24847,34.68671,33.12495,33.987823,34.850693,35.713566,36.57644,37.439312,32.722794,28.010181,23.301472,18.58886,13.8762455,13.911386,13.950429,13.985569,14.024612,14.063657,17.550287,21.036919,24.52355,28.014086,31.500717,31.239122,30.973623,30.712029,30.450434,30.188839,26.975515,23.762192,20.548868,17.33945,14.126127,13.286681,12.4511385,11.611692,10.77615,9.936704,11.0260315,12.111456,13.200784,14.286208,15.375536,0.13665408,0.24597734,0.3513962,0.46071947,0.5661383,0.6754616,0.6832704,0.6910792,0.698888,0.7066968,0.7106012,0.92924774,1.1439898,1.358732,1.5734742,1.7882162,1.8780174,1.9678187,2.05762,2.1474214,2.2372224,2.2489357,2.260649,2.2762666,2.2879796,2.2996929,2.358259,2.4207294,2.4792955,2.541766,2.6003318,2.7682211,2.9400148,3.1118085,3.279698,3.4514916,3.3655949,3.2836022,3.2016098,3.1196175,3.0376248,3.4475873,3.8575494,4.267512,4.677474,5.087436,5.2592297,5.4271193,5.5989127,5.7668023,5.938596,5.6262436,5.3177958,5.009348,4.6969957,4.388548,4.165997,3.9434462,3.7208953,3.4983444,3.2757936,3.6232853,3.9746814,4.3260775,4.6735697,5.024966,5.3841705,5.743376,6.1064854,6.46569,6.824895,6.559396,6.2938967,6.028397,5.7668023,5.5013027,6.8951745,8.289046,9.686822,11.080693,12.4745655,12.252014,12.029464,11.806912,11.584361,11.361811,10.510651,9.663396,8.812236,7.9610763,7.113821,7.0747766,7.0357327,7.000593,6.9615493,6.9264097,7.0513506,7.180196,7.309041,7.433982,7.562827,7.6252975,7.687768,7.7502384,7.812709,7.8751793,7.355894,6.8405128,6.321227,5.805846,5.2865605,5.8487945,6.4110284,6.9732623,7.5394006,8.101635,7.7970915,7.4964523,7.191909,6.89127,6.5867267,7.0357327,7.480835,7.929841,8.378847,8.823949,9.171441,9.518932,9.866425,10.213917,10.561408,9.807858,9.054309,8.296855,7.5433054,6.785851,7.28171,7.7775693,8.273428,8.769287,9.261242,9.839094,10.413041,10.986988,11.560935,12.138786,11.642927,11.147068,10.651209,10.159255,9.663396,10.174872,10.686349,11.20173,11.713207,12.224684,12.521418,12.818152,13.118792,13.415526,13.712261,11.732729,9.753197,7.773665,5.794133,3.8106966,3.3655949,2.9165885,2.4714866,2.0224805,1.5734742,2.241127,2.9087796,3.5764325,4.2440853,4.911738,5.2436123,5.579391,5.911265,6.2431393,6.575013,7.320754,8.066495,8.8083315,9.554072,10.299813,13.169549,16.039284,18.90902,21.778755,24.64849,24.234625,23.820759,23.40689,22.98912,22.575254,28.170261,33.76527,39.36028,44.955288,50.550297,48.102234,45.654175,43.206116,40.758057,38.3139,39.91861,41.52332,43.12803,44.73274,46.337444,39.719482,33.09762,26.475752,19.85779,13.235924,11.666354,10.096785,8.527214,6.957645,5.388075,6.0635366,6.7389984,7.4144597,8.086017,8.761478,9.390087,10.018696,10.6434,11.272009,11.900618,11.029937,10.159255,9.288573,8.421796,7.551114,7.941554,8.335898,8.726339,9.120684,9.511124,9.218294,8.921559,8.628729,8.331994,8.039165,8.128965,8.218767,8.308568,8.398369,8.488171,8.070399,7.6526284,7.2348576,6.817086,6.3993154,5.2279944,4.056674,2.8814487,1.7101282,0.5388075,1.0659018,1.5929961,2.1200905,2.6471848,3.174279,3.9239242,4.6696653,5.4193106,6.165051,6.910792,11.525795,16.140799,20.755802,25.370806,29.98581,35.94002,41.894238,47.844543,53.79876,59.74907,55.85638,51.959785,48.06319,44.1705,40.27391,34.09324,27.908667,21.727999,15.543426,9.362757,11.709302,14.051944,16.398489,18.74113,21.087677,19.924164,18.756748,17.593237,16.42582,15.262308,14.426766,13.591225,12.755682,11.924045,11.088503,10.674636,10.260769,9.850807,9.43694,9.023073,10.323239,11.619501,12.915763,14.215929,15.51219,14.641508,13.770826,12.90405,12.033368,11.162686,12.322293,13.481901,14.641508,15.801116,16.960724,17.975868,18.987108,19.998348,21.013493,22.024733,20.568392,19.115953,17.65961,16.20327,14.750832,13.396004,12.041177,10.686349,9.331521,7.9766936,8.39056,8.8083315,9.226103,9.643873,10.061645,9.007456,7.9532676,6.899079,5.840986,4.786797,4.7087092,4.6267166,4.548629,4.466636,4.388548,5.446641,6.5008297,7.558923,8.617016,9.675109,9.636065,9.600925,9.561881,9.526741,9.487698,9.6243515,9.757101,9.893755,10.0265045,10.163159,9.136301,8.113348,7.08649,6.0635366,5.036679,5.1499066,5.263134,5.376362,5.4856853,5.5989127,12.767395,19.935879,27.10436,34.26894,41.43742,38.274857,35.11229,31.949724,28.787157,25.624592,23.008642,20.396597,17.780647,15.164699,12.548749,11.588266,10.6238785,9.663396,8.699008,7.7385254,10.19049,12.642454,15.0944195,17.546383,19.998348,21.665527,23.328804,24.995983,26.659258,28.326439,25.886187,23.445936,21.005684,18.565434,16.125181,20.310701,24.49622,28.68174,32.863354,37.048874,33.65595,30.259117,26.866192,23.469362,20.076437,18.397543,16.71865,15.043662,13.364769,11.685876,12.494087,13.302299,14.11051,14.918721,15.723028,13.743496,11.760059,9.776623,7.793187,5.813655,5.5832953,5.35684,5.1303844,4.903929,4.6735697,4.853172,5.02887,5.2084727,5.3841705,5.563773,5.5169206,5.473972,5.4271193,5.3841705,5.337318,4.6384296,3.9356375,3.2367494,2.5378613,1.8389735,1.5695697,1.3040704,1.0346665,0.76916724,0.4997635,0.5036679,0.5114767,0.5153811,0.5192855,0.5231899,0.6637484,0.80040246,0.93705654,1.0737107,1.2142692,1.5110037,1.8077383,2.1044729,2.4012074,2.7018464,2.5690966,2.4402514,2.3114061,2.1786566,2.0498111,1.6515622,1.2494087,0.8511597,0.44900626,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,1.3040704,2.6081407,3.9161155,5.2201858,6.524256,6.001066,5.473972,4.950782,4.423688,3.900498,3.1235218,2.3465457,1.5656652,0.78868926,0.011713207,0.11713207,0.22255093,0.3279698,0.43338865,0.5388075,0.43338865,0.3279698,0.22255093,0.11713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.07027924,0.08980125,0.10932326,0.12884527,0.14836729,0.15227169,0.15617609,0.15617609,0.16008049,0.1639849,0.23426414,0.30844778,0.37872702,0.45291066,0.5231899,0.5427119,0.5583295,0.57785153,0.59346914,0.61299115,0.58956474,0.5661383,0.5466163,0.5231899,0.4997635,0.44510186,0.39044023,0.3357786,0.28111696,0.22645533,0.1835069,0.14055848,0.09761006,0.05466163,0.011713207,0.093705654,0.1717937,0.25378615,0.3318742,0.41386664,0.5114767,0.61299115,0.7106012,0.81211567,0.9136301,0.8433509,0.77697605,0.7106012,0.6442264,0.57394713,0.5349031,0.4958591,0.45681506,0.41386664,0.37482262,0.39044023,0.40605783,0.42167544,0.43338865,0.44900626,0.38263142,0.31625658,0.24597734,0.1796025,0.113227665,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.1717937,0.1717937,0.1678893,0.1639849,0.1639849,0.25378615,0.3435874,0.43338865,0.5231899,0.61299115,0.7418364,0.8667773,0.9956226,1.1205635,1.2494087,1.3821584,1.5149081,1.6476578,1.7804074,1.9131571,2.6471848,3.3812122,4.1191444,4.853172,5.5871997,5.056201,4.5291066,3.998108,3.4671092,2.9361105,4.9781127,7.016211,9.058213,11.096312,13.138313,13.856724,14.571229,15.289639,16.008049,16.72646,21.044727,25.359093,29.677362,33.995632,38.3139,37.665768,37.01764,36.369507,35.721375,35.073246,36.47102,37.864895,39.258766,40.65654,42.05041,37.65796,33.269413,28.880863,24.48841,20.099863,20.271656,20.439547,20.61134,20.779228,20.951023,23.719244,26.48356,29.251781,32.020004,34.788223,34.63205,34.475872,34.3236,34.167423,34.01125,31.161034,28.310822,25.460608,22.614298,19.764084,19.119858,18.475632,17.83531,17.191084,16.55076,17.405825,18.264793,19.123762,19.978827,20.837795,0.21083772,0.31625658,0.41777104,0.5192855,0.62079996,0.7262188,0.7418364,0.75354964,0.76916724,0.78478485,0.80040246,0.98000497,1.1596074,1.33921,1.5188124,1.698415,1.815547,1.9365835,2.0537157,2.1708477,2.2879796,2.338737,2.3855898,2.436347,2.4871042,2.5378613,2.5690966,2.6042364,2.6354716,2.6667068,2.7018464,2.8658314,3.0298162,3.193801,3.3616903,3.5256753,3.4475873,3.3694992,3.2914112,3.213323,3.1391394,3.506153,3.8770714,4.2479897,4.618908,4.985922,5.0132523,5.040583,5.0718184,5.099149,5.12648,4.903929,4.6852827,4.466636,4.2440853,4.025439,3.9044023,3.7833657,3.6662338,3.5451972,3.4241607,3.78727,4.1503797,4.513489,4.8765984,5.2358036,5.7316628,6.2275214,6.7233806,7.2192397,7.7111945,7.2192397,6.727285,6.2353306,5.743376,5.251421,6.239235,7.230953,8.218767,9.2104845,10.198298,10.042123,9.885946,9.725866,9.56969,9.413514,8.85128,8.289046,7.726812,7.1606736,6.5984397,6.473499,6.348558,6.223617,6.098676,5.9737353,6.266566,6.559396,6.852226,7.1450562,7.437886,7.3988423,7.363703,7.3246584,7.2856145,7.250475,6.89127,6.5281606,6.168956,5.8097506,5.4505453,5.9268827,6.3993154,6.8756523,7.348085,7.824422,7.531592,7.238762,6.9459314,6.6531014,6.364176,6.5086384,6.6531014,6.7975645,6.942027,7.08649,7.570636,8.050878,8.535024,9.019169,9.499411,9.140205,8.781001,8.421796,8.058686,7.699481,8.050878,8.406178,8.757574,9.108971,9.464272,9.526741,9.589212,9.651682,9.714153,9.776623,9.597021,9.421323,9.24172,9.066022,8.886419,9.43694,9.987461,10.537982,11.088503,11.639023,11.896713,12.154405,12.408191,12.665881,12.923572,11.10412,9.280765,7.4574084,5.6340523,3.8106966,3.3421683,2.87364,2.4012074,1.9326792,1.4641509,2.0732377,2.6823244,3.2914112,3.9044023,4.513489,4.927356,5.3412223,5.758993,6.17286,6.5867267,7.629202,8.667773,9.706344,10.748819,11.787391,14.465811,17.14423,19.818747,22.497166,25.175587,24.457176,23.738766,23.02426,22.305851,21.58744,26.58898,31.590519,36.595963,41.5975,46.59904,44.74445,42.885956,41.02746,39.168964,37.314373,38.42322,39.532074,40.640923,41.753677,42.86253,36.77166,30.680794,24.59383,18.502962,12.412095,11.174399,9.932799,8.691199,7.453504,6.211904,6.824895,7.437886,8.050878,8.663869,9.276859,10.131924,10.983084,11.838148,12.693212,13.548276,12.521418,11.49456,10.467703,9.440845,8.413987,10.096785,11.783486,13.466284,15.152986,16.835783,16.30869,15.781594,15.254499,14.727406,14.200311,13.2671585,12.334006,11.400854,10.471607,9.538455,8.866898,8.191436,7.519879,6.8483214,6.1767645,5.040583,3.9083066,2.77603,1.6437533,0.5114767,0.92924774,1.3470187,1.7647898,2.182561,2.6003318,3.5569105,4.513489,5.473972,6.4305506,7.387129,11.455516,15.523903,19.588387,23.656773,27.72516,31.731077,35.73309,39.739006,43.744923,47.75084,45.123177,42.495514,39.86785,37.24019,34.612526,30.44653,26.284435,22.118439,17.952442,13.786445,16.738173,19.693806,22.645533,25.597261,28.548988,25.93304,23.313187,20.697237,18.081287,15.461433,14.555612,13.645885,12.740065,11.834243,10.924518,10.986988,11.0494585,11.111929,11.174399,11.23687,12.83377,14.426766,16.023666,17.616663,19.213564,18.74894,18.284315,17.815788,17.351164,16.88654,16.95682,17.027098,17.097378,17.167656,17.237936,17.487818,17.7377,17.987581,18.237463,18.487345,17.175465,15.867491,14.555612,13.247637,11.935758,11.354002,10.768341,10.182681,9.597021,9.01136,9.323712,9.63216,9.940608,10.25296,10.561408,9.327617,8.093826,6.8561306,5.6223392,4.388548,4.3026514,4.2167544,4.1308575,4.0488653,3.9629683,5.2279944,6.493021,7.758047,9.023073,10.2881,9.686822,9.089449,8.488171,7.8868923,7.2856145,8.956698,10.627783,12.298867,13.966047,15.637131,13.274967,10.912805,8.550641,6.1884775,3.8263142,4.025439,4.224563,4.423688,4.6267166,4.825841,10.198298,15.570756,20.943214,26.315672,31.68813,29.46262,27.23711,25.0116,22.78609,20.560583,18.994917,17.429253,15.859682,14.294017,12.724447,12.025558,11.326671,10.6238785,9.924991,9.226103,10.518459,11.810817,13.103174,14.395531,15.687888,17.643993,19.596195,21.5523,23.508406,25.460608,23.258524,21.052536,18.84655,16.640562,14.438479,17.10909,19.775797,22.44641,25.11702,27.78763,28.459188,29.130745,29.806208,30.477764,31.14932,27.83058,24.515741,21.197,17.878258,14.56342,16.191557,17.815788,19.443924,21.07206,22.700195,20.084246,17.468296,14.856251,12.240301,9.6243515,8.956698,8.289046,7.621393,6.9537406,6.2860875,6.629675,6.9732623,7.3168497,7.656533,8.00012,7.3597984,6.719476,6.0791545,5.4388323,4.7985106,4.1620927,3.5256753,2.8892577,2.2489357,1.6125181,1.4524376,1.2923572,1.1322767,0.97219616,0.81211567,0.7340276,0.6559396,0.58175594,0.5036679,0.42557985,0.5231899,0.62470436,0.7262188,0.8238289,0.92534333,1.1439898,1.3665408,1.5851873,1.8038338,2.0263848,2.077142,2.1318035,2.182561,2.233318,2.2879796,1.8389735,1.3860629,0.93705654,0.48805028,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,1.43682,2.8697357,4.3065557,5.7394714,7.1762915,6.5125427,5.8487945,5.1889505,4.5252023,3.8614538,3.096191,2.3270237,1.5617609,0.79259366,0.023426414,0.10932326,0.19522011,0.28111696,0.3631094,0.44900626,0.3631094,0.28111696,0.19522011,0.10932326,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.05075723,0.06637484,0.08199245,0.09761006,0.113227665,0.11713207,0.12103647,0.12884527,0.13274968,0.13665408,0.20693332,0.27721256,0.3474918,0.41777104,0.48805028,0.4958591,0.5075723,0.5192855,0.5270943,0.5388075,0.5192855,0.4958591,0.47633708,0.45681506,0.43729305,0.39044023,0.3435874,0.29673457,0.24597734,0.19912452,0.1639849,0.12884527,0.093705654,0.058566034,0.023426414,0.08589685,0.14446288,0.20693332,0.26549935,0.3240654,0.44900626,0.57394713,0.698888,0.8238289,0.94876975,0.8784905,0.80430686,0.7340276,0.659844,0.58566034,0.5466163,0.5036679,0.46071947,0.41777104,0.37482262,0.39434463,0.40996224,0.42557985,0.44510186,0.46071947,0.39044023,0.31625658,0.24597734,0.1717937,0.10151446,0.113227665,0.12494087,0.13665408,0.14836729,0.1639849,0.15617609,0.15227169,0.14836729,0.14055848,0.13665408,0.21864653,0.29673457,0.37872702,0.45681506,0.5388075,0.679366,0.8238289,0.96438736,1.1088502,1.2494087,1.4016805,1.5539521,1.7062237,1.8584955,2.0107672,2.7213683,3.4280653,4.134762,4.841459,5.548156,5.0132523,4.478349,3.9434462,3.408543,2.87364,4.466636,6.0596323,7.6526284,9.245625,10.838621,11.6585455,12.482374,13.306203,14.126127,14.949956,19.096432,23.24681,27.393286,31.53976,35.686237,35.95564,36.221138,36.490543,36.756042,37.025448,38.95422,40.879093,42.807865,44.73664,46.66151,42.593124,38.52864,34.460255,30.391867,26.32348,26.628023,26.928663,27.233206,27.533844,27.838388,29.884295,31.934107,33.98001,36.02592,38.07573,38.028877,37.97812,37.931267,37.884415,37.837563,35.350456,32.863354,30.37625,27.889145,25.398136,24.953035,24.504028,24.058928,23.60992,23.160913,23.789522,24.41813,25.04674,25.671444,26.300053,0.28892577,0.38653582,0.48414588,0.58175594,0.679366,0.77307165,0.79649806,0.8199245,0.8433509,0.8667773,0.8862993,1.0307622,1.1791295,1.3235924,1.4680552,1.6125181,1.756981,1.901444,2.0459068,2.194274,2.338737,2.4246337,2.514435,2.6003318,2.6862288,2.77603,2.7799344,2.7838387,2.7916477,2.795552,2.7994564,2.959537,3.1196175,3.279698,3.4397783,3.5998588,3.5256753,3.455396,3.3812122,3.310933,3.2367494,3.5686235,3.8965936,4.2284675,4.5564375,4.8883114,4.7711797,4.657952,4.5408196,4.4275923,4.3143644,4.181615,4.0527697,3.9239242,3.7911747,3.6623292,3.6467118,3.6271896,3.611572,3.59205,3.5764325,3.951255,4.3260775,4.7009,5.0757227,5.4505453,6.0791545,6.7116675,7.3402762,7.968885,8.601398,7.8790836,7.1606736,6.4383593,5.7199492,5.001539,5.5832953,6.168956,6.754616,7.3402762,7.9259367,7.832231,7.7385254,7.648724,7.5550184,7.461313,7.1880045,6.910792,6.6374836,6.364176,6.086963,5.8761253,5.661383,5.4505453,5.2358036,5.024966,5.481781,5.938596,6.3993154,6.8561306,7.3129454,7.1762915,7.0357327,6.899079,6.7624245,6.6257706,6.422742,6.2197127,6.016684,5.813655,5.610626,6.001066,6.387602,6.774138,7.1606736,7.551114,7.266093,6.984976,6.703859,6.4188375,6.13772,5.9815445,5.8214636,5.6652875,5.5091114,5.349031,5.9659266,6.5867267,7.2036223,7.8205175,8.437413,8.472553,8.507692,8.542832,8.577971,8.6131115,8.823949,9.030883,9.24172,9.452558,9.663396,9.21439,8.761478,8.312472,7.8634663,7.4105554,7.551114,7.6916723,7.832231,7.9727893,8.113348,8.699008,9.288573,9.874233,10.4637985,11.0494585,11.268105,11.486752,11.701493,11.92014,12.138786,10.471607,8.8083315,7.141152,5.477876,3.8106966,3.3187418,2.8267872,2.3348327,1.8428779,1.3509232,1.901444,2.455869,3.0063896,3.5608149,4.1113358,4.6110992,5.1069584,5.606722,6.1025805,6.5984397,7.9337454,9.269051,10.604357,11.939662,13.274967,15.758167,18.245272,20.728472,23.215576,25.698776,24.679728,23.660677,22.641628,21.618675,20.599627,25.0116,29.41967,33.831646,38.239716,42.65169,41.38276,40.11383,38.8488,37.579872,36.31094,36.927837,37.54083,38.157722,38.770714,39.38761,33.82774,28.267872,22.708004,17.148134,11.588266,10.67854,9.768814,8.859089,7.9493628,7.0357327,7.5862536,8.136774,8.687295,9.237816,9.788337,10.869856,11.951375,13.036799,14.118319,15.199838,14.016804,12.829865,11.6468315,10.459893,9.276859,12.252014,15.231073,18.206228,21.185287,24.164345,23.402987,22.641628,21.884174,21.122816,20.361458,18.409256,16.453152,14.4970455,12.54094,10.588739,9.659492,8.734148,7.8049,6.8756523,5.950309,4.8570766,3.7638438,2.6706111,1.5812829,0.48805028,0.79649806,1.1010414,1.4094892,1.717937,2.0263848,3.193801,4.3612175,5.5286336,6.6960497,7.8634663,11.381332,14.903104,18.420969,21.942741,25.460608,27.518227,29.575848,31.633467,33.691086,35.748707,34.389977,33.031242,31.668606,30.309875,28.951143,26.803722,24.6563,22.508879,20.361458,18.214037,21.770947,25.331762,28.892576,32.453392,36.014206,31.941916,27.873528,23.801235,19.73285,15.660558,14.684457,13.704452,12.720543,11.740538,10.764437,11.29934,11.838148,12.376955,12.911859,13.450665,15.344301,17.234032,19.127666,21.021301,22.911032,22.852467,22.7939,22.73143,22.672863,22.614298,21.591345,20.572296,19.553246,18.534197,17.511244,16.999767,16.48829,15.976814,15.461433,14.949956,13.786445,12.619028,11.455516,10.2881,9.124588,9.308095,9.495506,9.679013,9.866425,10.049932,10.25296,10.455989,10.6590185,10.858143,11.061172,9.647778,8.234385,6.817086,5.4036927,3.9863946,3.8965936,3.8067923,3.716991,3.6271896,3.5373883,5.009348,6.481308,7.9532676,9.4291315,10.901091,9.737579,8.574067,7.4105554,6.250948,5.087436,8.292951,11.498465,14.703979,17.909492,21.111103,17.413633,13.712261,10.010887,6.3134184,2.612045,2.900971,3.1859922,3.474918,3.7638438,4.0488653,7.629202,11.205634,14.782067,18.3585,21.938837,20.650383,19.36193,18.073479,16.788929,15.500477,14.981192,14.458001,13.938716,13.419431,12.900145,12.4628525,12.025558,11.588266,11.150972,10.71368,10.84643,10.979179,11.108025,11.240774,11.373524,13.618555,15.863586,18.108618,20.35365,22.59868,20.630861,18.659138,16.69132,14.719597,12.751778,13.903577,15.059279,16.214983,17.370686,18.526388,23.266333,28.006277,32.746223,37.486168,42.22611,37.26752,32.30893,27.354242,22.39565,17.437061,19.88512,22.333181,24.78124,27.229301,29.673458,26.4289,23.180437,19.931974,16.683512,13.438952,12.330102,11.221252,10.116306,9.007456,7.898606,8.406178,8.913751,9.421323,9.928895,10.436467,9.202676,7.968885,6.7311897,5.4973984,4.263607,3.6857557,3.1118085,2.5378613,1.9639144,1.3860629,1.3353056,1.2806439,1.2298868,1.1791295,1.1244678,0.96438736,0.80430686,0.6442264,0.48414588,0.3240654,0.38653582,0.44900626,0.5114767,0.57394713,0.63641757,0.78088045,0.92143893,1.0659018,1.2064602,1.3509232,1.5851873,1.8194515,2.0537157,2.2918842,2.5261483,2.0263848,1.5266213,1.0268579,0.5231899,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,1.5656652,3.1313305,4.6969957,6.2587566,7.824422,7.0240197,6.223617,5.423215,4.6267166,3.8263142,3.06886,2.3114061,1.5539521,0.79649806,0.039044023,0.10151446,0.1678893,0.23426414,0.29673457,0.3631094,0.29673457,0.23426414,0.1678893,0.10151446,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.03513962,0.046852827,0.05466163,0.06637484,0.07418364,0.08199245,0.08980125,0.09761006,0.10541886,0.113227665,0.1796025,0.24597734,0.31625658,0.38263142,0.44900626,0.45291066,0.45681506,0.45681506,0.46071947,0.46071947,0.44510186,0.42557985,0.40996224,0.39434463,0.37482262,0.3357786,0.29673457,0.25378615,0.21474212,0.1756981,0.14836729,0.12103647,0.093705654,0.06637484,0.039044023,0.078088045,0.11713207,0.15617609,0.19912452,0.23816854,0.38653582,0.5388075,0.6871748,0.8355421,0.9878138,0.9097257,0.8316377,0.75354964,0.679366,0.60127795,0.5544251,0.5114767,0.46462387,0.42167544,0.37482262,0.39434463,0.41386664,0.43338865,0.45681506,0.47633708,0.39824903,0.32016098,0.24207294,0.1639849,0.08589685,0.10151446,0.113227665,0.12494087,0.13665408,0.14836729,0.14055848,0.13665408,0.12884527,0.12103647,0.113227665,0.1835069,0.25378615,0.3240654,0.39434463,0.46071947,0.62079996,0.77697605,0.93315214,1.0932326,1.2494087,1.4212024,1.5969005,1.7686942,1.9404879,2.1122816,2.7916477,3.4710135,4.154284,4.83365,5.5130157,4.9742084,4.4314966,3.892689,3.3538816,2.8111696,3.959064,5.1030536,6.2470436,7.3910336,8.538928,9.464272,10.393518,11.318862,12.24811,13.173453,17.152039,21.130625,25.109211,29.083893,33.062477,34.245514,35.428547,36.61158,37.79071,38.973743,41.433517,43.897194,46.356968,48.816742,51.276516,47.52829,43.783966,40.039646,36.295322,32.551003,32.98439,33.421684,33.855072,34.28846,34.725754,36.05325,37.38075,38.708244,40.03574,41.36324,41.421803,41.484276,41.54284,41.601406,41.663876,39.535976,37.411983,35.287987,33.163994,31.036093,30.786211,30.532425,30.278639,30.028757,29.774971,30.173222,30.57147,30.965815,31.364063,31.762312,0.3631094,0.45681506,0.5466163,0.64032197,0.7340276,0.8238289,0.8550641,0.8862993,0.9136301,0.94486535,0.97610056,1.0854238,1.1947471,1.3040704,1.4133936,1.5266213,1.698415,1.8702087,2.0420024,2.2137961,2.3855898,2.514435,2.639376,2.7643168,2.8892577,3.0141985,2.9907722,2.9673457,2.9439192,2.9243972,2.900971,3.0532427,3.2094188,3.3655949,3.521771,3.6740425,3.6076677,3.541293,3.4710135,3.4046388,3.338264,3.6271896,3.9161155,4.2089458,4.4978714,4.786797,4.5291066,4.271416,4.0137253,3.7560349,3.4983444,3.4593005,3.4202564,3.3812122,3.338264,3.2992198,3.3851168,3.4710135,3.5569105,3.638903,3.7247996,4.1113358,4.5017757,4.8883114,5.2748475,5.661383,6.426646,7.191909,7.957172,8.722435,9.487698,8.538928,7.5940623,6.6452928,5.6965227,4.7516575,4.93126,5.1108627,5.290465,5.4700675,5.64967,5.6223392,5.5950084,5.5676775,5.5403466,5.5130157,5.5247293,5.5364423,5.548156,5.563773,5.575486,5.2748475,4.9742084,4.6735697,4.376835,4.0761957,4.6969957,5.3217,5.9425,6.5633,7.1880045,6.949836,6.7116675,6.473499,6.239235,6.001066,5.9542136,5.911265,5.8644123,5.8214636,5.774611,6.0752497,6.375889,6.676528,6.9732623,7.2739015,7.000593,6.7311897,6.4578815,6.184573,5.911265,5.45445,4.9937305,4.533011,4.0722914,3.611572,4.365122,5.1186714,5.8683167,6.621866,7.375416,7.8049,8.234385,8.663869,9.093353,9.526741,9.593117,9.659492,9.725866,9.796145,9.86252,8.898132,7.9376497,6.9732623,6.012779,5.0483923,5.5091114,5.9659266,6.422742,6.8795567,7.336372,7.9610763,8.58578,9.21439,9.839094,10.4637985,10.639496,10.819098,10.994797,11.174399,11.350098,9.8429985,8.335898,6.8287997,5.3217,3.8106966,3.2992198,2.7838387,2.2684577,1.7530766,1.2376955,1.7335546,2.2294137,2.7213683,3.2172275,3.7130866,4.290938,4.872694,5.45445,6.0323014,6.6140575,8.242193,9.874233,11.502369,13.134409,14.762545,17.054428,19.346313,21.638197,23.933987,26.22587,24.902277,23.578686,22.258997,20.935406,19.611813,23.430319,27.248823,31.063425,34.88193,38.700436,38.02107,37.345608,36.66624,35.99078,35.311413,35.43245,35.553486,35.67062,35.791656,35.912693,30.883821,25.851048,20.822178,15.793307,10.764437,10.182681,9.600925,9.023073,8.441318,7.8634663,8.351517,8.835662,9.323712,9.811763,10.299813,11.611692,12.919667,14.231546,15.539521,16.8514,15.5082855,14.165172,12.822057,11.478943,10.135828,14.407245,18.678661,22.946173,27.217588,31.489004,30.493382,29.501663,28.509945,27.518227,26.526508,23.54745,20.568392,17.593237,14.614178,11.639023,10.455989,9.272955,8.089922,6.9068875,5.7238536,4.6735697,3.619381,2.5690966,1.5149081,0.46071947,0.659844,0.8589685,1.0541886,1.2533131,1.4485333,2.8267872,4.2050414,5.5832953,6.9615493,8.335898,11.311053,14.282304,17.253553,20.228708,23.199959,23.309282,23.418604,23.531832,23.641155,23.750479,23.656773,23.563068,23.473267,23.37956,23.285854,23.15701,23.028164,22.899319,22.76657,22.637724,26.803722,30.973623,35.13962,39.30952,43.475517,37.95079,32.429966,26.90914,21.38441,15.863586,14.809398,13.759113,12.704925,11.650736,10.600452,11.611692,12.626837,13.638077,14.649317,15.664462,17.850927,20.041296,22.231667,24.422035,26.612406,26.955994,27.303486,27.647072,27.99066,28.338152,26.22587,24.117493,22.009115,19.896833,17.788456,16.511717,15.238882,13.962143,12.689307,11.412568,10.393518,9.370565,8.351517,7.3324676,6.3134184,7.266093,8.2226715,9.17925,10.131924,11.088503,11.182208,11.275913,11.373524,11.46723,11.560935,9.967939,8.371038,6.7780423,5.181142,3.5881457,3.49444,3.39683,3.3031244,3.2094188,3.1118085,4.7907014,6.473499,8.152391,9.8312845,11.514082,9.788337,8.062591,6.336845,4.6110992,2.8892577,7.629202,12.369146,17.10909,21.849035,26.58898,21.548395,16.511717,11.475039,6.4383593,1.4016805,1.7765031,2.1513257,2.5261483,2.900971,3.2757936,5.056201,6.8405128,8.62092,10.405232,12.185639,11.838148,11.486752,11.139259,10.787864,10.436467,10.963562,11.490656,12.021654,12.548749,13.075843,12.900145,12.724447,12.548749,12.376955,12.201257,11.170495,10.143637,9.116779,8.089922,7.0630636,9.597021,12.130978,14.668839,17.202797,19.736753,18.003199,16.26574,14.532186,12.798631,11.061172,10.701966,10.342762,9.983557,9.620447,9.261242,18.069574,26.877905,35.686237,44.494568,53.298996,46.700554,40.106018,33.50758,26.90914,20.310701,23.578686,26.84667,30.114655,33.38264,36.650623,32.76965,28.888672,25.0116,21.130625,17.24965,15.7035055,14.153459,12.607315,11.061172,9.511124,10.186585,10.858143,11.5297,12.201257,12.8767185,11.045554,9.21439,7.3832245,5.5559645,3.7247996,3.213323,2.7018464,2.1864653,1.6749885,1.1635119,1.2181735,1.2728351,1.3274968,1.3821584,1.43682,1.1947471,0.95267415,0.7106012,0.46852827,0.22645533,0.24988174,0.27330816,0.30063897,0.3240654,0.3513962,0.41386664,0.48024148,0.5466163,0.60908675,0.6754616,1.0932326,1.5110037,1.9287747,2.3465457,2.7643168,2.2137961,1.6632754,1.1127546,0.5622339,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,1.6945106,3.3890212,5.083532,6.7819467,8.476458,7.5394006,6.5984397,5.661383,4.7243266,3.78727,3.0415294,2.2918842,1.5461433,0.79649806,0.05075723,0.093705654,0.14055848,0.1835069,0.23035973,0.27330816,0.23035973,0.1835069,0.14055848,0.093705654,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.015617609,0.023426414,0.027330816,0.031235218,0.039044023,0.046852827,0.058566034,0.06637484,0.078088045,0.08589685,0.15227169,0.21864653,0.28111696,0.3474918,0.41386664,0.40605783,0.40215343,0.39824903,0.39434463,0.38653582,0.3709182,0.359205,0.3435874,0.3279698,0.31235218,0.28111696,0.24597734,0.21474212,0.1835069,0.14836729,0.12884527,0.10932326,0.08980125,0.07027924,0.05075723,0.07027924,0.08980125,0.10932326,0.12884527,0.14836729,0.3240654,0.4997635,0.6754616,0.8511597,1.0268579,0.94096094,0.8589685,0.77697605,0.6949836,0.61299115,0.5661383,0.5192855,0.46852827,0.42167544,0.37482262,0.39824903,0.42167544,0.44119745,0.46462387,0.48805028,0.40605783,0.3240654,0.23816854,0.15617609,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.13665408,0.12884527,0.11713207,0.10932326,0.09761006,0.08589685,0.14836729,0.20693332,0.26940376,0.3279698,0.38653582,0.5583295,0.7340276,0.9058213,1.077615,1.2494087,1.4407244,1.6359446,1.8272603,2.018576,2.2137961,2.8658314,3.5178664,4.169902,4.8219366,5.473972,4.93126,4.3846436,3.8419318,3.2953155,2.7486992,3.4475873,4.1464753,4.841459,5.5403466,6.239235,7.269997,8.300759,9.335425,10.366188,11.400854,15.207646,19.014439,22.821232,26.628023,30.43872,32.535385,34.63205,36.72871,38.82928,40.925945,43.916718,46.911392,49.902164,52.892937,55.887615,52.46345,49.043198,45.619038,42.19878,38.77462,39.340755,39.9108,40.476936,41.04698,41.61312,42.2183,42.82739,43.436474,44.041656,44.650745,44.818634,44.986523,45.15441,45.318398,45.486286,43.7254,41.96061,40.199726,38.43884,36.67405,36.61939,36.56082,36.50226,36.44369,36.38903,36.55692,36.7209,36.888794,37.056683,37.22457,0.43729305,0.5231899,0.61299115,0.698888,0.78868926,0.8745861,0.9136301,0.94876975,0.9878138,1.0268579,1.0619974,1.1361811,1.2142692,1.2884527,1.3626363,1.43682,1.6359446,1.8389735,2.0380979,2.2372224,2.436347,2.6003318,2.7643168,2.9243972,3.0883822,3.2484627,3.2016098,3.1508527,3.1000953,3.049338,2.998581,3.1508527,3.2992198,3.4514916,3.5998588,3.7482262,3.6857557,3.6232853,3.5608149,3.4983444,3.435874,3.6857557,3.9356375,4.1894236,4.4393053,4.689187,4.2870336,3.8887846,3.4866312,3.0883822,2.6862288,2.736986,2.787743,2.8385005,2.8892577,2.9361105,3.1235218,3.310933,3.4983444,3.6857557,3.873167,4.2753205,4.6735697,5.0757227,5.473972,5.8761253,6.774138,7.676055,8.574067,9.475985,10.373997,9.198771,8.023546,6.8483214,5.6730967,4.5017757,4.2753205,4.0488653,3.8263142,3.5998588,3.3734035,3.4124475,3.4514916,3.4866312,3.5256753,3.5608149,3.8614538,4.1620927,4.462732,4.7633705,5.0640097,4.6735697,4.2870336,3.900498,3.513962,3.1235218,3.912211,4.7009,5.4856853,6.2743745,7.0630636,6.7233806,6.387602,6.0518236,5.7121406,5.376362,5.4856853,5.5989127,5.7121406,5.825368,5.938596,6.1494336,6.364176,6.575013,6.785851,7.000593,6.7389984,6.473499,6.211904,5.950309,5.688714,4.9234514,4.1620927,3.4007344,2.639376,1.8741131,2.7643168,3.6506162,4.5369153,5.423215,6.3134184,7.137247,7.9610763,8.78881,9.612638,10.436467,10.362284,10.2881,10.213917,10.135828,10.061645,8.58578,7.113821,5.6379566,4.1620927,2.6862288,3.4632049,4.2362766,5.0132523,5.786324,6.5633,7.223144,7.8868923,8.550641,9.21439,9.874233,10.010887,10.151445,10.2881,10.424754,10.561408,9.21439,7.8634663,6.5125427,5.1616197,3.8106966,3.2757936,2.736986,2.1981785,1.6632754,1.1244678,1.5617609,1.999054,2.436347,2.87364,3.310933,3.9746814,4.6384296,5.298274,5.9620223,6.6257706,8.550641,10.475512,12.400381,14.325252,16.250122,18.35069,20.45126,22.551826,24.64849,26.74906,25.124828,23.500597,21.876366,20.24823,18.623999,21.849035,25.074072,28.299107,31.524143,34.74918,34.663284,34.573483,34.487587,34.401688,34.311886,33.937065,33.56224,33.18742,32.812595,32.437775,27.935999,23.438128,18.936352,14.438479,9.936704,9.686822,9.43694,9.187058,8.937177,8.687295,9.112875,9.538455,9.964035,10.38571,10.81129,12.349625,13.887959,15.426293,16.960724,18.499058,16.999767,15.500477,14.001186,12.501896,10.998701,16.562475,22.126247,27.686117,33.24989,38.813663,37.58768,36.3617,35.135715,33.91364,32.687656,28.685644,24.687536,20.685524,16.687416,12.689307,11.248583,9.811763,8.374943,6.9381227,5.5013027,4.4861584,3.474918,2.463678,1.4485333,0.43729305,0.5231899,0.61299115,0.698888,0.78868926,0.8745861,2.463678,4.0488653,5.6379566,7.223144,8.812236,11.23687,13.661504,16.086138,18.51077,20.93931,19.100336,17.261362,15.426293,13.58732,11.748346,12.923572,14.098797,15.274021,16.449247,17.624472,19.514202,21.400028,23.285854,25.175587,27.061413,31.836496,36.61158,41.386665,46.161747,50.936832,43.96357,36.986404,30.01314,23.035973,16.062712,14.938243,13.813775,12.689307,11.560935,10.436467,11.924045,13.411622,14.899199,16.386776,17.874353,20.361458,22.848562,25.335667,27.826675,30.31378,31.063425,31.81307,32.562714,33.31236,34.062004,30.860395,27.66269,24.46108,21.263374,18.061766,16.023666,13.989473,11.951375,9.913278,7.8751793,7.000593,6.126007,5.251421,4.376835,3.4983444,5.22409,6.949836,8.675582,10.401327,12.123169,12.111456,12.099743,12.08803,12.076316,12.0606985,10.2881,8.511597,6.7389984,4.9624953,3.1859922,3.0883822,2.9868677,2.8892577,2.787743,2.6862288,4.575959,6.461786,8.351517,10.237343,12.123169,9.839094,7.551114,5.263134,2.9751544,0.6871748,6.9615493,13.235924,19.514202,25.788576,32.06295,25.687063,19.311174,12.939189,6.5633,0.18741131,0.6481308,1.1127546,1.5734742,2.0380979,2.4988174,2.4871042,2.475391,2.463678,2.4480603,2.436347,3.0259118,3.611572,4.2011366,4.786797,5.376362,6.949836,8.52331,10.100689,11.674163,13.251541,13.337439,13.423335,13.513136,13.599033,13.688834,11.498465,9.311999,7.125534,4.939069,2.7486992,5.575486,8.398369,11.225157,14.051944,16.874826,15.375536,13.8762455,12.373051,10.87376,9.37447,7.5003567,5.6262436,3.7482262,1.8741131,0.0,12.8767185,25.749533,38.62625,51.499065,64.375786,56.137497,47.899208,39.66092,31.426535,23.188246,27.276154,31.364063,35.451973,39.535976,43.623886,39.110397,34.60081,30.087324,25.573835,21.06425,19.073006,17.085665,15.098324,13.110983,11.123642,11.963089,12.798631,13.638077,14.473619,15.313066,12.888432,10.4637985,8.039165,5.610626,3.1859922,2.736986,2.2879796,1.8389735,1.3860629,0.93705654,1.1010414,1.261122,1.4251068,1.5890918,1.7491722,1.4251068,1.1010414,0.77307165,0.44900626,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.60127795,1.1986516,1.7999294,2.4012074,2.998581,2.4012074,1.7999294,1.1986516,0.60127795,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.8233559,3.6506162,5.473972,7.3012323,9.124588,8.050878,6.9732623,5.899552,4.825841,3.7482262,3.0141985,2.2762666,1.5383345,0.80040246,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.37482262,0.3631094,0.3513962,0.3357786,0.3240654,0.31235218,0.30063897,0.28892577,0.27330816,0.26159495,0.24988174,0.22645533,0.19912452,0.1756981,0.14836729,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.26159495,0.46071947,0.6637484,0.8628729,1.0619974,0.97610056,0.8862993,0.80040246,0.7106012,0.62470436,0.57394713,0.5231899,0.47633708,0.42557985,0.37482262,0.39824903,0.42557985,0.44900626,0.47633708,0.4997635,0.41386664,0.3240654,0.23816854,0.14836729,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.113227665,0.1639849,0.21083772,0.26159495,0.31235218,0.4997635,0.6871748,0.8745861,1.0619974,1.2494087,1.4641509,1.6749885,1.8858263,2.1005683,2.3114061,2.9361105,3.5608149,4.1894236,4.814128,5.4388323,4.8883114,4.337791,3.78727,3.2367494,2.6862288,2.9361105,3.1859922,3.435874,3.6857557,3.9356375,5.0757227,6.211904,7.348085,8.488171,9.6243515,13.263254,16.902157,20.537155,24.17606,27.811058,30.825256,33.839455,36.849747,39.86395,42.87424,46.399918,49.92559,53.451267,56.973038,60.498714,57.398617,54.298523,51.198425,48.09833,44.998238,45.701027,46.399918,47.098804,47.801598,48.500484,48.387257,48.27403,48.1608,48.05148,47.93825,48.21156,48.488773,48.76208,49.03929,49.3126,47.91092,46.513145,45.111465,43.713688,42.312008,42.44866,42.58922,42.725872,42.86253,42.999184,42.93671,42.87424,42.81177,42.749302,42.68683,0.48805028,0.5661383,0.6481308,0.7262188,0.80821127,0.8862993,0.92924774,0.97219616,1.0151446,1.0580931,1.1010414,1.2064602,1.3118792,1.4133936,1.5188124,1.6242313,1.7843118,1.9443923,2.1044729,2.2645533,2.4246337,2.5612879,2.6940374,2.8306916,2.9634414,3.1000953,3.0415294,2.9868677,2.9283018,2.8697357,2.8111696,3.135235,3.4593005,3.7794614,4.1035266,4.423688,4.263607,4.1035266,3.9434462,3.7833657,3.6232853,3.7989833,3.970777,4.142571,4.3143644,4.4861584,4.0996222,3.7130866,3.3265507,2.9361105,2.5495746,2.612045,2.6745155,2.736986,2.7994564,2.8619268,3.0415294,3.2172275,3.39683,3.5725281,3.7482262,4.185519,4.618908,5.056201,5.4895897,5.9268827,6.6648145,7.406651,8.144583,8.886419,9.6243515,8.495979,7.363703,6.2353306,5.1030536,3.9746814,3.7794614,3.5842414,3.3890212,3.193801,2.998581,3.0922866,3.1859922,3.2757936,3.3694992,3.4632049,3.6662338,3.873167,4.0761957,4.283129,4.4861584,4.4861584,4.4861584,4.4861584,4.4861584,4.4861584,5.0483923,5.610626,6.1767645,6.7389984,7.3012323,6.89127,6.481308,6.0713453,5.661383,5.251421,5.349031,5.4505453,5.548156,5.64967,5.7511845,5.930787,6.114294,6.297801,6.481308,6.66091,6.348558,6.0323014,5.716045,5.4036927,5.087436,4.5291066,3.9668727,3.408543,2.8463092,2.2879796,2.951728,3.611572,4.2753205,4.939069,5.5989127,6.4110284,7.2192397,8.031356,8.839567,9.651682,9.522837,9.393991,9.269051,9.140205,9.01136,7.9259367,6.8366084,5.7511845,4.661856,3.5764325,3.9863946,4.4002614,4.814128,5.22409,5.6379566,6.2040954,6.7663293,7.3324676,7.898606,8.460839,8.749765,9.0386915,9.323712,9.612638,9.901564,8.796618,7.6916723,6.5867267,5.481781,4.376835,3.873167,3.3694992,2.8658314,2.366068,1.8623998,2.25284,2.6432803,3.0337205,3.4241607,3.8106966,4.4041657,4.9937305,5.5832953,6.17286,6.7624245,8.683391,10.604357,12.521418,14.442384,16.36335,18.623999,20.880743,23.141392,25.40204,27.66269,26.284435,24.906181,23.531832,22.153578,20.775324,23.44984,26.124355,28.79887,31.473387,34.151806,33.91364,33.679375,33.44511,33.210846,32.97658,32.746223,32.51586,32.285503,32.05514,31.824783,27.631454,23.442032,19.248703,15.055375,10.862047,10.651209,10.436467,10.22563,10.010887,9.80005,10.174872,10.549695,10.924518,11.29934,11.674163,12.810344,13.946525,15.078801,16.214983,17.351164,17.323833,17.300406,17.273075,17.24965,17.226223,20.775324,24.324427,27.873528,31.426535,34.975636,33.636425,32.30112,30.96191,29.626604,28.287394,24.804668,21.321941,17.839214,14.356487,10.87376,9.608734,8.343708,7.0786815,5.813655,4.548629,3.7599394,2.97125,2.1786566,1.3899672,0.60127795,0.76916724,0.93315214,1.1010414,1.2689307,1.43682,3.6740425,5.9073606,8.140678,10.377901,12.611219,13.790349,14.965574,16.144703,17.323833,18.499058,17.671324,16.843592,16.015858,15.188125,14.364296,14.96167,15.559043,16.156416,16.75379,17.351164,19.330696,21.310228,23.289759,25.26929,27.248823,31.258644,35.26456,39.274384,43.2803,47.286217,41.433517,35.576912,29.724215,23.86761,18.011007,16.773312,15.531713,14.294017,13.052417,11.810817,13.384291,14.957765,16.531239,18.10081,19.674282,20.67381,21.669432,22.668959,23.664581,24.664108,25.546503,26.4289,27.311295,28.19369,29.076084,26.366428,23.656773,20.943214,18.233559,15.523903,13.774731,12.025558,10.276386,8.52331,6.774138,6.1455293,5.5169206,4.884407,4.2557983,3.6232853,4.93126,6.2353306,7.5394006,8.843472,10.151445,10.377901,10.604357,10.8308115,11.061172,11.287627,9.901564,8.519405,7.1333427,5.74728,4.3612175,4.40807,4.4510183,4.4978714,4.5408196,4.5876727,5.7238536,6.8561306,7.9923115,9.128492,10.260769,8.488171,6.719476,4.9468775,3.174279,1.4016805,6.3993154,11.393045,16.394585,21.388315,26.38595,21.927124,17.468296,13.005564,8.546737,4.087909,4.814128,5.5364423,6.262661,6.98888,7.7111945,7.4300776,7.1489606,6.8639393,6.5828223,6.3017054,6.606249,6.914696,7.223144,7.531592,7.8361354,9.183154,10.526268,11.873287,13.216402,14.56342,14.743023,14.922626,15.102228,15.281831,15.461433,12.950902,10.444276,7.9337454,5.423215,2.912684,5.4505453,7.988407,10.526268,13.06413,15.598087,14.422862,13.243732,12.068507,10.889378,9.714153,8.183627,6.657006,5.1303844,3.6037633,2.0732377,12.076316,22.079395,32.082474,42.085552,52.08863,45.56047,39.03231,32.50415,25.975988,19.451733,22.911032,26.370333,29.829634,33.288933,36.748234,33.148376,29.544611,25.94085,22.34099,18.737226,17.440966,16.148607,14.852346,13.556085,12.263727,12.2793455,12.291059,12.306676,12.322293,12.337912,10.545791,8.75367,6.9615493,5.169429,3.3734035,2.8502135,2.3231194,1.7999294,1.2767396,0.74964523,0.8784905,1.0112402,1.1400855,1.2689307,1.4016805,2.084951,2.7682211,3.455396,4.138666,4.825841,3.8692627,2.9165885,1.9600099,1.0034313,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.48024148,0.96048295,1.4407244,1.9209659,2.4012074,1.9209659,1.4407244,0.96048295,0.48024148,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.4602464,2.920493,4.380739,5.840986,7.3012323,6.813182,6.3251314,5.8370814,5.349031,4.860981,3.9278288,2.9907722,2.05762,1.1205635,0.18741131,0.1796025,0.1717937,0.1639849,0.15617609,0.14836729,0.12884527,0.10932326,0.08980125,0.07027924,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.10932326,0.1639849,0.22255093,0.28111696,0.3357786,0.3631094,0.39434463,0.42167544,0.44900626,0.47633708,0.45681506,0.44119745,0.42167544,0.40605783,0.38653582,0.3357786,0.28111696,0.23035973,0.1756981,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.06637484,0.06637484,0.07027924,0.07418364,0.07418364,0.26549935,0.45681506,0.6442264,0.8355421,1.0268579,0.92924774,0.8355421,0.7418364,0.6442264,0.5505207,0.5114767,0.47633708,0.43729305,0.39824903,0.3631094,0.39824903,0.43729305,0.47633708,0.5114767,0.5505207,0.45291066,0.3553006,0.25769055,0.16008049,0.062470436,0.07418364,0.08199245,0.093705654,0.10151446,0.113227665,0.10932326,0.10151446,0.09761006,0.093705654,0.08589685,0.12103647,0.15617609,0.19131571,0.22645533,0.26159495,0.42948425,0.59737355,0.76526284,0.93315214,1.1010414,1.358732,1.620327,1.8819219,2.1396124,2.4012074,2.9048753,3.408543,3.9161155,4.4197836,4.9234514,4.579864,4.2362766,3.8887846,3.5451972,3.2016098,3.3890212,3.5764325,3.7638438,3.951255,4.138666,5.0913405,6.044015,6.996689,7.9493628,8.898132,11.818625,14.735214,17.651802,20.568392,23.488884,26.28834,29.087797,31.887253,34.68671,37.486168,40.871284,44.2564,47.641518,51.026634,54.41175,52.71724,51.022728,49.328217,47.63371,45.939198,46.485813,47.036335,47.586853,48.137375,48.687897,48.1569,47.6259,47.098804,46.567806,46.036808,45.564373,45.09194,44.61951,44.147076,43.674644,42.378384,41.078217,39.781956,38.485695,37.18943,37.290947,37.396366,37.501785,37.6072,37.71262,37.759476,37.806328,37.85318,37.90394,37.95079,0.5388075,0.60908675,0.6832704,0.75354964,0.8277333,0.9019169,0.94876975,0.9956226,1.0424755,1.0893283,1.1361811,1.2728351,1.4055848,1.542239,1.678893,1.8116426,1.9326792,2.0537157,2.1708477,2.2918842,2.4129205,2.5183394,2.6276627,2.7330816,2.8424048,2.951728,2.8853533,2.8189783,2.7565079,2.690133,2.6237583,3.1196175,3.6154766,4.1113358,4.60329,5.099149,4.841459,4.5837684,4.3260775,4.068387,3.8106966,3.9083066,4.0020123,4.095718,4.193328,4.2870336,3.912211,3.5373883,3.1625657,2.787743,2.4129205,2.4871042,2.5612879,2.639376,2.7135596,2.787743,2.9556324,3.1235218,3.2914112,3.4593005,3.6232853,4.095718,4.564246,5.036679,5.505207,5.9737353,6.5554914,7.1333427,7.715099,8.296855,8.874706,7.7892823,6.703859,5.618435,4.5369153,3.4514916,3.2836022,3.1196175,2.9556324,2.7916477,2.6237583,2.7721257,2.920493,3.06886,3.213323,3.3616903,3.4710135,3.5842414,3.6935644,3.802888,3.912211,4.298747,4.689187,5.0757227,5.462259,5.8487945,6.1884775,6.524256,6.8639393,7.1997175,7.5394006,7.055255,6.571109,6.0908675,5.606722,5.12648,5.212377,5.298274,5.388075,5.473972,5.563773,5.716045,5.8683167,6.0205884,6.17286,6.3251314,5.958118,5.591104,5.22409,4.853172,4.4861584,4.1308575,3.7716527,3.416352,3.057147,2.7018464,3.1391394,3.5764325,4.0137253,4.4510183,4.8883114,5.6809053,6.477403,7.2739015,8.066495,8.862993,8.683391,8.503788,8.324185,8.140678,7.9610763,7.262188,6.5633,5.8644123,5.1616197,4.462732,4.513489,4.564246,4.6110992,4.661856,4.7126136,5.181142,5.645766,6.114294,6.5828223,7.0513506,7.4886436,7.9259367,8.36323,8.800523,9.237816,8.378847,7.5159745,6.657006,5.7980375,4.939069,4.4705405,4.0020123,3.533484,3.06886,2.6003318,2.9439192,3.2836022,3.6271896,3.970777,4.3143644,4.829746,5.349031,5.8644123,6.3836975,6.899079,8.81614,10.729298,12.6463585,14.559516,16.476578,18.893402,21.314133,23.734861,26.15559,28.57632,27.444044,26.315672,25.183395,24.055023,22.926651,25.050644,27.17464,29.298634,31.426535,33.55053,33.167896,32.785267,32.402634,32.020004,31.637371,31.551476,31.465578,31.383585,31.297688,31.211792,27.326912,23.442032,19.557152,15.672271,11.787391,11.611692,11.435994,11.2642,11.088503,10.912805,11.23687,11.560935,11.888905,12.212971,12.537036,13.271063,14.001186,14.735214,15.469242,16.199366,17.651802,19.100336,20.548868,22.001307,23.44984,24.988174,26.526508,28.06094,29.599274,31.137608,29.689075,28.236637,26.788103,25.335667,23.887133,20.92369,17.956347,14.992905,12.025558,9.062118,7.968885,6.8756523,5.786324,4.6930914,3.5998588,3.0337205,2.463678,1.8975395,1.3314011,0.76135844,1.0112402,1.2572175,1.5031948,1.7530766,1.999054,4.884407,7.7658563,10.647305,13.528754,16.414106,16.343828,16.273548,16.20327,16.13299,16.062712,16.246218,16.42582,16.609327,16.792833,16.976341,16.995863,17.015385,17.034906,17.054428,17.073952,19.147188,21.220427,23.293663,25.366901,27.436235,30.67689,33.91754,37.158195,40.39885,43.6356,38.903465,34.167423,29.431385,24.69925,19.96321,18.608381,17.253553,15.8987255,14.543899,13.189071,14.844538,16.503908,18.159374,19.818747,21.474213,20.982258,20.490303,19.998348,19.506393,19.010534,20.025679,21.040823,22.05597,23.071114,24.086258,21.868557,19.646952,17.429253,15.207646,12.986042,11.525795,10.061645,8.601398,7.137247,5.6730967,5.290465,4.903929,4.521298,4.134762,3.7482262,4.6345253,5.520825,6.4032197,7.289519,8.175818,8.644346,9.108971,9.577498,10.046027,10.510651,9.518932,8.52331,7.5276875,6.532065,5.5364423,5.727758,5.919074,6.1064854,6.297801,6.4891167,6.871748,7.2543793,7.633106,8.015738,8.398369,7.141152,5.883934,4.6267166,3.3694992,2.1122816,5.833177,9.554072,13.271063,16.991959,20.712854,18.167183,15.621513,13.075843,10.534078,7.988407,8.976221,9.964035,10.951848,11.935758,12.923572,12.373051,11.818625,11.268105,10.71368,10.163159,10.19049,10.217821,10.2451515,10.272482,10.299813,11.416472,12.529227,13.645885,14.75864,15.875299,16.148607,16.421915,16.69132,16.964628,17.237936,14.40334,11.572648,8.738052,5.9073606,3.076669,5.3256044,7.57454,9.823476,12.076316,14.325252,13.470188,12.615124,11.760059,10.904996,10.049932,8.870802,7.6916723,6.5086384,5.3295093,4.1503797,11.279819,18.409256,25.538694,32.668133,39.801476,34.983444,30.165411,25.34738,20.529346,15.711315,18.54591,21.376602,24.211199,27.04189,29.876486,27.18245,24.48841,21.798277,19.10424,16.414106,15.808925,15.207646,14.606369,14.001186,13.399908,12.591698,11.783486,10.979179,10.170968,9.362757,8.203149,7.043542,5.883934,4.7243266,3.5608149,2.9634414,2.3621633,1.7608855,1.1635119,0.5622339,0.659844,0.75745404,0.8550641,0.95267415,1.0502841,2.7447948,4.4393053,6.133816,7.8283267,9.526741,7.629202,5.7316628,3.8341231,1.9365835,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.359205,0.71841,1.0815194,1.4407244,1.7999294,1.4407244,1.0815194,0.71841,0.359205,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0932326,2.1903696,3.2836022,4.380739,5.473972,5.575486,5.6730967,5.774611,5.8761253,5.9737353,4.841459,3.7091823,2.5769055,1.4446288,0.31235218,0.27330816,0.23426414,0.19131571,0.15227169,0.113227665,0.09761006,0.08199245,0.06637484,0.05075723,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.08980125,0.14055848,0.19522011,0.24597734,0.30063897,0.3670138,0.43338865,0.5036679,0.5700427,0.63641757,0.61689556,0.59346914,0.5700427,0.5466163,0.5231899,0.44510186,0.3631094,0.28502136,0.20693332,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.06637484,0.07418364,0.078088045,0.08199245,0.08589685,0.26940376,0.44900626,0.62860876,0.80821127,0.9878138,0.8862993,0.78088045,0.679366,0.57785153,0.47633708,0.44900626,0.42557985,0.39824903,0.37482262,0.3513962,0.39824903,0.44900626,0.4997635,0.5505207,0.60127795,0.49195468,0.38653582,0.27721256,0.1717937,0.062470436,0.07027924,0.078088045,0.08589685,0.093705654,0.10151446,0.10151446,0.10541886,0.10932326,0.10932326,0.113227665,0.13274968,0.15227169,0.1717937,0.19131571,0.21083772,0.359205,0.5075723,0.6559396,0.80430686,0.94876975,1.2572175,1.5656652,1.8741131,2.1786566,2.4871042,2.87364,3.2562714,3.6428072,4.029343,4.4119744,4.271416,4.1308575,3.9942036,3.853645,3.7130866,3.8380275,3.9629683,4.087909,4.21285,4.337791,5.1069584,5.872221,6.6413884,7.406651,8.175818,10.373997,12.572175,14.766449,16.964628,19.162806,21.751425,24.33614,26.924759,29.513376,32.09809,35.346554,38.59111,41.83567,45.080227,48.324787,48.035862,47.74303,47.454105,47.16518,46.876255,47.2745,47.676655,48.074905,48.473152,48.87531,47.926537,46.981674,46.0329,45.084133,44.139267,42.91719,41.699017,40.476936,39.258766,38.036686,36.841938,35.647194,34.452446,33.257698,32.06295,32.133232,32.207413,32.281597,32.351875,32.42606,32.582237,32.738415,32.898495,33.05467,33.210846,0.58566034,0.6520352,0.71841,0.78088045,0.8472553,0.9136301,0.96438736,1.0190489,1.0698062,1.1205635,1.175225,1.33921,1.5031948,1.6710842,1.8350691,1.999054,2.0810463,2.1591344,2.241127,2.3192148,2.4012074,2.4792955,2.5612879,2.639376,2.7213683,2.7994564,2.7291772,2.6549935,2.5808098,2.5105307,2.436347,3.1039999,3.7716527,4.4393053,5.1069584,5.774611,5.4193106,5.0640097,4.7087092,4.3534083,3.998108,4.01763,4.0332475,4.0527697,4.068387,4.087909,3.7247996,3.3616903,2.998581,2.639376,2.2762666,2.3621633,2.4480603,2.5378613,2.6237583,2.7135596,2.8697357,3.0259118,3.1859922,3.3421683,3.4983444,4.0059166,4.5095844,5.0132523,5.520825,6.0244927,6.446168,6.8639393,7.2856145,7.703386,8.125061,7.08649,6.044015,5.0054436,3.9668727,2.9243972,2.7916477,2.6549935,2.5183394,2.3855898,2.2489357,2.4519646,2.6549935,2.8580225,3.0610514,3.2640803,3.2757936,3.2914112,3.3070288,3.3226464,3.338264,4.1113358,4.8883114,5.661383,6.4383593,7.211431,7.3246584,7.437886,7.551114,7.6643414,7.773665,7.2192397,6.6648145,6.1103897,5.5559645,5.001539,5.0757227,5.1499066,5.22409,5.298274,5.376362,5.4973984,5.618435,5.743376,5.8644123,5.989353,5.5676775,5.1460023,4.728231,4.3065557,3.8887846,3.7326086,3.5764325,3.4241607,3.2679846,3.1118085,3.3265507,3.5373883,3.7482262,3.9629683,4.173806,4.9546866,5.735567,6.5164475,7.2934237,8.074304,7.843944,7.60968,7.37932,7.1450562,6.910792,6.5984397,6.2860875,5.9737353,5.661383,5.349031,5.036679,4.7243266,4.4119744,4.0996222,3.78727,4.1581883,4.5291066,4.8961205,5.267039,5.6379566,6.223617,6.813182,7.3988423,7.988407,8.574067,7.9610763,7.3441806,6.7311897,6.114294,5.5013027,5.067914,4.6345253,4.2011366,3.7716527,3.338264,3.631094,3.9278288,4.220659,4.5173936,4.814128,5.2592297,5.704332,6.1494336,6.590631,7.0357327,8.94889,10.858143,12.767395,14.676648,16.585901,19.16671,21.74752,24.328331,26.90914,29.486046,28.603651,27.721256,26.838861,25.956467,25.074072,26.65145,28.224924,29.798397,31.375776,32.94925,32.41825,31.891157,31.360159,30.82916,30.29816,30.360632,30.419197,30.481668,30.540234,30.5988,27.022367,23.445936,19.865599,16.289165,12.712734,12.576079,12.439425,12.298867,12.162213,12.025558,12.298867,12.576079,12.849388,13.1266,13.399908,13.731783,14.059752,14.391626,14.719597,15.051471,17.975868,20.900265,23.824663,26.74906,29.673458,29.201025,28.724688,28.24835,27.775917,27.29958,25.73782,24.17606,22.610394,21.048632,19.486872,17.03881,14.590752,12.146595,9.698535,7.250475,6.329036,5.4115014,4.4900627,3.5686235,2.6510892,2.3035975,1.9600099,1.6164225,1.2689307,0.92534333,1.2533131,1.5812829,1.9092526,2.233318,2.5612879,6.0908675,9.6243515,13.153932,16.683512,20.21309,18.893402,17.57762,16.261835,14.942147,13.626364,14.817206,16.008049,17.202797,18.393639,19.588387,19.030056,18.471727,17.913397,17.358973,16.800642,18.963682,21.130625,23.293663,25.460608,27.623646,30.099037,32.570522,35.04201,37.513496,39.988888,36.373413,32.757935,29.142458,25.526981,21.911505,20.44345,18.97149,17.503435,16.031475,14.56342,16.304783,18.046146,19.791414,21.532778,23.274141,21.290705,19.311174,17.327738,15.344301,13.360865,14.508759,15.656653,16.804546,17.952442,19.100336,17.370686,15.641035,13.911386,12.181735,10.44818,9.272955,8.101635,6.9264097,5.7511845,4.575959,4.435401,4.2948427,4.154284,4.0137253,3.873167,4.3416953,4.806319,5.270943,5.735567,6.2001905,6.9068875,7.6135845,8.324185,9.030883,9.737579,9.132397,8.527214,7.9220324,7.3168497,6.7116675,7.0474463,7.3832245,7.719003,8.050878,8.386656,8.015738,7.648724,7.277806,6.9068875,6.5359693,5.794133,5.0522966,4.31046,3.5686235,2.8267872,5.267039,7.7111945,10.151445,12.595602,15.035853,14.407245,13.778636,13.146122,12.517513,11.888905,13.138313,14.387722,15.637131,16.88654,18.135948,17.316025,16.492195,15.668366,14.848442,14.024612,13.770826,13.520945,13.2671585,13.013372,12.763491,13.645885,14.532186,15.418485,16.300879,17.18718,17.554192,17.917301,18.284315,18.647425,19.014439,15.855778,12.70102,9.546264,6.3915067,3.2367494,5.2006636,7.1606736,9.124588,11.088503,13.048512,12.517513,11.986515,11.4516115,10.920613,10.38571,9.554072,8.722435,7.890797,7.0591593,6.223617,10.48332,14.739119,18.998821,23.25462,27.510418,24.406418,21.298513,18.19061,15.0827055,11.974802,14.180789,16.382872,18.58886,20.794846,23.000834,21.216522,19.436115,17.651802,15.871395,14.087084,14.176885,14.2666855,14.356487,14.446288,14.53609,12.907954,11.275913,9.647778,8.015738,6.387602,5.860508,5.3334136,4.806319,4.279225,3.7482262,3.076669,2.4012074,1.7257458,1.0502841,0.37482262,0.44119745,0.5036679,0.5700427,0.63641757,0.698888,3.4046388,6.1103897,8.81614,11.521891,14.223738,11.385237,8.546737,5.704332,2.8658314,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.23816854,0.48024148,0.71841,0.96048295,1.1986516,0.96048295,0.71841,0.48024148,0.23816854,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7301232,1.4602464,2.1903696,2.920493,3.6506162,4.337791,5.024966,5.7121406,6.3993154,7.08649,5.758993,4.4275923,3.096191,1.7686942,0.43729305,0.3631094,0.29283017,0.21864653,0.14836729,0.07418364,0.06637484,0.05466163,0.046852827,0.03513962,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.07418364,0.12103647,0.1678893,0.21474212,0.26159495,0.3709182,0.47633708,0.58566034,0.6910792,0.80040246,0.77307165,0.74574083,0.71841,0.6910792,0.6637484,0.5544251,0.44900626,0.339683,0.23426414,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.07027924,0.078088045,0.08589685,0.093705654,0.10151446,0.26940376,0.44119745,0.60908675,0.78088045,0.94876975,0.8394465,0.7301232,0.62079996,0.5114767,0.39824903,0.38653582,0.37482262,0.3631094,0.3513962,0.3357786,0.39824903,0.46071947,0.5231899,0.58566034,0.6481308,0.5309987,0.41386664,0.29673457,0.1796025,0.062470436,0.06637484,0.07418364,0.078088045,0.08199245,0.08589685,0.09761006,0.10932326,0.11713207,0.12884527,0.13665408,0.14055848,0.14836729,0.15227169,0.15617609,0.1639849,0.28892577,0.41777104,0.5466163,0.6715572,0.80040246,1.1557031,1.5110037,1.8663043,2.2216048,2.5769055,2.8385005,3.1039999,3.3694992,3.6349986,3.900498,3.9668727,4.029343,4.095718,4.1581883,4.224563,4.2870336,4.349504,4.4119744,4.474445,4.5369153,5.1186714,5.704332,6.2860875,6.8678436,7.4495993,8.929368,10.405232,11.881096,13.360865,14.836729,17.210606,19.588387,21.962263,24.33614,26.71392,29.81792,32.92192,36.02592,39.133823,42.237823,43.35058,44.467236,45.583897,46.69665,47.81331,48.06319,48.313072,48.562954,48.812836,49.062717,47.69618,46.33354,44.967,43.604362,42.237823,40.270004,38.302185,36.334366,34.36655,32.39873,31.305498,30.21617,29.122936,28.029703,26.936472,26.975515,27.018463,27.057508,27.096552,27.135595,27.404999,27.670498,27.939903,28.205402,28.474806,0.63641757,0.6949836,0.75354964,0.80821127,0.8667773,0.92534333,0.98390937,1.038571,1.097137,1.1557031,1.2142692,1.4055848,1.6008049,1.796025,1.9912452,2.1864653,2.2294137,2.2684577,2.3075018,2.3465457,2.3855898,2.4402514,2.4910088,2.5456703,2.5964274,2.6510892,2.5690966,2.4910088,2.4090161,2.330928,2.2489357,3.0883822,3.9317331,4.7711797,5.610626,6.4500723,5.997162,5.5442514,5.0913405,4.6384296,4.1894236,4.126953,4.068387,4.0059166,3.9473507,3.8887846,3.5373883,3.1859922,2.8385005,2.4871042,2.135708,2.2372224,2.338737,2.436347,2.5378613,2.639376,2.7838387,2.9322062,3.0805733,3.2289407,3.3734035,3.9161155,4.454923,4.9937305,5.5364423,6.0752497,6.336845,6.5945354,6.8561306,7.113821,7.375416,6.379793,5.3841705,4.388548,3.39683,2.4012074,2.2957885,2.1903696,2.084951,1.979532,1.8741131,2.1318035,2.3894942,2.6471848,2.9048753,3.1625657,3.0805733,3.0024853,2.9243972,2.8424048,2.7643168,3.9239242,5.087436,6.250948,7.4144597,8.574067,8.460839,8.351517,8.238289,8.125061,8.011833,7.3832245,6.75852,6.1299114,5.5013027,4.8765984,4.939069,5.001539,5.0640097,5.12648,5.1889505,5.278752,5.3724575,5.466163,5.5559645,5.64967,5.1772375,4.704805,4.2323723,3.7599394,3.2875066,3.3343596,3.3812122,3.4280653,3.4788225,3.5256753,3.513962,3.4983444,3.4866312,3.474918,3.4632049,4.2284675,4.9937305,5.758993,6.524256,7.2856145,7.000593,6.715572,6.4305506,6.1455293,5.8644123,5.938596,6.012779,6.086963,6.1611466,6.239235,5.563773,4.8883114,4.21285,3.5373883,2.8619268,3.135235,3.408543,3.6818514,3.951255,4.224563,4.9624953,5.700427,6.4383593,7.1762915,7.914223,7.5433054,7.172387,6.801469,6.4305506,6.0635366,5.6652875,5.267039,4.8687897,4.474445,4.0761957,4.322173,4.5681505,4.8180323,5.0640097,5.3138914,5.6848097,6.055728,6.4305506,6.801469,7.1762915,9.081639,10.983084,12.888432,14.79378,16.69913,19.44002,22.18091,24.921799,27.658785,30.399675,29.763258,29.130745,28.494328,27.861814,27.225397,28.24835,29.275208,30.29816,31.32502,32.351875,31.672512,30.993145,30.317684,29.638317,28.962856,29.165884,29.372818,29.575848,29.78278,29.98581,26.717825,23.445936,20.177952,16.906061,13.638077,13.536563,13.438952,13.337439,13.235924,13.138313,13.360865,13.58732,13.813775,14.036326,14.262781,14.188598,14.118319,14.044135,13.973856,13.899672,18.299932,22.700195,27.100456,31.500717,35.900978,33.413876,30.926771,28.435762,25.948658,23.461554,21.786564,20.111576,18.436588,16.761599,15.086611,13.157836,11.229061,9.296382,7.367607,5.4388323,4.689187,3.9434462,3.193801,2.4480603,1.698415,1.5773785,1.456342,1.3314011,1.2103647,1.0893283,1.4953861,1.901444,2.3114061,2.717464,3.1235218,7.3012323,11.478943,15.656653,19.834364,24.012074,21.446882,18.88169,16.316498,13.751305,11.186112,13.388195,15.594183,17.796265,19.998348,22.200432,21.06425,19.931974,18.795792,17.65961,16.52343,18.784079,21.040823,23.297567,25.554314,27.811058,29.51728,31.223505,32.925823,34.63205,36.338272,33.843357,31.348446,28.853533,26.35862,23.863707,22.278519,20.693333,19.108145,17.522957,15.93777,17.76503,19.59229,21.41955,23.24681,25.074072,21.603058,18.12814,14.657126,11.186112,7.7111945,8.991838,10.272482,11.553126,12.83377,14.11051,12.872814,11.631214,10.393518,9.151918,7.914223,7.0240197,6.13772,5.251421,4.3612175,3.474918,3.5803368,3.6857557,3.7911747,3.8965936,3.998108,4.044961,4.0918136,4.134762,4.181615,4.224563,5.173333,6.1181984,7.066968,8.015738,8.960603,8.745861,8.531119,8.316377,8.101635,7.8868923,8.367134,8.847376,9.327617,9.807858,10.2881,9.163632,8.043069,6.918601,5.7980375,4.6735697,4.447114,4.220659,3.9942036,3.7638438,3.5373883,4.7009,5.8683167,7.0318284,8.1992445,9.362757,10.647305,11.931853,13.216402,14.50095,15.789403,17.300406,18.81141,20.326319,21.837322,23.348326,22.258997,21.165764,20.072533,18.9793,17.886066,17.355068,16.82407,16.289165,15.758167,15.223265,15.879204,16.535143,17.191084,17.843119,18.499058,18.955873,19.416592,19.873407,20.330223,20.787037,17.308216,13.833297,10.354475,6.8756523,3.4007344,5.0757227,6.7507114,8.4257,10.100689,11.775677,11.564839,11.354002,11.143164,10.936231,10.725393,10.241247,9.753197,9.269051,8.784905,8.300759,9.686822,11.06898,12.455043,13.841106,15.223265,13.825488,12.431617,11.033841,9.636065,8.238289,9.815667,11.393045,12.970425,14.547803,16.125181,15.250595,14.379913,13.509232,12.634645,11.763964,12.544845,13.325725,14.11051,14.89139,15.676175,13.224211,10.768341,8.316377,5.8644123,3.4124475,3.5178664,3.6232853,3.7287042,3.8341231,3.9356375,3.1859922,2.436347,1.6867018,0.93705654,0.18741131,0.21864653,0.25378615,0.28502136,0.31625658,0.3513962,4.0644827,7.7814736,11.49456,15.211552,18.924637,15.141272,11.361811,7.578445,3.795079,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.12103647,0.23816854,0.359205,0.48024148,0.60127795,0.48024148,0.359205,0.23816854,0.12103647,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3631094,0.7301232,1.0932326,1.4602464,1.8233559,3.1000953,4.376835,5.64967,6.9264097,8.1992445,6.6726236,5.1460023,3.619381,2.0888553,0.5622339,0.45681506,0.3513962,0.24597734,0.14055848,0.039044023,0.031235218,0.027330816,0.023426414,0.015617609,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.05466163,0.09761006,0.14055848,0.1835069,0.22645533,0.3709182,0.5192855,0.6676528,0.8160201,0.96438736,0.92924774,0.8980125,0.8667773,0.8316377,0.80040246,0.6637484,0.5309987,0.39434463,0.26159495,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.07418364,0.08199245,0.093705654,0.10151446,0.113227665,0.27330816,0.43338865,0.59346914,0.75354964,0.9136301,0.79649806,0.679366,0.5583295,0.44119745,0.3240654,0.3240654,0.3240654,0.3240654,0.3240654,0.3240654,0.39824903,0.47633708,0.5505207,0.62470436,0.698888,0.57394713,0.44510186,0.31625658,0.19131571,0.062470436,0.06637484,0.06637484,0.07027924,0.07418364,0.07418364,0.093705654,0.10932326,0.12884527,0.14446288,0.1639849,0.15227169,0.14055848,0.13274968,0.12103647,0.113227665,0.21864653,0.3279698,0.43338865,0.5427119,0.6481308,1.0541886,1.456342,1.8584955,2.260649,2.6628022,2.8072653,2.951728,3.096191,3.240654,3.3890212,3.6584249,3.9278288,4.1972322,4.466636,4.73604,4.73604,4.73604,4.73604,4.73604,4.73604,5.134289,5.532538,5.930787,6.329036,6.7233806,7.480835,8.238289,8.995743,9.753197,10.510651,12.67369,14.836729,16.999767,19.162806,21.325846,24.289286,27.256632,30.220074,33.183514,36.15086,38.6692,41.191444,43.70978,46.228123,48.750366,48.851883,48.94949,49.051006,49.148617,49.25013,47.465816,45.68541,43.9011,42.120693,40.33638,37.62282,34.905357,32.191795,29.478237,26.760773,25.772959,24.78124,23.793427,22.801708,21.813896,21.821705,21.82561,21.833418,21.841227,21.849035,22.227762,22.60649,22.981312,23.360039,23.738766,0.6871748,0.737932,0.78868926,0.8394465,0.8862993,0.93705654,0.999527,1.0619974,1.1244678,1.1869383,1.2494087,1.475864,1.698415,1.9248703,2.1513257,2.3738766,2.3738766,2.3738766,2.3738766,2.3738766,2.3738766,2.4012074,2.4246337,2.4480603,2.475391,2.4988174,2.4129205,2.3231194,2.2372224,2.1513257,2.0615244,3.076669,4.087909,5.099149,6.114294,7.125534,6.575013,6.0244927,5.473972,4.9234514,4.376835,4.2362766,4.0996222,3.9629683,3.8263142,3.6857557,3.349977,3.0141985,2.6745155,2.338737,1.999054,2.1122816,2.2255092,2.338737,2.4480603,2.5612879,2.7018464,2.8385005,2.9751544,3.1118085,3.2484627,3.8263142,4.4002614,4.9742084,5.548156,6.126007,6.223617,6.3251314,6.426646,6.524256,6.6257706,5.6730967,4.7243266,3.775557,2.8267872,1.8741131,1.7999294,1.7257458,1.6515622,1.5734742,1.4992905,1.8116426,2.1239948,2.436347,2.7486992,3.0610514,2.8892577,2.7135596,2.5378613,2.3621633,2.1864653,3.736513,5.2865605,6.8366084,8.386656,9.936704,9.600925,9.261242,8.925464,8.58578,8.250002,7.551114,6.8483214,6.1494336,5.4505453,4.7516575,4.7985106,4.8492675,4.900025,4.950782,5.001539,5.0640097,5.12648,5.1889505,5.251421,5.3138914,4.786797,4.263607,3.736513,3.213323,2.6862288,2.9361105,3.1859922,3.435874,3.6857557,3.9356375,3.7013733,3.4632049,3.2250361,2.9868677,2.7486992,3.4983444,4.251894,5.001539,5.7511845,6.5008297,6.1611466,5.825368,5.4856853,5.1499066,4.814128,5.2748475,5.735567,6.2001905,6.66091,7.125534,6.086963,5.0483923,4.0137253,2.9751544,1.9365835,2.1122816,2.2879796,2.463678,2.639376,2.8111696,3.7013733,4.5876727,5.473972,6.364176,7.250475,7.125534,7.000593,6.8756523,6.7507114,6.6257706,6.262661,5.899552,5.5364423,5.173333,4.814128,5.0132523,5.212377,5.4115014,5.610626,5.813655,6.114294,6.4110284,6.7116675,7.012306,7.3129454,9.21439,11.111929,13.013372,14.9109125,16.812357,19.713327,22.614298,25.511364,28.412334,31.313307,30.926771,30.53633,30.149794,29.763258,29.376722,29.849155,30.325493,30.80183,31.274261,31.750599,30.926771,30.099037,29.275208,28.45138,27.623646,27.975042,28.326439,28.673931,29.025326,29.376722,26.41328,23.44984,20.486399,17.526861,14.56342,14.50095,14.438479,14.376009,14.313539,14.251068,14.426766,14.59856,14.774258,14.949956,15.125654,14.649317,14.176885,13.700547,13.224211,12.751778,18.623999,24.500124,30.37625,36.24847,42.124596,37.626724,33.12495,28.623173,24.125301,19.623526,17.839214,16.050997,14.262781,12.4745655,10.686349,9.276859,7.8634663,6.4500723,5.036679,3.6232853,3.049338,2.475391,1.901444,1.3235924,0.74964523,0.8511597,0.94876975,1.0502841,1.1517987,1.2494087,1.737459,2.2255092,2.7135596,3.2016098,3.6857557,8.511597,13.337439,18.163279,22.98912,27.811058,24.00036,20.18576,16.375063,12.564366,8.749765,11.963089,15.176412,18.38583,21.599154,24.812477,23.098444,21.388315,19.674282,17.964155,16.250122,18.600573,20.951023,23.301472,25.651922,27.998468,28.93943,29.876486,30.813543,31.750599,32.687656,31.313307,29.938957,28.560703,27.186354,25.812004,24.113588,22.411268,20.712854,19.010534,17.31212,19.225277,21.138433,23.05159,24.960844,26.874,21.911505,16.94901,11.986515,7.0240197,2.0615244,3.474918,4.8883114,6.3017054,7.7111945,9.124588,8.374943,7.6252975,6.8756523,6.126007,5.376362,4.775084,4.173806,3.5764325,2.9751544,2.3738766,2.7252727,3.076669,3.4241607,3.775557,4.123049,3.7482262,3.3734035,2.998581,2.6237583,2.2489357,3.435874,4.6267166,5.813655,7.000593,8.187531,8.36323,8.538928,8.710721,8.886419,9.062118,9.686822,10.311526,10.936231,11.560935,12.185639,10.311526,8.437413,6.5633,4.689187,2.8111696,3.1000953,3.3890212,3.6740425,3.9629683,4.251894,4.138666,4.025439,3.912211,3.7989833,3.6857557,6.8873653,10.088976,13.286681,16.48829,19.685997,21.4625,23.239002,25.0116,26.788103,28.560703,27.198067,25.839334,24.476698,23.114061,21.751425,20.93931,20.12329,19.311174,18.499058,17.686943,18.112522,18.538101,18.963682,19.389261,19.810938,20.361458,20.911978,21.4625,22.01302,22.563541,18.760653,14.96167,11.162686,7.363703,3.5608149,4.950782,6.336845,7.726812,9.112875,10.498938,10.612165,10.725393,10.838621,10.951848,11.061172,10.924518,10.787864,10.651209,10.510651,10.373997,8.886419,7.3988423,5.911265,4.423688,2.9361105,3.2484627,3.5608149,3.873167,4.1894236,4.5017757,5.4505453,6.3993154,7.348085,8.300759,9.249529,9.288573,9.323712,9.362757,9.4018,9.43694,10.912805,12.388668,13.860628,15.336493,16.812357,13.536563,10.260769,6.98888,3.7130866,0.43729305,1.175225,1.9131571,2.6510892,3.3890212,4.123049,3.2992198,2.475391,1.6515622,0.8238289,0.0,0.0,0.0,0.0,0.0,0.0,4.7243266,9.448653,14.176885,18.90121,23.625538,18.90121,14.176885,9.448653,4.7243266,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.8623998,3.7247996,5.5871997,7.4495993,9.311999,7.5862536,5.8644123,4.138666,2.4129205,0.6871748,0.5505207,0.41386664,0.27330816,0.13665408,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.37482262,0.5622339,0.74964523,0.93705654,1.1244678,1.0893283,1.0502841,1.0112402,0.97610056,0.93705654,0.77307165,0.61299115,0.44900626,0.28892577,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.27330816,0.42557985,0.57394713,0.7262188,0.8745861,0.74964523,0.62470436,0.4997635,0.37482262,0.24988174,0.26159495,0.27330816,0.28892577,0.30063897,0.31235218,0.39824903,0.48805028,0.57394713,0.6637484,0.74964523,0.61299115,0.47633708,0.3357786,0.19912452,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.14836729,0.23816854,0.3240654,0.41386664,0.4997635,0.94876975,1.4016805,1.8506867,2.2996929,2.7486992,2.77603,2.7994564,2.8267872,2.8502135,2.87364,3.349977,3.8263142,4.298747,4.775084,5.251421,5.1889505,5.12648,5.0640097,5.001539,4.939069,5.1499066,5.3607445,5.575486,5.786324,6.001066,6.036206,6.0752497,6.114294,6.1494336,6.1884775,8.136774,10.088976,12.037272,13.985569,15.93777,18.764557,21.58744,24.414227,27.23711,30.063898,33.987823,37.911747,41.83567,45.7635,49.687424,49.636665,49.585907,49.539055,49.4883,49.437542,47.23546,45.03728,42.8391,40.63702,38.43884,34.975636,31.51243,28.049225,24.586021,21.12672,20.236517,19.350218,18.463919,17.573715,16.687416,16.663988,16.636658,16.613232,16.585901,16.562475,17.050524,17.538574,18.026625,18.51077,18.998821,0.58566034,0.6442264,0.7027924,0.76135844,0.8160201,0.8745861,0.92924774,0.98000497,1.0307622,1.0854238,1.1361811,1.3157835,1.4992905,1.678893,1.8584955,2.0380979,2.0654287,2.0927596,2.1200905,2.1474214,2.174752,2.1786566,2.1864653,2.1903696,2.194274,2.1981785,2.1239948,2.0459068,1.9678187,1.8897307,1.8116426,3.1781836,4.5408196,5.9073606,7.2739015,8.636538,7.9064145,7.172387,6.4383593,5.708236,4.9742084,4.728231,4.478349,4.2323723,3.9863946,3.736513,3.408543,3.076669,2.7486992,2.416825,2.0888553,2.1591344,2.233318,2.3035975,2.377781,2.4480603,2.639376,2.8306916,3.018103,3.2094188,3.4007344,4.0605783,4.7204223,5.380266,6.04011,6.699954,6.649197,6.5945354,6.5437784,6.4891167,6.4383593,5.520825,4.60329,3.6857557,2.7682211,1.8506867,1.7647898,1.678893,1.5969005,1.5110037,1.4251068,1.6593709,1.8897307,2.1239948,2.3543546,2.5886188,2.6432803,2.697942,2.7526035,2.8072653,2.8619268,4.1035266,5.3412223,6.5828223,7.824422,9.062118,8.706817,8.351517,7.996216,7.6409154,7.2856145,6.7819467,6.278279,5.7707067,5.267039,4.7633705,4.786797,4.806319,4.829746,4.853172,4.8765984,4.83365,4.7907014,4.747753,4.704805,4.661856,4.251894,3.8380275,3.4241607,3.0141985,2.6003318,2.7994564,2.998581,3.2016098,3.4007344,3.5998588,3.3694992,3.1391394,2.9087796,2.67842,2.4480603,3.0220075,3.5959544,4.165997,4.7399445,5.3138914,5.181142,5.0522966,4.9234514,4.7907014,4.661856,5.0718184,5.477876,5.883934,6.2938967,6.699954,6.262661,5.825368,5.388075,4.950782,4.513489,4.3729305,4.2323723,4.0918136,3.951255,3.8106966,4.318269,4.825841,5.3334136,5.840986,6.348558,6.5828223,6.813182,7.0474463,7.28171,7.5120697,7.988407,8.468649,8.944985,9.421323,9.901564,10.61607,11.330575,12.045081,12.759586,13.4740925,12.915763,12.353529,11.795199,11.23687,10.674636,12.041177,13.411622,14.778163,16.144703,17.511244,20.127193,22.743143,25.359093,27.971138,30.587088,30.930676,31.274261,31.613945,31.957533,32.30112,31.707651,31.114182,30.520712,29.931149,29.337679,28.716879,28.092175,27.471375,26.84667,26.22587,26.596788,26.971611,27.34253,27.713448,28.08827,25.210726,22.337086,19.463446,16.585901,13.712261,13.6810255,13.653695,13.622459,13.591225,13.563893,13.353056,13.142218,12.93138,12.724447,12.513609,12.166118,11.818625,11.471134,11.123642,10.77615,15.383345,19.994444,24.605543,29.216642,33.823837,30.278639,26.729538,23.184341,19.635239,16.086138,16.066616,16.043188,16.019762,15.996336,15.976814,13.376482,10.780055,8.183627,5.5832953,2.9868677,2.5964274,2.2059872,1.815547,1.4290112,1.038571,1.2181735,1.4016805,1.5851873,1.7686942,1.9482968,3.049338,4.1464753,5.2436123,6.3407493,7.437886,10.58093,13.727879,16.870922,20.01787,23.160913,20.138906,17.1169,14.0948925,11.072885,8.050878,11.377428,14.703979,18.034433,21.360985,24.687536,23.613825,22.544018,21.470308,20.396597,19.326792,20.693333,22.063778,23.434223,24.804668,26.175114,26.65145,27.131691,27.608028,28.084366,28.560703,27.444044,26.327385,25.210726,24.094067,22.973503,21.48983,20.006157,18.51858,17.034906,15.551234,17.01148,18.475632,19.935879,21.400028,22.86418,18.94416,15.024139,11.10412,7.1841,3.2640803,4.0761957,4.8883114,5.700427,6.5125427,7.3246584,7.0201154,6.715572,6.4110284,6.1064854,5.801942,5.2318993,4.6657605,4.095718,3.5295796,2.9634414,3.240654,3.521771,3.802888,4.084005,4.3612175,3.912211,3.4632049,3.0141985,2.5612879,2.1122816,3.2289407,4.3416953,5.4583545,6.571109,7.687768,7.621393,7.558923,7.492548,7.426173,7.363703,8.699008,10.034314,11.365715,12.70102,14.036326,11.732729,9.4291315,7.1216297,4.8180323,2.514435,2.7486992,2.9829633,3.2172275,3.4514916,3.6857557,3.6076677,3.5256753,3.4475873,3.3655949,3.2875066,5.899552,8.507692,11.115833,13.727879,16.33602,17.725986,19.11205,20.502016,21.888079,23.274141,22.364416,21.45469,20.544964,19.635239,18.725513,17.811884,16.894348,15.980719,15.063184,14.149553,16.808453,19.471254,22.130152,24.78905,27.447948,25.815908,24.183868,22.551826,20.919786,19.287746,16.585901,13.884054,11.178304,8.476458,5.774611,6.4891167,7.1997175,7.914223,8.624825,9.339331,9.24172,9.148014,9.054309,8.956698,8.862993,8.75367,8.648251,8.538928,8.433509,8.324185,7.1294384,5.9346914,4.7399445,3.5451972,2.35045,2.8619268,3.3734035,3.8887846,4.4002614,4.911738,5.4115014,5.9073606,6.4032197,6.902983,7.3988423,7.4300776,7.461313,7.4886436,7.519879,7.551114,8.730244,9.909373,11.088503,12.271536,13.450665,10.865952,8.281238,5.6965227,3.1118085,0.5231899,1.3353056,2.1435168,2.9556324,3.7638438,4.575959,3.6584249,2.7447948,1.8311646,0.9136301,0.0,0.0,0.0,0.0,0.0,0.0,3.7833657,7.570636,11.354002,15.141272,18.924637,15.18422,11.443803,7.703386,3.9668727,0.22645533,0.19912452,0.1717937,0.14055848,0.113227665,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.5031948,3.0102942,4.513489,6.0205884,7.523783,6.1455293,4.7633705,3.3851168,2.0068626,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.07027924,0.12884527,0.1835069,0.24207294,0.30063897,0.42557985,0.5505207,0.6754616,0.80040246,0.92534333,0.92924774,0.93315214,0.94096094,0.94486535,0.94876975,0.8316377,0.7145056,0.59737355,0.48024148,0.3631094,0.30454338,0.24597734,0.19131571,0.13274968,0.07418364,0.078088045,0.08589685,0.08980125,0.093705654,0.10151446,0.24597734,0.39434463,0.5427119,0.6910792,0.8394465,0.7301232,0.62079996,0.5153811,0.40605783,0.30063897,0.30454338,0.30844778,0.31625658,0.32016098,0.3240654,0.40605783,0.48805028,0.57394713,0.6559396,0.737932,0.60908675,0.48414588,0.3553006,0.22645533,0.10151446,0.093705654,0.08980125,0.08589685,0.078088045,0.07418364,0.10541886,0.13665408,0.1639849,0.19522011,0.22645533,0.19131571,0.16008049,0.12884527,0.093705654,0.062470436,0.12884527,0.19912452,0.26549935,0.3318742,0.39824903,0.77697605,1.1557031,1.53443,1.9092526,2.2879796,2.3894942,2.4910088,2.5964274,2.697942,2.7994564,3.232845,3.6662338,4.095718,4.5291066,4.9624953,5.1772375,5.3919797,5.606722,5.8214636,6.036206,6.0713453,6.1025805,6.133816,6.168956,6.2001905,6.168956,6.133816,6.1025805,6.0713453,6.036206,7.6838636,9.327617,10.971371,12.619028,14.262781,16.683512,19.10424,21.521065,23.941795,26.362524,29.833538,33.308456,36.77947,40.250484,43.7254,44.41648,45.111465,45.802544,46.49362,47.188606,45.127083,43.065556,41.00794,38.94641,36.888794,33.874596,30.860395,27.850101,24.835903,21.82561,21.044727,20.263847,19.486872,18.705992,17.92511,17.893875,17.858736,17.827501,17.796265,17.761126,18.296028,18.827028,19.36193,19.89293,20.423927,0.48805028,0.5544251,0.61689556,0.6832704,0.74574083,0.81211567,0.8550641,0.8980125,0.94096094,0.98390937,1.0268579,1.1596074,1.2962615,1.4290112,1.5656652,1.698415,1.7530766,1.8116426,1.8663043,1.9209659,1.9756275,1.9600099,1.9443923,1.9287747,1.9131571,1.901444,1.8311646,1.7647898,1.698415,1.6281357,1.5617609,3.279698,4.997635,6.715572,8.433509,10.151445,9.2339115,8.320281,7.406651,6.4891167,5.575486,5.2162814,4.860981,4.5017757,4.1464753,3.78727,3.4632049,3.1430438,2.8189783,2.4988174,2.174752,2.2059872,2.241127,2.2723622,2.3035975,2.338737,2.5808098,2.822883,3.0649557,3.3070288,3.5491016,4.2948427,5.040583,5.786324,6.5281606,7.2739015,7.0708723,6.8639393,6.66091,6.453977,6.250948,5.364649,4.478349,3.5959544,2.7096553,1.8233559,1.7296503,1.6359446,1.5383345,1.4446288,1.3509232,1.5031948,1.6554666,1.8077383,1.9600099,2.1122816,2.397303,2.6823244,2.9673457,3.252367,3.5373883,4.466636,5.395884,6.329036,7.2582836,8.187531,7.816613,7.4417906,7.0708723,6.6960497,6.3251314,6.016684,5.704332,5.395884,5.083532,4.775084,4.7711797,4.7633705,4.759466,4.755562,4.7516575,4.60329,4.454923,4.3065557,4.1581883,4.0137253,3.7130866,3.4124475,3.1118085,2.8111696,2.514435,2.6628022,2.8111696,2.9634414,3.1118085,3.2640803,3.0415294,2.8189783,2.5964274,2.3738766,2.1513257,2.5456703,2.9400148,3.3343596,3.7287042,4.123049,4.2011366,4.279225,4.357313,4.435401,4.513489,4.8648853,5.2162814,5.571582,5.9229784,6.2743745,6.4383593,6.5984397,6.7624245,6.9264097,7.08649,6.6335793,6.1767645,5.7238536,5.267039,4.814128,4.939069,5.067914,5.196759,5.3217,5.4505453,6.04011,6.629675,7.2192397,7.8088045,8.398369,9.718058,11.033841,12.353529,13.6693125,14.989,16.218887,17.448774,18.678661,19.908546,21.138433,19.717232,18.296028,16.87873,15.457528,14.036326,14.871868,15.70741,16.542952,17.378494,18.214037,20.54106,22.871988,25.202917,27.533844,29.860868,30.93458,32.00829,33.078094,34.151806,35.225517,33.566147,31.906775,30.2435,28.58413,26.924759,26.503082,26.085312,25.663635,25.245865,24.82419,25.218534,25.616783,26.011127,26.405472,26.799816,24.012074,21.22433,18.436588,15.648844,12.861101,12.8650055,12.86891,12.86891,12.872814,12.8767185,12.2793455,11.685876,11.088503,10.495033,9.901564,9.679013,9.460366,9.24172,9.019169,8.800523,12.146595,15.488764,18.834837,22.18091,25.523077,22.930555,20.334127,17.741604,15.145176,12.548749,14.294017,16.03538,17.776743,19.518106,21.263374,17.48001,13.696643,9.913278,6.133816,2.35045,2.1435168,1.9404879,1.7335546,1.5305257,1.3235924,1.5890918,1.8545911,2.1200905,2.3855898,2.6510892,4.357313,6.0635366,7.773665,9.479889,11.186112,12.654168,14.118319,15.582469,17.04662,18.51077,16.281357,14.048039,11.814721,9.581403,7.348085,10.791768,14.235451,17.679134,21.118912,24.562595,24.129206,23.695818,23.266333,22.832945,22.399555,22.789995,23.180437,23.570877,23.961317,24.351757,24.367374,24.386896,24.402514,24.41813,24.437654,23.578686,22.715813,21.856844,20.997875,20.138906,18.866072,17.597141,16.32821,15.059279,13.786445,14.801589,15.812829,16.82407,17.839214,18.850454,15.97291,13.095366,10.217821,7.3402762,4.462732,4.6735697,4.8883114,5.099149,5.3138914,5.5247293,5.6652875,5.805846,5.9464045,6.083059,6.223617,5.688714,5.153811,4.618908,4.084005,3.5491016,3.7599394,3.970777,4.181615,4.388548,4.5993857,4.0761957,3.5491016,3.0259118,2.4988174,1.9756275,3.018103,4.0605783,5.1030536,6.1455293,7.1880045,6.883461,6.578918,6.2743745,5.9659266,5.661383,7.70729,9.753197,11.799104,13.841106,15.8870125,13.153932,10.416945,7.6838636,4.9468775,2.2137961,2.3933985,2.5769055,2.7604125,2.9439192,3.1235218,3.076669,3.0298162,2.9829633,2.9361105,2.8892577,4.9078336,6.9264097,8.94889,10.967466,12.986042,13.989473,14.989,15.988527,16.988054,17.987581,17.530766,17.073952,16.613232,16.156416,15.699601,14.6805525,13.665408,12.6463585,11.631214,10.612165,15.5082855,20.400501,25.296621,30.192743,35.088863,31.270357,27.455757,23.641155,19.826555,16.011953,14.407245,12.802535,11.197825,9.593117,7.988407,8.023546,8.062591,8.101635,8.136774,8.175818,7.871275,7.570636,7.266093,6.9654536,6.66091,6.5867267,6.5086384,6.4305506,6.3524623,6.2743745,5.3724575,4.4705405,3.5686235,2.6667068,1.7608855,2.475391,3.1859922,3.900498,4.6110992,5.3256044,5.368553,5.4154058,5.4583545,5.505207,5.548156,5.571582,5.5950084,5.618435,5.6418614,5.661383,6.547683,7.433982,8.316377,9.202676,10.088976,8.191436,6.297801,4.4041657,2.5066261,0.61299115,1.4953861,2.377781,3.260176,4.142571,5.024966,4.0215344,3.0141985,2.0107672,1.0034313,0.0,0.0,0.0,0.0,0.0,0.0,2.8463092,5.688714,8.535024,11.381332,14.223738,11.471134,8.714626,5.958118,3.2055142,0.44900626,0.39434463,0.339683,0.28502136,0.23035973,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1478943,2.2957885,3.4436827,4.591577,5.735567,4.7009,3.6662338,2.631567,1.5969005,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.10151446,0.1796025,0.25769055,0.3357786,0.41386664,0.47633708,0.5388075,0.60127795,0.6637484,0.7262188,0.77307165,0.8199245,0.8667773,0.9136301,0.96438736,0.8902037,0.8160201,0.74574083,0.6715572,0.60127795,0.4958591,0.39434463,0.29283017,0.19131571,0.08589685,0.08589685,0.08199245,0.078088045,0.078088045,0.07418364,0.21864653,0.3631094,0.5114767,0.6559396,0.80040246,0.7106012,0.62079996,0.5309987,0.44119745,0.3513962,0.3474918,0.3435874,0.3435874,0.339683,0.3357786,0.41386664,0.49195468,0.5700427,0.6481308,0.7262188,0.60908675,0.49195468,0.3709182,0.25378615,0.13665408,0.12884527,0.11713207,0.10932326,0.09761006,0.08589685,0.12103647,0.15617609,0.19131571,0.22645533,0.26159495,0.22255093,0.1835069,0.14055848,0.10151446,0.062470436,0.10932326,0.15617609,0.20693332,0.25378615,0.30063897,0.60518235,0.9097257,1.2142692,1.5188124,1.8233559,2.0068626,2.1864653,2.366068,2.5456703,2.7252727,3.1157131,3.506153,3.8965936,4.283129,4.6735697,5.169429,5.661383,6.153338,6.6452928,7.137247,6.98888,6.844417,6.6960497,6.547683,6.3993154,6.297801,6.196286,6.0908675,5.989353,5.8878384,7.2270484,8.566258,9.909373,11.248583,12.587793,14.602465,16.617136,18.631807,20.646479,22.66115,25.683159,28.701262,31.723269,34.74137,37.76338,39.196293,40.633114,42.06603,43.50285,44.935764,43.018703,41.097736,39.176773,37.255806,35.338745,32.773552,30.212265,27.650976,25.085785,22.524496,21.85294,21.181383,20.50592,19.834364,19.162806,19.123762,19.080814,19.041769,19.002726,18.963682,19.541533,20.119385,20.693333,21.271183,21.849035,0.38653582,0.46071947,0.5309987,0.60518235,0.679366,0.74964523,0.78088045,0.8160201,0.8472553,0.8784905,0.9136301,1.0034313,1.0932326,1.183034,1.2728351,1.3626363,1.4446288,1.5266213,1.6086137,1.6906061,1.7765031,1.7413634,1.7062237,1.6710842,1.6359446,1.6008049,1.542239,1.4836729,1.4290112,1.3704453,1.3118792,3.3812122,5.4505453,7.523783,9.593117,11.66245,10.565312,9.468176,8.371038,7.2739015,6.1767645,5.708236,5.239708,4.7711797,4.3065557,3.8380275,3.521771,3.2094188,2.893162,2.5769055,2.260649,2.2567444,2.2489357,2.241127,2.233318,2.2255092,2.5183394,2.815074,3.1118085,3.4046388,3.7013733,4.5291066,5.3607445,6.1884775,7.0201154,7.8517528,7.492548,7.1333427,6.7780423,6.4188375,6.0635366,5.2084727,4.357313,3.506153,2.6510892,1.7999294,1.6945106,1.5890918,1.4836729,1.3782539,1.2767396,1.3470187,1.4212024,1.4914817,1.5656652,1.6359446,2.1513257,2.6667068,3.182088,3.697469,4.21285,4.83365,5.4505453,6.0713453,6.6921453,7.3129454,6.9225054,6.532065,6.141625,5.7511845,5.3607445,5.2475166,5.134289,5.017157,4.903929,4.786797,4.755562,4.7243266,4.689187,4.657952,4.6267166,4.3729305,4.1191444,3.8692627,3.6154766,3.3616903,3.174279,2.9868677,2.7994564,2.612045,2.4246337,2.5261483,2.6237583,2.7252727,2.8267872,2.9243972,2.7096553,2.494913,2.280171,2.0654287,1.8506867,2.069333,2.2840753,2.5027218,2.7213683,2.9361105,3.2211318,3.506153,3.7911747,4.0761957,4.3612175,4.661856,4.958591,5.2553253,5.55206,5.8487945,6.6140575,7.375416,8.136774,8.898132,9.663396,8.894228,8.121157,7.3519893,6.5828223,5.813655,5.559869,5.3060827,5.056201,4.802415,4.548629,5.4973984,6.446168,7.3910336,8.339804,9.288573,11.443803,13.602938,15.762072,17.917301,20.076437,21.821705,23.566973,25.308336,27.053604,28.79887,26.5187,24.23853,21.958359,19.678188,17.40192,17.70256,18.003199,18.307743,18.608381,18.912924,20.958832,23.000834,25.04674,27.092648,29.138554,30.938484,32.742317,34.54615,36.34608,38.149914,35.42074,32.695465,29.966288,27.241014,24.511837,24.29319,24.07845,23.859802,23.641155,23.426414,23.844185,24.25805,24.675823,25.093594,25.511364,22.813423,20.111576,17.413633,14.711788,12.013845,12.0489855,12.084125,12.119265,12.154405,12.185639,11.205634,10.22563,9.245625,8.265619,7.2856145,7.195813,7.1021075,7.008402,6.918601,6.824895,8.905942,10.983084,13.06413,15.145176,17.226223,15.582469,13.938716,12.298867,10.655114,9.01136,12.521418,16.02757,19.533724,23.043781,26.549934,21.583536,16.617136,11.6468315,6.6804323,1.7140326,1.6906061,1.6710842,1.6515622,1.6320401,1.6125181,1.9600099,2.3075018,2.6549935,3.0024853,3.349977,5.6691923,7.984503,10.303718,12.619028,14.938243,14.723501,14.508759,14.294017,14.079274,13.860628,12.419904,10.979179,9.534551,8.093826,6.649197,10.206107,13.763018,17.323833,20.880743,24.437654,24.644587,24.85152,25.058455,25.26929,25.476225,24.88666,24.29319,23.703627,23.114061,22.524496,22.0833,21.638197,21.197,20.755802,20.310701,19.709423,19.108145,18.502962,17.901684,17.300406,16.246218,15.188125,14.133936,13.079747,12.025558,12.587793,13.150026,13.712261,14.274494,14.836729,13.001659,11.166591,9.331521,7.4964523,5.661383,5.2748475,4.8883114,4.5017757,4.1113358,3.7247996,4.31046,4.8961205,5.481781,6.0635366,6.649197,6.1494336,5.645766,5.142098,4.6384296,4.138666,4.279225,4.415879,4.5564375,4.6969957,4.8375545,4.2362766,3.638903,3.0376248,2.436347,1.8389735,2.8072653,3.775557,4.747753,5.716045,6.688241,6.141625,5.5989127,5.0522966,4.50568,3.9629683,6.719476,9.47208,12.228588,14.981192,17.7377,14.571229,11.408664,8.242193,5.0757227,1.9131571,2.0420024,2.1708477,2.3035975,2.4324427,2.5612879,2.5456703,2.533957,2.5183394,2.5027218,2.4871042,3.9161155,5.349031,6.7780423,8.207053,9.636065,10.249056,10.862047,11.475039,12.08803,12.70102,12.693212,12.689307,12.685403,12.681499,12.67369,11.553126,10.436467,9.315904,8.19534,7.0747766,14.204215,21.333654,28.466997,35.596436,42.725872,36.72871,30.73155,24.730484,18.733322,12.73616,12.228588,11.721016,11.213444,10.705871,10.198298,9.561881,8.925464,8.289046,7.648724,7.012306,6.5008297,5.9932575,5.481781,4.9742084,4.462732,4.415879,4.369026,4.318269,4.271416,4.224563,3.6154766,3.0063896,2.3933985,1.7843118,1.175225,2.0888553,2.998581,3.912211,4.825841,5.735567,5.3295093,4.9234514,4.513489,4.1074314,3.7013733,3.7130866,3.7287042,3.7443218,3.7599394,3.775557,4.365122,4.9546866,5.5442514,6.133816,6.7233806,5.520825,4.3143644,3.1118085,1.9053483,0.698888,1.6554666,2.6081407,3.5647192,4.521298,5.473972,4.380739,3.2836022,2.1903696,1.0932326,0.0,0.0,0.0,0.0,0.0,0.0,1.9053483,3.8106966,5.716045,7.621393,9.526741,7.7541428,5.985449,4.2167544,2.4441557,0.6754616,0.59346914,0.5114767,0.42557985,0.3435874,0.26159495,0.21083772,0.15617609,0.10541886,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.78868926,1.5812829,2.3699722,3.1586614,3.951255,3.260176,2.5690966,1.8780174,1.1908426,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.13665408,0.23426414,0.3318742,0.42557985,0.5231899,0.5231899,0.5231899,0.5231899,0.5231899,0.5231899,0.61689556,0.7066968,0.79649806,0.8862993,0.97610056,0.94876975,0.92143893,0.8941081,0.8667773,0.8394465,0.6910792,0.5427119,0.39434463,0.24597734,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.19131571,0.3357786,0.47633708,0.62079996,0.76135844,0.6910792,0.61689556,0.5466163,0.47243267,0.39824903,0.39044023,0.37872702,0.3709182,0.359205,0.3513962,0.42167544,0.4958591,0.5661383,0.64032197,0.7106012,0.60518235,0.4958591,0.39044023,0.28111696,0.1756981,0.16008049,0.14446288,0.12884527,0.113227665,0.10151446,0.14055848,0.1796025,0.21864653,0.26159495,0.30063897,0.25378615,0.20693332,0.15617609,0.10932326,0.062470436,0.08980125,0.11713207,0.14446288,0.1717937,0.19912452,0.43338865,0.6637484,0.8980125,1.1283722,1.3626363,1.620327,1.8780174,2.135708,2.3933985,2.6510892,2.998581,3.3460727,3.6935644,4.041056,4.388548,5.1577153,5.9268827,6.6960497,7.4691215,8.238289,7.910319,7.5823493,7.2543793,6.9264097,6.5984397,6.426646,6.2548523,6.083059,5.911265,5.735567,6.774138,7.8088045,8.843472,9.878138,10.912805,12.521418,14.133936,15.74255,17.351164,18.963682,21.528873,24.097971,26.663162,29.23226,31.801357,33.97611,36.154766,38.33342,40.508175,42.68683,40.90642,39.126015,37.345608,35.569103,33.788696,31.676416,29.564135,27.451853,25.339571,23.223385,22.66115,22.095013,21.528873,20.96664,20.400501,20.35365,20.306797,20.256039,20.209187,20.162333,20.783133,21.407837,22.028637,22.653341,23.274141,0.28892577,0.3670138,0.44900626,0.5270943,0.60908675,0.6871748,0.7106012,0.7340276,0.75354964,0.77697605,0.80040246,0.8433509,0.8902037,0.93315214,0.98000497,1.0268579,1.1361811,1.2455044,1.3548276,1.4641509,1.5734742,1.5188124,1.4641509,1.4094892,1.3548276,1.3001659,1.2533131,1.2064602,1.1557031,1.1088502,1.0619974,3.4866312,5.9073606,8.331994,10.752724,13.173453,11.896713,10.61607,9.335425,8.054782,6.774138,6.196286,5.618435,5.040583,4.466636,3.8887846,3.5803368,3.2718892,2.9634414,2.6588979,2.35045,2.3035975,2.2567444,2.2059872,2.1591344,2.1122816,2.4597735,2.8072653,3.154757,3.5022488,3.8497405,4.7633705,5.6809053,6.5945354,7.5081654,8.4257,7.914223,7.406651,6.8951745,6.3836975,5.8761253,5.056201,4.2362766,3.416352,2.5964274,1.7765031,1.6593709,1.5461433,1.4290112,1.3157835,1.1986516,1.1908426,1.1869383,1.1791295,1.1713207,1.1635119,1.9092526,2.6510892,3.39683,4.142571,4.8883114,5.196759,5.5091114,5.8175592,6.126007,6.4383593,6.028397,5.6223392,5.2162814,4.806319,4.4002614,4.478349,4.560342,4.6384296,4.7204223,4.7985106,4.7399445,4.6813784,4.618908,4.560342,4.5017757,4.142571,3.7833657,3.4280653,3.06886,2.7135596,2.639376,2.5612879,2.4871042,2.4129205,2.338737,2.3855898,2.436347,2.4871042,2.5378613,2.5886188,2.3816853,2.1708477,1.9639144,1.756981,1.5500476,1.5890918,1.6281357,1.6710842,1.7101282,1.7491722,2.241127,2.7330816,3.2289407,3.7208953,4.21285,4.454923,4.6969957,4.939069,5.181142,5.423215,6.785851,8.148487,9.511124,10.87376,12.236397,11.150972,10.069453,8.98403,7.898606,6.813182,6.180669,5.548156,4.9156423,4.283129,3.6506162,4.9546866,6.2587566,7.5667315,8.870802,10.174872,13.173453,16.168129,19.16671,22.16529,25.163872,27.420616,29.681267,31.941916,34.202564,36.46321,33.324074,30.18103,27.04189,23.90275,20.76361,20.53325,20.30289,20.072533,19.842173,19.611813,21.372698,23.133583,24.894468,26.65145,28.412334,30.946293,33.476345,36.010303,38.54426,41.07431,37.279232,33.484154,29.689075,25.893995,22.098917,22.0833,22.071587,22.05597,22.04035,22.024733,22.46593,22.903223,23.344421,23.785618,24.226816,21.610867,18.998821,16.386776,13.774731,11.162686,11.229061,11.29934,11.365715,11.43209,11.498465,10.135828,8.769287,7.406651,6.04011,4.6735697,4.7087092,4.743849,4.7789884,4.814128,4.8492675,5.6652875,6.481308,7.2934237,8.109444,8.925464,8.234385,7.5433054,6.8561306,6.165051,5.473972,10.748819,16.019762,21.29461,26.565554,31.836496,25.687063,19.533724,13.380386,7.2270484,1.0737107,1.2415999,1.4055848,1.5695697,1.7335546,1.901444,2.330928,2.7604125,3.1898966,3.619381,4.0488653,6.9771667,9.905469,12.83377,15.758167,18.68647,16.792833,14.899199,13.001659,11.108025,9.2104845,8.55845,7.9064145,7.2543793,6.602344,5.950309,9.6243515,13.29449,16.968533,20.63867,24.312714,25.159967,26.007223,26.854479,27.701735,28.548988,26.97942,25.40985,23.84028,22.27071,20.701141,19.799223,18.893402,17.991486,17.08957,16.187653,15.844065,15.4965725,15.152986,14.809398,14.461906,13.622459,12.783013,11.943566,11.10412,10.260769,10.373997,10.487225,10.600452,10.71368,10.823003,10.034314,9.24172,8.449126,7.656533,6.8639393,5.8761253,4.8883114,3.900498,2.912684,1.9248703,2.9556324,3.9863946,5.0132523,6.044015,7.0747766,6.606249,6.133816,5.6652875,5.196759,4.7243266,4.794606,4.8648853,4.9351645,5.0054436,5.0757227,4.4002614,3.7247996,3.049338,2.3738766,1.698415,2.5964274,3.49444,4.3924527,5.290465,6.1884775,5.4036927,4.618908,3.8341231,3.049338,2.260649,5.727758,9.190963,12.658072,16.121277,19.588387,15.992432,12.396477,8.800523,5.2084727,1.6125181,1.6906061,1.7686942,1.8467822,1.9209659,1.999054,2.018576,2.0341935,2.0537157,2.069333,2.0888553,2.9283018,3.767748,4.607195,5.446641,6.2860875,6.5125427,6.7389984,6.9615493,7.1880045,7.4105554,7.859562,8.308568,8.75367,9.202676,9.651682,8.4257,7.2036223,5.9815445,4.759466,3.5373883,12.90405,22.266806,31.633467,40.996223,50.362885,42.183163,34.00344,25.823717,17.643993,9.464272,10.053836,10.6434,11.232965,11.82253,12.412095,11.100216,9.788337,8.476458,7.1606736,5.8487945,5.134289,4.415879,3.697469,2.979059,2.260649,2.2450314,2.2294137,2.2098918,2.194274,2.174752,1.8584955,1.5383345,1.2220778,0.9058213,0.58566034,1.698415,2.8111696,3.9239242,5.036679,6.1494336,5.290465,4.4314966,3.5686235,2.7096553,1.8506867,1.8584955,1.8663043,1.8741131,1.8819219,1.8858263,2.182561,2.4792955,2.7721257,3.06886,3.3616903,2.8463092,2.330928,1.815547,1.3040704,0.78868926,1.815547,2.8424048,3.8692627,4.8961205,5.9268827,4.7399445,3.5569105,2.3699722,1.183034,0.0,0.0,0.0,0.0,0.0,0.0,0.96438736,1.9287747,2.893162,3.8614538,4.825841,4.041056,3.2562714,2.4714866,1.6867018,0.9019169,0.78868926,0.679366,0.5700427,0.46071947,0.3513962,0.28111696,0.21083772,0.14055848,0.07027924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.43338865,0.8667773,1.2962615,1.7296503,2.1630387,1.815547,1.4719596,1.1283722,0.78088045,0.43729305,0.3513962,0.26159495,0.1756981,0.08589685,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.1678893,0.28502136,0.40215343,0.5192855,0.63641757,0.57394713,0.5114767,0.44900626,0.38653582,0.3240654,0.45681506,0.58956474,0.7223144,0.8550641,0.9878138,1.0034313,1.0229534,1.038571,1.0580931,1.0737107,0.8823949,0.6910792,0.4958591,0.30454338,0.113227665,0.093705654,0.078088045,0.058566034,0.042948425,0.023426414,0.1639849,0.30454338,0.44510186,0.58566034,0.7262188,0.6715572,0.61689556,0.5583295,0.5036679,0.44900626,0.43338865,0.41386664,0.39824903,0.37872702,0.3631094,0.42948425,0.4958591,0.5661383,0.63251317,0.698888,0.60127795,0.5036679,0.40605783,0.30844778,0.21083772,0.19131571,0.1717937,0.15227169,0.13274968,0.113227665,0.15617609,0.20302892,0.24597734,0.29283017,0.3357786,0.28111696,0.22645533,0.1717937,0.11713207,0.062470436,0.07027924,0.078088045,0.08589685,0.093705654,0.10151446,0.26159495,0.42167544,0.58175594,0.7418364,0.9019169,1.2337911,1.5695697,1.9053483,2.241127,2.5769055,2.8814487,3.1859922,3.4905357,3.795079,4.0996222,5.1460023,6.196286,7.2426662,8.289046,9.339331,8.831758,8.324185,7.816613,7.309041,6.801469,6.559396,6.3134184,6.0713453,5.8292727,5.5871997,6.3173227,7.0474463,7.7775693,8.507692,9.237816,10.444276,11.6468315,12.853292,14.055848,15.262308,17.378494,19.490776,21.606962,23.723148,25.839334,28.755922,31.676416,34.59691,37.517403,40.437893,38.798046,37.158195,35.51835,33.878498,32.23865,30.575375,28.912098,27.248823,25.589453,23.926178,23.469362,23.008642,22.551826,22.095013,21.638197,21.583536,21.528873,21.474213,21.415646,21.360985,22.028637,22.696291,23.363943,24.031595,24.69925,0.18741131,0.27330816,0.3631094,0.44900626,0.5388075,0.62470436,0.63641757,0.6481308,0.6637484,0.6754616,0.6871748,0.6871748,0.6871748,0.6871748,0.6871748,0.6871748,0.8238289,0.96438736,1.1010414,1.2376955,1.3743496,1.3001659,1.2259823,1.1517987,1.0737107,0.999527,0.96438736,0.92534333,0.8862993,0.8511597,0.81211567,3.5881457,6.364176,9.136301,11.912332,14.688361,13.224211,11.763964,10.299813,8.835662,7.375416,6.688241,6.001066,5.3138914,4.6267166,3.9356375,3.638903,3.338264,3.0376248,2.736986,2.436347,2.35045,2.260649,2.174752,2.0888553,1.999054,2.4012074,2.7994564,3.2016098,3.5998588,3.998108,5.001539,6.001066,7.000593,8.00012,8.999647,8.335898,7.676055,7.012306,6.348558,5.688714,4.900025,4.1113358,3.3265507,2.5378613,1.7491722,1.6242313,1.4992905,1.3743496,1.2494087,1.1244678,1.038571,0.94876975,0.8628729,0.77307165,0.6871748,1.6632754,2.639376,3.611572,4.5876727,5.563773,5.563773,5.563773,5.563773,5.563773,5.563773,5.138193,4.7126136,4.2870336,3.8614538,3.435874,3.7130866,3.9863946,4.263607,4.5369153,4.814128,4.7243266,4.6384296,4.548629,4.462732,4.376835,3.912211,3.4514916,2.9868677,2.5261483,2.0615244,2.1005683,2.135708,2.174752,2.2137961,2.2489357,2.2489357,2.2489357,2.2489357,2.2489357,2.2489357,2.0498111,1.8506867,1.6515622,1.4485333,1.2494087,1.1127546,0.97610056,0.8394465,0.698888,0.5622339,1.261122,1.9639144,2.6628022,3.3616903,4.0605783,4.251894,4.4393053,4.6267166,4.814128,5.001539,6.9615493,8.925464,10.889378,12.849388,14.813302,13.411622,12.013845,10.612165,9.21439,7.812709,6.801469,5.786324,4.775084,3.7638438,2.7486992,4.4119744,6.0752497,7.7385254,9.4018,11.061172,14.899199,18.737226,22.575254,26.41328,30.251308,33.023434,35.799465,38.575493,41.351524,44.12365,40.12554,36.12353,32.125423,28.12341,24.125301,23.363943,22.59868,21.837322,21.075964,20.310701,21.786564,23.262428,24.738293,26.214157,27.686117,30.950197,34.214275,37.474453,40.738533,43.99871,39.13773,34.27675,29.411861,24.55088,19.685997,19.873407,20.06082,20.24823,20.435642,20.623053,21.087677,21.548395,22.01302,22.47374,22.938364,20.412214,17.886066,15.363823,12.837675,10.311526,10.413041,10.510651,10.612165,10.71368,10.81129,9.062118,7.3129454,5.563773,3.8106966,2.0615244,2.2255092,2.3855898,2.5495746,2.7135596,2.87364,2.4246337,1.9756275,1.5266213,1.0737107,0.62470436,0.8862993,1.1517987,1.4133936,1.6749885,1.9365835,8.976221,16.011953,23.05159,30.087324,37.12306,29.786684,22.450314,15.113941,7.773665,0.43729305,0.78868926,1.1361811,1.4875772,1.8389735,2.1864653,2.7018464,3.213323,3.7247996,4.2362766,4.7516575,8.289046,11.826434,15.363823,18.90121,22.4386,18.862167,15.285735,11.713207,8.136774,4.564246,4.7009,4.8375545,4.9742084,5.1108627,5.251421,9.0386915,12.825961,16.613232,20.400501,24.187773,25.67535,27.162926,28.650503,30.13808,31.625658,29.076084,26.526508,23.97303,21.423454,18.87388,17.511244,16.148607,14.785972,13.423335,12.0606985,11.974802,11.888905,11.799104,11.713207,11.623405,10.998701,10.373997,9.749292,9.124588,8.499884,8.164105,7.824422,7.4886436,7.1489606,6.813182,7.0630636,7.3129454,7.562827,7.812709,8.062591,6.473499,4.8883114,3.2992198,1.7140326,0.12494087,1.6008049,3.076669,4.548629,6.0244927,7.5003567,7.0630636,6.6257706,6.1884775,5.7511845,5.3138914,5.3138914,5.3138914,5.3138914,5.3138914,5.3138914,4.564246,3.8106966,3.0610514,2.3114061,1.5617609,2.3894942,3.213323,4.037152,4.860981,5.688714,4.661856,3.638903,2.612045,1.5890918,0.5622339,4.73604,8.913751,13.087557,17.261362,21.439074,17.413633,13.388195,9.362757,5.337318,1.3118792,1.33921,1.3626363,1.3860629,1.4133936,1.43682,1.4875772,1.5383345,1.5890918,1.6359446,1.6867018,1.9365835,2.1864653,2.436347,2.6862288,2.9361105,2.77603,2.612045,2.4480603,2.2879796,2.1239948,3.0259118,3.9239242,4.825841,5.7238536,6.6257706,5.298274,3.9746814,2.6510892,1.3235924,0.0,11.599979,23.199959,34.79994,46.399918,57.999897,47.63761,37.27533,26.913044,16.55076,6.1884775,7.8751793,9.561881,11.248583,12.939189,14.625891,12.63855,10.651209,8.663869,6.676528,4.689187,3.7638438,2.8385005,1.9131571,0.9878138,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,1.3118792,2.6237583,3.9356375,5.251421,6.5633,5.251421,3.9356375,2.6237583,1.3118792,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1756981,0.3513962,0.5231899,0.698888,0.8745861,1.9756275,3.076669,4.173806,5.2748475,6.375889,5.099149,3.8263142,2.5495746,1.2767396,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.3240654,0.5231899,0.7262188,0.92534333,1.1244678,0.9878138,0.8511597,0.7106012,0.57394713,0.43729305,0.3513962,0.26159495,0.1756981,0.08589685,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.19912452,0.3357786,0.47633708,0.61299115,0.74964523,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.30063897,0.47633708,0.6481308,0.8238289,0.999527,1.0619974,1.1244678,1.1869383,1.2494087,1.3118792,1.0737107,0.8394465,0.60127795,0.3631094,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.13665408,0.27330816,0.41386664,0.5505207,0.6871748,0.6481308,0.61299115,0.57394713,0.5388075,0.4997635,0.47633708,0.44900626,0.42557985,0.39824903,0.37482262,0.43729305,0.4997635,0.5622339,0.62470436,0.6871748,0.60127795,0.5114767,0.42557985,0.3357786,0.24988174,0.22645533,0.19912452,0.1756981,0.14836729,0.12494087,0.1756981,0.22645533,0.27330816,0.3240654,0.37482262,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.8511597,1.261122,1.6749885,2.0888553,2.4988174,2.7643168,3.0259118,3.2875066,3.5491016,3.8106966,5.138193,6.461786,7.7892823,9.112875,10.436467,9.749292,9.062118,8.374943,7.687768,7.000593,6.688241,6.375889,6.0635366,5.7511845,5.4388323,5.8644123,6.2860875,6.7116675,7.137247,7.562827,8.36323,9.163632,9.964035,10.760532,11.560935,13.224211,14.8874855,16.55076,18.214037,19.873407,23.53964,27.201971,30.8643,34.52663,38.188957,36.685764,35.186474,33.687183,32.187893,30.688602,29.474333,28.263968,27.049698,25.839334,24.625065,24.273668,23.926178,23.574781,23.223385,22.875893,22.813423,22.750952,22.688482,22.62601,22.563541,23.274141,23.988647,24.69925,25.413754,26.124355,0.14836729,0.22645533,0.30454338,0.38263142,0.46071947,0.5388075,0.5583295,0.58175594,0.60518235,0.62860876,0.6481308,0.63641757,0.62470436,0.61299115,0.60127795,0.58566034,0.71841,0.8472553,0.97610056,1.1088502,1.2376955,1.183034,1.1283722,1.0737107,1.0190489,0.96438736,1.0229534,1.0815194,1.1439898,1.2025559,1.261122,3.4827268,5.704332,7.9220324,10.143637,12.361338,11.615597,10.87376,10.128019,9.382278,8.636538,7.6955767,6.75852,5.8175592,4.8765984,3.9356375,3.619381,3.3031244,2.9868677,2.6667068,2.35045,2.2567444,2.1591344,2.0654287,1.9717231,1.8741131,2.2840753,2.6940374,3.1039999,3.513962,3.9239242,4.7243266,5.5247293,6.3251314,7.125534,7.9259367,7.328563,6.735094,6.141625,5.5442514,4.950782,4.31046,3.6701381,3.0298162,2.3894942,1.7491722,1.6125181,1.475864,1.33921,1.1986516,1.0619974,1.1478943,1.2337911,1.3157835,1.4016805,1.4875772,2.3738766,3.2640803,4.1503797,5.036679,5.9268827,5.8644123,5.805846,5.743376,5.6848097,5.6262436,5.196759,4.7711797,4.3416953,3.9161155,3.4866312,3.7247996,3.9629683,4.2011366,4.4393053,4.6735697,4.533011,4.388548,4.2479897,4.1035266,3.9629683,3.8263142,3.6857557,3.5491016,3.4124475,3.2757936,3.1157131,2.959537,2.803361,2.6432803,2.4871042,2.3738766,2.2567444,2.1435168,2.0263848,1.9131571,1.7491722,1.5890918,1.4251068,1.261122,1.1010414,1.2572175,1.4133936,1.5734742,1.7296503,1.8858263,2.6159496,3.3460727,4.0761957,4.806319,5.5364423,5.9425,6.348558,6.7507114,7.1567693,7.562827,9.460366,11.357906,13.2554455,15.152986,17.050524,16.43363,15.816733,15.195933,14.579038,13.962143,12.458947,10.955752,9.456462,7.9532676,6.4500723,8.484266,10.514555,12.548749,14.579038,16.613232,19.959305,23.305378,26.655354,30.001427,33.351402,34.59691,35.83851,37.08401,38.329517,39.57502,36.209427,32.84383,29.478237,26.116547,22.750952,21.997402,21.243853,20.494207,19.740658,18.987108,20.15062,21.314133,22.47374,23.63725,24.800762,27.631454,30.466051,33.29674,36.13134,38.96203,34.432922,29.903816,25.370806,20.8417,16.312593,17.526861,18.74113,19.959305,21.173573,22.387842,21.888079,21.388315,20.888552,20.388788,19.889025,19.151093,18.417065,17.683039,16.94901,16.211079,15.816733,15.418485,15.020235,14.621986,14.223738,12.993851,11.760059,10.526268,9.296382,8.062591,7.027924,5.9932575,4.958591,3.9239242,2.8892577,3.3616903,3.8341231,4.3065557,4.7789884,5.251421,8.39056,11.533605,14.676648,17.819693,20.962736,23.340517,25.722202,28.103888,30.481668,32.863354,26.948185,21.033014,15.117846,9.202676,3.2875066,3.0727646,2.8580225,2.6432803,2.4285383,2.2137961,3.7638438,5.3138914,6.8639393,8.413987,9.964035,11.924045,13.887959,15.851873,17.811884,19.775797,17.530766,15.285735,13.040704,10.795672,8.550641,7.8790836,7.211431,6.5398736,5.8683167,5.2006636,8.659965,12.119265,15.578565,19.041769,22.50107,23.453745,24.410322,25.366901,26.319576,27.276154,26.405472,25.53479,24.664108,23.793427,22.926651,20.935406,18.94416,16.95682,14.965574,12.974329,12.786918,12.595602,12.404286,12.216875,12.025558,11.810817,11.599979,11.389141,11.174399,10.963562,10.0226,9.081639,8.140678,7.2036223,6.262661,7.3129454,8.36323,9.413514,10.4637985,11.514082,10.104593,8.699008,7.289519,5.883934,4.474445,4.7789884,5.083532,5.388075,5.6965227,6.001066,6.2040954,6.4110284,6.6140575,6.8209906,7.0240197,6.7233806,6.426646,6.126007,5.825368,5.5247293,4.786797,4.0488653,3.310933,2.5769055,1.8389735,2.4246337,3.0141985,3.5998588,4.1894236,4.775084,4.3455997,3.9161155,3.4866312,3.0532427,2.6237583,6.6726236,10.721489,14.766449,18.815315,22.86418,18.709896,14.559516,10.405232,6.250948,2.1005683,1.9131571,1.7257458,1.5383345,1.3509232,1.1635119,1.3899672,1.6164225,1.8467822,2.0732377,2.2996929,2.4441557,2.5886188,2.7330816,2.8814487,3.0259118,2.8189783,2.6081407,2.4012074,2.194274,1.9873407,3.9824903,5.9776397,7.9727893,9.967939,11.963089,9.612638,7.262188,4.911738,2.5612879,0.21083772,9.515028,18.81922,28.119505,37.423695,46.72398,39.383705,32.04343,24.703154,17.366781,10.0265045,10.561408,11.096312,11.631214,12.166118,12.70102,12.232492,11.763964,11.29934,10.8308115,10.362284,8.335898,6.3056097,4.279225,2.25284,0.22645533,0.19912452,0.1756981,0.14836729,0.12494087,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,1.1010414,2.1981785,3.2992198,4.4002614,5.5013027,4.4705405,3.4436827,2.416825,1.3899672,0.3631094,0.42167544,0.47633708,0.5349031,0.59346914,0.6481308,0.5192855,0.39044023,0.26159495,0.12884527,0.0,0.14055848,0.28111696,0.42167544,0.5583295,0.698888,1.5812829,2.463678,3.3460727,4.2284675,5.1108627,4.1035266,3.096191,2.0888553,1.0815194,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.3318742,0.47243267,0.61689556,0.75745404,0.9019169,0.79259366,0.6832704,0.57785153,0.46852827,0.3631094,0.29283017,0.22255093,0.15227169,0.08199245,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.30063897,0.30063897,0.30063897,0.30063897,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.21083772,0.359205,0.5036679,0.6520352,0.80040246,0.659844,0.5192855,0.37872702,0.23816854,0.10151446,0.25378615,0.40996224,0.5661383,0.71841,0.8745861,0.96829176,1.0580931,1.1517987,1.2455044,1.33921,1.116659,0.8980125,0.679366,0.45681506,0.23816854,0.19131571,0.14055848,0.093705654,0.046852827,0.0,0.11713207,0.23426414,0.3513962,0.46852827,0.58566034,0.58566034,0.58175594,0.58175594,0.57785153,0.57394713,0.5466163,0.5192855,0.49195468,0.46462387,0.43729305,0.4958591,0.5583295,0.61689556,0.679366,0.737932,0.64032197,0.5427119,0.44510186,0.3474918,0.24988174,0.23426414,0.21864653,0.20693332,0.19131571,0.1756981,0.24988174,0.3240654,0.39824903,0.47633708,0.5505207,0.46462387,0.37872702,0.29673457,0.21083772,0.12494087,0.10151446,0.078088045,0.058566034,0.03513962,0.011713207,0.08589685,0.15617609,0.23035973,0.30063897,0.37482262,0.7223144,1.0698062,1.4172981,1.7647898,2.1122816,2.338737,2.5690966,2.795552,3.0220075,3.2484627,4.3260775,5.4036927,6.481308,7.558923,8.636538,8.437413,8.238289,8.039165,7.8361354,7.6370106,7.172387,6.707763,6.2431393,5.7785153,5.3138914,5.8487945,6.3836975,6.918601,7.453504,7.988407,8.902037,9.815667,10.733202,11.6468315,12.564366,13.884054,15.207646,16.531239,17.850927,19.174519,22.106726,25.03893,27.971138,30.903343,33.839455,32.61738,31.399202,30.177126,28.958952,27.736874,27.045794,26.350811,25.65973,24.968653,24.273668,24.3908,24.504028,24.62116,24.734388,24.85152,24.941322,25.035027,25.128733,25.218534,25.31224,25.687063,26.061886,26.436708,26.811531,27.186354,0.113227665,0.1796025,0.24597734,0.31625658,0.38263142,0.44900626,0.48414588,0.5153811,0.5466163,0.58175594,0.61299115,0.58566034,0.5622339,0.5388075,0.5114767,0.48805028,0.60908675,0.7340276,0.8550641,0.97610056,1.1010414,1.0659018,1.0307622,0.9956226,0.96048295,0.92534333,1.0815194,1.2415999,1.397776,1.5539521,1.7140326,3.377308,5.040583,6.707763,8.371038,10.0382185,10.010887,9.983557,9.956225,9.928895,9.901564,8.706817,7.5159745,6.321227,5.1303844,3.9356375,3.6037633,3.2679846,2.9322062,2.5964274,2.260649,2.1591344,2.05762,1.9561055,1.8506867,1.7491722,2.1708477,2.5886188,3.0102942,3.4280653,3.8497405,4.4510183,5.0483923,5.64967,6.250948,6.8483214,6.321227,5.794133,5.267039,4.7399445,4.21285,3.7208953,3.2289407,2.7330816,2.241127,1.7491722,1.6008049,1.4485333,1.3001659,1.1517987,0.999527,1.2572175,1.5149081,1.7725986,2.0302892,2.2879796,3.0883822,3.8887846,4.689187,5.4856853,6.2860875,6.168956,6.0479193,5.9268827,5.805846,5.688714,5.2592297,4.825841,4.396357,3.9668727,3.5373883,3.736513,3.9356375,4.138666,4.337791,4.5369153,4.3416953,4.142571,3.9434462,3.7482262,3.5491016,3.736513,3.9239242,4.1113358,4.298747,4.4861584,4.134762,3.7833657,3.4280653,3.076669,2.7252727,2.494913,2.2645533,2.0341935,1.8038338,1.5734742,1.4485333,1.3235924,1.1986516,1.0737107,0.94876975,1.4016805,1.8545911,2.3075018,2.7604125,3.213323,3.970777,4.732136,5.493494,6.250948,7.012306,7.633106,8.257811,8.878611,9.503315,10.124115,11.959184,13.790349,15.621513,17.456583,19.287746,19.451733,19.615717,19.783606,19.947592,20.111576,18.12033,16.129086,14.133936,12.142691,10.151445,12.552653,14.95386,17.358973,19.76018,22.161386,25.01941,27.877432,30.735455,33.593475,36.4515,36.166477,35.88146,35.596436,35.311413,35.026394,32.293312,29.564135,26.834957,24.10578,21.376602,20.630861,19.889025,19.147188,18.405352,17.663515,18.51077,19.36193,20.21309,21.06425,21.911505,24.316618,26.717825,29.119032,31.524143,33.92535,29.728119,25.530886,21.333654,17.136421,12.939189,15.180316,17.421442,19.666473,21.9076,24.148727,22.688482,21.22433,19.764084,18.299932,16.835783,17.893875,18.948065,20.002253,21.056442,22.11063,21.216522,20.322414,19.428307,18.534197,17.636185,16.921679,16.207174,15.492668,14.778163,14.063657,11.8303385,9.597021,7.363703,5.134289,2.900971,4.2948427,5.688714,7.08649,8.480362,9.874233,15.8987255,21.919313,27.943808,33.964394,39.988888,37.708717,35.43245,33.156185,30.876013,28.599747,24.10578,19.615717,15.12175,10.631687,6.13772,5.35684,4.575959,3.7989833,3.018103,2.2372224,4.825841,7.4105554,9.999174,12.587793,15.176412,15.562947,15.949483,16.33602,16.72646,17.112995,16.199366,15.281831,14.3682,13.450665,12.537036,11.061172,9.581403,8.105539,6.6257706,5.1499066,8.281238,11.416472,14.547803,17.679134,20.81437,21.236044,21.657719,22.079395,22.50107,22.926651,23.734861,24.543072,25.355188,26.163399,26.975515,24.355661,21.739712,19.123762,16.503908,13.887959,13.595129,13.302299,13.009468,12.716639,12.423808,12.626837,12.825961,13.025085,13.224211,13.423335,11.881096,10.338858,8.796618,7.2543793,5.7121406,7.562827,9.413514,11.2642,13.110983,14.96167,13.735687,12.5058,11.279819,10.053836,8.823949,7.9610763,7.094299,6.2314262,5.364649,4.5017757,5.349031,6.196286,7.043542,7.890797,8.738052,8.136774,7.5394006,6.9381227,6.336845,5.735567,5.0132523,4.2870336,3.5608149,2.8385005,2.1122816,2.463678,2.8111696,3.1625657,3.513962,3.8614538,4.029343,4.193328,4.357313,4.521298,4.689187,8.609207,12.529227,16.449247,20.369267,24.289286,20.006157,15.726933,11.447707,7.168483,2.8892577,2.4871042,2.0888553,1.6867018,1.2884527,0.8862993,1.2923572,1.698415,2.1005683,2.5066261,2.912684,2.951728,2.9907722,3.0337205,3.0727646,3.1118085,2.8619268,2.6081407,2.3543546,2.1005683,1.8506867,4.939069,8.031356,11.119738,14.212025,17.300406,13.923099,10.549695,7.1762915,3.7989833,0.42557985,7.4300776,14.434575,21.439074,28.443571,35.448067,31.133703,26.815435,22.497166,18.178898,13.860628,13.243732,12.626837,12.009941,11.393045,10.77615,11.826434,12.880623,13.930907,14.985096,16.039284,12.907954,9.776623,6.649197,3.5178664,0.38653582,0.3240654,0.26159495,0.19912452,0.13665408,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.8862993,1.7765031,2.6628022,3.5491016,4.4393053,3.6935644,2.951728,2.2098918,1.4680552,0.7262188,0.8394465,0.95657855,1.0698062,1.1869383,1.3001659,1.038571,0.78088045,0.5192855,0.26159495,0.0,0.10541886,0.21083772,0.31625658,0.42167544,0.5231899,1.1908426,1.8545911,2.5183394,3.1859922,3.8497405,3.1118085,2.3699722,1.6281357,0.8902037,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.3357786,0.42167544,0.5036679,0.58956474,0.6754616,0.59737355,0.5192855,0.44119745,0.3631094,0.28892577,0.23426414,0.1835069,0.12884527,0.078088045,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.08980125,0.13665408,0.1796025,0.22645533,0.22645533,0.22645533,0.22645533,0.22645533,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.21864653,0.37872702,0.5349031,0.6910792,0.8511597,0.6949836,0.5388075,0.38653582,0.23035973,0.07418364,0.21083772,0.3435874,0.48024148,0.61689556,0.74964523,0.8706817,0.9956226,1.116659,1.2415999,1.3626363,1.1596074,0.95657855,0.75354964,0.5544251,0.3513962,0.28111696,0.21083772,0.14055848,0.07027924,0.0,0.09761006,0.19522011,0.29283017,0.39044023,0.48805028,0.5192855,0.5544251,0.58566034,0.61689556,0.6481308,0.62079996,0.58956474,0.5583295,0.5309987,0.4997635,0.5583295,0.61689556,0.6715572,0.7301232,0.78868926,0.679366,0.57394713,0.46462387,0.359205,0.24988174,0.24597734,0.23816854,0.23426414,0.23035973,0.22645533,0.3240654,0.42557985,0.5231899,0.62470436,0.7262188,0.61689556,0.5114767,0.40215343,0.29673457,0.18741131,0.15617609,0.12103647,0.08980125,0.058566034,0.023426414,0.08199245,0.14055848,0.19912452,0.25378615,0.31235218,0.59346914,0.8784905,1.1596074,1.4407244,1.7257458,1.9170616,2.1083772,2.3035975,2.494913,2.6862288,3.5178664,4.349504,5.1772375,6.008875,6.8366084,7.125534,7.4144597,7.699481,7.988407,8.273428,7.656533,7.039637,6.422742,5.805846,5.1889505,5.833177,6.477403,7.1216297,7.7658563,8.413987,9.440845,10.471607,11.502369,12.533132,13.563893,14.543899,15.527808,16.511717,17.491722,18.475632,20.677715,22.879797,25.08188,27.283962,29.486046,28.548988,27.608028,26.667067,25.726107,24.78905,24.613352,24.441559,24.269764,24.097971,23.926178,24.504028,25.085785,25.663635,26.245392,26.823244,27.073126,27.319103,27.568985,27.814962,28.06094,28.099983,28.139027,28.174168,28.213211,28.24835,0.07418364,0.13274968,0.19131571,0.24597734,0.30454338,0.3631094,0.40605783,0.44900626,0.48805028,0.5309987,0.57394713,0.5388075,0.4997635,0.46071947,0.42557985,0.38653582,0.5036679,0.61689556,0.7340276,0.8472553,0.96438736,0.94876975,0.93315214,0.91753453,0.9019169,0.8862993,1.1439898,1.397776,1.6515622,1.9092526,2.1630387,3.2718892,4.380739,5.493494,6.602344,7.7111945,8.402273,9.093353,9.784432,10.471607,11.162686,9.718058,8.273428,6.8287997,5.3841705,3.9356375,3.5842414,3.232845,2.8814487,2.5261483,2.174752,2.0654287,1.9561055,1.8467822,1.7335546,1.6242313,2.0537157,2.4831998,2.9165885,3.3460727,3.775557,4.173806,4.575959,4.9742084,5.376362,5.774611,5.3138914,4.853172,4.396357,3.9356375,3.474918,3.1313305,2.7838387,2.4402514,2.096664,1.7491722,1.5890918,1.4251068,1.261122,1.1010414,0.93705654,1.3665408,1.796025,2.2294137,2.6588979,3.0883822,3.7989833,4.513489,5.22409,5.938596,6.649197,6.4695945,6.289992,6.1103897,5.930787,5.7511845,5.3177958,4.884407,4.4510183,4.0215344,3.5881457,3.7482262,3.912211,4.0761957,4.2362766,4.4002614,4.1464753,3.8965936,3.6428072,3.3890212,3.1391394,3.6506162,4.1620927,4.6735697,5.1889505,5.700427,5.153811,4.60329,4.056674,3.5100577,2.9634414,2.6159496,2.2723622,1.9287747,1.5812829,1.2376955,1.1517987,1.0619974,0.97610056,0.8862993,0.80040246,1.5461433,2.2957885,3.0415294,3.7911747,4.5369153,5.3256044,6.1181984,6.9068875,7.699481,8.488171,9.327617,10.167064,11.00651,11.845957,12.689307,14.454097,16.222792,17.991486,19.756275,21.52497,22.47374,23.418604,24.367374,25.316145,26.26101,23.781713,21.298513,18.815315,16.332115,13.848915,16.62104,19.393166,22.169195,24.941322,27.713448,30.079515,32.449486,34.815556,37.18162,39.551594,37.73605,35.9205,34.104954,32.289406,30.47386,28.3811,26.284435,24.191677,22.095013,19.998348,19.268225,18.534197,17.804073,17.070047,16.33602,16.874826,17.413633,17.948538,18.487345,19.026152,20.997875,22.969599,24.941322,26.913044,28.888672,25.023314,21.157955,17.292597,13.427239,9.561881,12.83377,16.101755,19.373644,22.641628,25.913517,23.488884,21.06425,18.635712,16.211079,13.786445,16.632753,19.479063,22.321468,25.167776,28.014086,26.620214,25.226343,23.836376,22.442505,21.048632,20.853413,20.654287,20.459068,20.259943,20.06082,16.632753,13.200784,9.772718,6.3407493,2.912684,5.2318993,7.5472097,9.866425,12.181735,14.50095,23.402987,32.305023,41.20706,50.1091,59.011135,52.076916,45.1427,38.20848,31.274261,24.33614,21.267279,18.19842,15.125654,12.056794,8.987934,7.6409154,6.297801,4.950782,3.6076677,2.260649,5.8878384,9.511124,13.138313,16.761599,20.388788,19.20185,18.011007,16.82407,15.637131,14.450192,14.864059,15.281831,15.695697,16.109564,16.52343,14.239355,11.955279,9.671205,7.3832245,5.099149,7.9064145,10.709775,13.513136,16.320402,19.123762,19.014439,18.905115,18.795792,18.68647,18.573242,21.06425,23.55526,26.046267,28.533371,31.02438,27.779821,24.535263,21.290705,18.046146,14.801589,14.40334,14.008995,13.614651,13.220306,12.825961,13.438952,14.051944,14.661031,15.274021,15.8870125,13.743496,11.596075,9.452558,7.309041,5.1616197,7.812709,10.4637985,13.110983,15.762072,18.41316,17.366781,16.316498,15.270117,14.223738,13.173453,11.139259,9.105066,7.0708723,5.036679,2.998581,4.4900627,5.9815445,7.4691215,8.960603,10.44818,9.550168,8.648251,7.7502384,6.8483214,5.950309,5.2358036,4.5252023,3.8106966,3.1000953,2.3855898,2.4988174,2.612045,2.7252727,2.8385005,2.951728,3.7091823,4.4705405,5.2318993,5.989353,6.7507114,10.541886,14.33306,18.12814,21.919313,25.714394,21.306324,16.898252,12.490183,8.082112,3.6740425,3.0610514,2.4519646,1.8389735,1.2259823,0.61299115,1.1947471,1.7765031,2.358259,2.9439192,3.5256753,3.4593005,3.39683,3.330455,3.2640803,3.2016098,2.900971,2.6042364,2.3075018,2.0107672,1.7140326,5.899552,10.081166,14.2666855,18.452206,22.637724,18.237463,13.837202,9.43694,5.036679,0.63641757,5.3451266,10.053836,14.75864,19.46735,24.17606,22.879797,21.583536,20.291178,18.994917,17.698656,15.929961,14.161267,12.388668,10.619974,8.85128,11.424281,13.993378,16.56638,19.13938,21.712381,17.48001,13.247637,9.0152645,4.7828927,0.5505207,0.44900626,0.3513962,0.24988174,0.14836729,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.6754616,1.3509232,2.0263848,2.7018464,3.3734035,2.9165885,2.4597735,2.0029583,1.5461433,1.0893283,1.261122,1.4329157,1.6047094,1.7765031,1.9482968,1.5617609,1.1713207,0.78088045,0.39044023,0.0,0.07027924,0.14055848,0.21083772,0.28111696,0.3513962,0.79649806,1.2455044,1.6906061,2.1396124,2.5886188,2.1161861,1.6437533,1.1713207,0.698888,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.339683,0.3670138,0.39434463,0.42167544,0.44900626,0.40215343,0.3553006,0.30844778,0.26159495,0.21083772,0.1756981,0.14055848,0.10932326,0.07418364,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.14836729,0.14836729,0.14836729,0.14836729,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.23035973,0.39824903,0.5661383,0.7340276,0.9019169,0.7301232,0.5583295,0.39044023,0.21864653,0.05075723,0.1639849,0.28111696,0.39434463,0.5114767,0.62470436,0.77697605,0.92924774,1.0815194,1.2337911,1.3860629,1.2025559,1.0190489,0.8316377,0.6481308,0.46071947,0.3709182,0.27721256,0.1835069,0.093705654,0.0,0.078088045,0.15617609,0.23426414,0.30844778,0.38653582,0.45681506,0.5231899,0.58956474,0.6559396,0.7262188,0.6910792,0.659844,0.62860876,0.59346914,0.5622339,0.61689556,0.6715572,0.7262188,0.78088045,0.8394465,0.71841,0.60127795,0.48414588,0.3670138,0.24988174,0.25378615,0.26159495,0.26549935,0.26940376,0.27330816,0.39824903,0.5231899,0.6481308,0.77307165,0.9019169,0.76916724,0.64032197,0.5114767,0.37872702,0.24988174,0.20693332,0.1639849,0.12103647,0.078088045,0.039044023,0.078088045,0.12103647,0.1639849,0.20693332,0.24988174,0.46852827,0.6832704,0.9019169,1.1205635,1.33921,1.4953861,1.6515622,1.8116426,1.9678187,2.1239948,2.7057507,3.2914112,3.873167,4.454923,5.036679,5.813655,6.5867267,7.363703,8.136774,8.913751,8.140678,7.3715115,6.602344,5.833177,5.0640097,5.8175592,6.571109,7.328563,8.082112,8.835662,9.983557,11.127546,12.271536,13.415526,14.56342,15.203742,15.847969,16.48829,17.132517,17.776743,19.248703,20.720663,22.192623,23.664581,25.136541,24.476698,23.816854,23.15701,22.497166,21.837322,22.184814,22.532305,22.879797,23.22729,23.574781,24.62116,25.663635,26.710016,27.756395,28.79887,29.201025,29.603178,30.009235,30.411388,30.813543,30.512903,30.212265,29.911625,29.610987,29.314253,0.039044023,0.08589685,0.13274968,0.1796025,0.22645533,0.27330816,0.3279698,0.37872702,0.43338865,0.48414588,0.5388075,0.48805028,0.43729305,0.38653582,0.3357786,0.28892577,0.39434463,0.5036679,0.60908675,0.71841,0.8238289,0.8316377,0.8355421,0.8394465,0.8433509,0.8511597,1.2025559,1.5539521,1.9092526,2.260649,2.612045,3.1664703,3.7208953,4.279225,4.83365,5.388075,6.79366,8.203149,9.608734,11.018223,12.423808,10.729298,9.030883,7.3324676,5.6340523,3.9356375,3.5686235,3.1977055,2.8267872,2.455869,2.0888553,1.9717231,1.8506867,1.7335546,1.6164225,1.4992905,1.9404879,2.3816853,2.8189783,3.260176,3.7013733,3.900498,4.0996222,4.298747,4.5017757,4.7009,4.3065557,3.9161155,3.521771,3.1313305,2.736986,2.541766,2.3426414,2.1435168,1.9482968,1.7491722,1.5734742,1.4016805,1.2259823,1.0502841,0.8745861,1.475864,2.0810463,2.6823244,3.2836022,3.8887846,4.513489,5.138193,5.7628975,6.387602,7.012306,6.774138,6.532065,6.2938967,6.0518236,5.813655,5.376362,4.942973,4.50568,4.0722914,3.638903,3.7638438,3.8887846,4.0137253,4.138666,4.263607,3.9551594,3.6467118,3.338264,3.0337205,2.7252727,3.5608149,4.4002614,5.2358036,6.0752497,6.910792,6.168956,5.4271193,4.6852827,3.9434462,3.2016098,2.7408905,2.280171,1.8194515,1.358732,0.9019169,0.8511597,0.80040246,0.74964523,0.698888,0.6481308,1.6906061,2.7330816,3.7794614,4.8219366,5.8644123,6.6843367,7.504261,8.324185,9.14411,9.964035,11.018223,12.076316,13.134409,14.192502,15.250595,16.952915,18.655233,20.357553,22.059874,23.762192,25.491842,27.221493,28.951143,30.680794,32.41435,29.439194,26.467943,23.496693,20.521538,17.550287,20.693333,23.836376,26.97942,30.118559,33.261604,35.13962,37.01764,38.895657,40.773674,42.65169,39.30562,35.959545,32.613472,29.271303,25.925232,24.464985,23.004738,21.54449,20.084246,18.623999,17.901684,17.17937,16.457056,15.734741,15.012426,15.238882,15.461433,15.687888,15.914344,16.136894,17.679134,19.221373,20.76361,22.305851,23.84809,20.31851,16.785025,13.251541,9.718058,6.1884775,10.48332,14.782067,19.080814,23.375656,27.674404,24.289286,20.900265,17.511244,14.126127,10.737106,15.371632,20.006157,24.644587,29.279112,33.91364,32.023907,30.134176,28.244446,26.350811,24.46108,24.78124,25.101402,25.421562,25.741724,26.061886,21.43517,16.808453,12.181735,7.551114,2.9243972,6.165051,9.405705,12.6463585,15.8870125,19.123762,30.907248,42.690735,54.47422,66.2538,78.037285,66.445114,54.852947,43.260777,31.668606,20.076437,18.42878,16.78112,15.133463,13.4858055,11.838148,9.928895,8.015738,6.1064854,4.1972322,2.2879796,6.949836,11.611692,16.273548,20.93931,25.601166,22.83685,20.076437,17.31212,14.551707,11.787391,13.532659,15.277926,17.023193,18.768461,20.51373,17.421442,14.329156,11.23687,8.140678,5.0483923,7.5276875,10.003078,12.482374,14.96167,17.437061,16.796738,16.152512,15.5082855,14.867964,14.223738,18.393639,22.563541,26.733442,30.903343,35.073246,31.203983,27.330816,23.45765,19.584482,15.711315,15.215456,14.7156925,14.219833,13.723974,13.224211,14.251068,15.274021,16.300879,17.323833,18.35069,15.601992,12.853292,10.108498,7.3597984,4.6110992,8.062591,11.514082,14.96167,18.41316,21.860748,20.99397,20.127193,19.260416,18.393639,17.526861,14.321347,11.115833,7.910319,4.704805,1.4992905,3.631094,5.7668023,7.898606,10.03041,12.162213,10.963562,9.761005,8.562354,7.363703,6.1611466,5.462259,4.7633705,4.0605783,3.3616903,2.6628022,2.5378613,2.4129205,2.2879796,2.1630387,2.0380979,3.3929255,4.747753,6.1025805,7.4574084,8.812236,12.47847,16.140799,19.807034,23.473267,27.135595,22.602585,18.069574,13.532659,8.995743,4.462732,3.638903,2.8111696,1.9873407,1.1635119,0.3357786,1.097137,1.8584955,2.6159496,3.377308,4.138666,3.9668727,3.7989833,3.6271896,3.4593005,3.2875066,2.9439192,2.6042364,2.260649,1.9170616,1.5734742,6.8561306,12.134882,17.413633,22.696291,27.975042,22.547922,17.124708,11.701493,6.2743745,0.8511597,3.260176,5.6691923,8.078208,10.491129,12.900145,14.625891,16.355541,18.081287,19.810938,21.536682,18.61619,15.6917925,12.771299,9.846903,6.9264097,11.018223,15.110037,19.20185,23.293663,27.389381,22.052063,16.71865,11.381332,6.0479193,0.7106012,0.57394713,0.43729305,0.30063897,0.1639849,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.46071947,0.92534333,1.3860629,1.8506867,2.3114061,2.1396124,1.9678187,1.796025,1.6242313,1.4485333,1.678893,1.9092526,2.1396124,2.3699722,2.6003318,2.0810463,1.5617609,1.038571,0.5192855,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.40605783,0.63641757,0.8667773,1.0932326,1.3235924,1.1205635,0.9136301,0.7106012,0.5036679,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.3435874,0.31625658,0.28502136,0.25378615,0.22645533,0.20693332,0.19131571,0.1717937,0.15617609,0.13665408,0.12103647,0.10151446,0.08589685,0.06637484,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.23816854,0.41777104,0.59346914,0.77307165,0.94876975,0.76526284,0.58175594,0.39434463,0.21083772,0.023426414,0.12103647,0.21474212,0.30844778,0.40605783,0.4997635,0.6832704,0.8667773,1.0463798,1.2298868,1.4133936,1.2455044,1.077615,0.9097257,0.7418364,0.57394713,0.46071947,0.3435874,0.23035973,0.113227665,0.0,0.058566034,0.113227665,0.1717937,0.23035973,0.28892577,0.39044023,0.49195468,0.59346914,0.698888,0.80040246,0.76526284,0.7301232,0.6949836,0.659844,0.62470436,0.679366,0.7301232,0.78088045,0.8355421,0.8862993,0.76135844,0.63251317,0.5036679,0.37872702,0.24988174,0.26549935,0.28111696,0.29673457,0.30844778,0.3240654,0.47633708,0.62470436,0.77307165,0.92534333,1.0737107,0.92143893,0.76916724,0.61689556,0.46462387,0.31235218,0.26159495,0.20693332,0.15617609,0.10151446,0.05075723,0.078088045,0.10541886,0.13274968,0.16008049,0.18741131,0.339683,0.49195468,0.6442264,0.79649806,0.94876975,1.0737107,1.1947471,1.3157835,1.4407244,1.5617609,1.8975395,2.233318,2.5690966,2.900971,3.2367494,4.5017757,5.7628975,7.0240197,8.289046,9.550168,8.628729,7.703386,6.7819467,5.860508,4.939069,5.801942,6.6687193,7.531592,8.398369,9.261242,10.522364,11.783486,13.040704,14.301826,15.562947,15.863586,16.168129,16.46877,16.773312,17.073952,17.815788,18.56153,19.303364,20.0452,20.787037,20.40831,20.025679,19.646952,19.268225,18.885593,19.756275,20.623053,21.48983,22.356607,23.223385,24.734388,26.245392,27.756395,29.263494,30.774498,31.332829,31.891157,32.449486,33.003914,33.56224,32.925823,32.289406,31.649084,31.012667,30.37625,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.24988174,0.31235218,0.37482262,0.43729305,0.4997635,0.43729305,0.37482262,0.31235218,0.24988174,0.18741131,0.28892577,0.38653582,0.48805028,0.58566034,0.6871748,0.7106012,0.737932,0.76135844,0.78868926,0.81211567,1.261122,1.7140326,2.1630387,2.612045,3.0610514,3.0610514,3.0610514,3.0610514,3.0610514,3.0610514,5.1889505,7.3129454,9.43694,11.560935,13.688834,11.736633,9.788337,7.8361354,5.8878384,3.9356375,3.5491016,3.1625657,2.77603,2.3855898,1.999054,1.8741131,1.7491722,1.6242313,1.4992905,1.3743496,1.8233559,2.2762666,2.7252727,3.174279,3.6232853,3.6232853,3.6232853,3.6232853,3.6232853,3.6232853,3.2992198,2.9751544,2.6510892,2.3231194,1.999054,1.9482968,1.901444,1.8506867,1.7999294,1.7491722,1.5617609,1.3743496,1.1869383,0.999527,0.81211567,1.5890918,2.3621633,3.1391394,3.912211,4.689187,5.22409,5.7628975,6.3017054,6.8366084,7.375416,7.0747766,6.774138,6.473499,6.1767645,5.8761253,5.4388323,5.001539,4.564246,4.123049,3.6857557,3.775557,3.8614538,3.951255,4.037152,4.123049,3.7638438,3.4007344,3.0376248,2.6745155,2.3114061,3.474918,4.6384296,5.801942,6.9615493,8.125061,7.1880045,6.250948,5.3138914,4.376835,3.435874,2.8619268,2.2879796,1.7140326,1.1361811,0.5622339,0.5505207,0.5388075,0.5231899,0.5114767,0.4997635,1.8389735,3.174279,4.513489,5.8487945,7.1880045,8.039165,8.886419,9.737579,10.588739,11.435994,12.712734,13.985569,15.262308,16.539047,17.811884,19.451733,21.087677,22.723621,24.36347,25.999414,28.51385,31.02438,33.538815,36.049347,38.56378,35.100574,31.637371,28.174168,24.710962,21.251661,24.761719,28.27568,31.785738,35.2997,38.813663,40.199726,41.58579,42.975754,44.36182,45.751785,40.875187,35.99859,31.125895,26.249296,21.376602,20.548868,5052.0,18.90121,18.073479,17.24965,16.539047,15.824542,15.113941,14.399435,13.688834,13.599033,13.513136,13.423335,13.337439,13.251541,14.364296,15.473146,16.585901,17.698656,18.81141,15.613705,12.412095,9.2104845,6.012779,2.8111696,8.136774,13.462379,18.787983,24.113588,29.439194,25.085785,20.73628,16.386776,12.037272,7.687768,14.11051,20.537155,26.963802,33.386543,39.81319,37.423695,35.038105,32.648613,30.263021,27.873528,28.712975,29.548515,30.387962,31.223505,32.06295,26.237583,20.412214,14.586847,8.761478,2.9361105,7.098203,11.2642,15.426293,19.588387,23.750479,38.41151,53.076443,67.73747,82.398506,97.06344,80.81332,64.563194,48.313072,32.06295,15.812829,15.586374,15.363823,15.137367,14.9109125,14.688361,12.212971,9.737579,7.262188,4.786797,2.3114061,8.011833,13.712261,19.412687,25.113115,30.813543,26.475752,22.13796,17.800169,13.462379,9.124588,12.201257,15.274021,18.35069,21.423454,24.500124,20.599627,16.69913,12.798631,8.898132,5.001539,7.1489606,9.300286,11.4516115,13.599033,15.750359,14.575133,13.399908,12.224684,11.0494585,9.874233,15.723028,21.575727,27.424522,33.273315,39.126015,34.62424,30.126368,25.624592,21.12672,16.624945,16.023666,15.426293,14.825015,14.223738,13.626364,15.063184,16.500004,17.936825,19.373644,20.81437,17.464392,14.114414,10.760532,7.4105554,4.0605783,8.312472,12.560462,16.812357,21.06425,25.31224,24.625065,23.937891,23.250715,22.563541,21.876366,17.49953,13.1266,8.749765,4.376835,0.0,2.77603,5.548156,8.324185,11.100216,13.8762455,12.373051,10.87376,9.37447,7.8751793,6.375889,5.688714,5.001539,4.3143644,3.6232853,2.9361105,2.5769055,2.2137961,1.8506867,1.4875772,1.1244678,3.076669,5.024966,6.9732623,8.925464,10.87376,14.411149,17.948538,21.485926,25.023314,28.560703,23.898846,19.23699,14.575133,9.913278,5.251421,4.21285,3.174279,2.135708,1.1010414,0.062470436,0.999527,1.9365835,2.87364,3.8106966,4.7516575,4.474445,4.2011366,3.9239242,3.6506162,3.3734035,2.9868677,2.6003318,2.2137961,1.8233559,1.43682,7.812709,14.188598,20.564487,26.936472,33.31236,26.862288,20.412214,13.962143,7.5120697,1.0619974,1.175225,1.2884527,1.4016805,1.5110037,1.6242313,6.375889,11.123642,15.875299,20.626957,25.37471,21.298513,17.226223,13.150026,9.073831,5.001539,10.612165,16.226696,21.837322,27.451853,33.062477,26.624119,20.18576,13.751305,7.3129454,0.8745861,0.698888,0.5231899,0.3513962,0.1756981,0.0,0.0,0.0,0.0,0.0,0.0,0.24988174,0.4997635,0.74964523,0.999527,1.2494087,1.3626363,1.475864,1.5890918,1.698415,1.8116426,2.1005683,2.3855898,2.6745155,2.9634414,3.2484627,2.6003318,1.9482968,1.3001659,0.6481308,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.3513962,0.26159495,0.1756981,0.08589685,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.24988174,0.43729305,0.62470436,0.81211567,0.999527,0.80040246,0.60127795,0.39824903,0.19912452,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.58566034,0.80040246,1.0112402,1.2259823,1.43682,1.2884527,1.1361811,0.9878138,0.8394465,0.6871748,0.5505207,0.41386664,0.27330816,0.13665408,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.3240654,0.46071947,0.60127795,0.737932,0.8745861,0.8394465,0.80040246,0.76135844,0.7262188,0.6871748,0.737932,0.78868926,0.8394465,0.8862993,0.93705654,0.80040246,0.6637484,0.5231899,0.38653582,0.24988174,0.27330816,0.30063897,0.3240654,0.3513962,0.37482262,0.5505207,0.7262188,0.9019169,1.0737107,1.2494087,1.0737107,0.9019169,0.7262188,0.5505207,0.37482262,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.21083772,0.30063897,0.38653582,0.47633708,0.5622339,0.6481308,0.737932,0.8238289,0.9136301,0.999527,1.0893283,1.175225,1.261122,1.3509232,1.43682,3.1859922,4.939069,6.688241,8.437413,10.186585,9.112875,8.039165,6.9615493,5.8878384,4.814128,5.786324,6.7624245,7.7385254,8.710721,9.686822,11.061172,12.439425,13.813775,15.188125,16.562475,16.52343,16.48829,16.449247,16.414106,16.375063,16.386776,16.398489,16.414106,16.42582,16.437534,16.33602,16.238409,16.136894,16.039284,15.93777,17.323833,18.7138,20.099863,21.485926,22.875893,24.85152,26.827148,28.79887,30.774498,32.750126,33.460728,34.175232,34.885834,35.600338,36.31094,35.338745,34.362644,33.386543,32.41435,31.438248,0.0,0.031235218,0.06637484,0.09761006,0.12884527,0.1639849,0.21083772,0.26159495,0.31235218,0.3631094,0.41386664,0.3631094,0.31235218,0.26159495,0.21083772,0.1639849,0.24597734,0.3279698,0.40996224,0.49195468,0.57394713,0.60908675,0.6442264,0.679366,0.7145056,0.74964523,1.2533131,1.7608855,2.2645533,2.7682211,3.2757936,3.4124475,3.5491016,3.6857557,3.8263142,3.9629683,5.5091114,7.0513506,8.597494,10.143637,11.685876,10.03041,8.371038,6.715572,5.056201,3.4007344,3.0805733,2.7643168,2.4480603,2.1318035,1.8116426,1.6906061,1.5734742,1.4524376,1.3314011,1.2142692,1.5969005,1.9756275,2.358259,2.7408905,3.1235218,3.2094188,3.2914112,3.3734035,3.455396,3.5373883,3.2289407,2.9165885,2.6081407,2.2957885,1.9873407,2.0380979,2.0927596,2.1435168,2.1981785,2.2489357,2.1513257,2.0498111,1.9482968,1.8506867,1.7491722,2.436347,3.1235218,3.8106966,4.5017757,5.1889505,5.700427,6.211904,6.7233806,7.238762,7.7502384,7.367607,6.984976,6.602344,6.2197127,5.8370814,5.4427366,5.0483923,4.6540475,4.2557983,3.8614538,3.9356375,4.0137253,4.087909,4.1620927,4.2362766,4.1581883,4.0761957,3.998108,3.9161155,3.8380275,4.892216,5.9464045,7.000593,8.058686,9.112875,8.335898,7.562827,6.785851,6.012779,5.2358036,4.548629,3.8614538,3.174279,2.4871042,1.7999294,1.7765031,1.7491722,1.7257458,1.698415,1.6749885,2.9634414,4.251894,5.5364423,6.824895,8.113348,8.827853,9.542359,10.256865,10.971371,11.685876,12.6463585,13.606842,14.567325,15.527808,16.48829,17.886066,19.283842,20.68162,22.079395,23.473267,26.284435,29.095606,31.906775,34.71404,37.52521,34.151806,30.774498,27.401094,24.023787,20.650383,23.711435,26.768581,29.829634,32.890686,35.951736,37.263615,38.5794,39.895184,41.210964,42.52675,39.446175,36.365604,33.28503,30.204456,27.123882,26.28053,25.433277,24.589926,23.746574,22.899319,21.411741,19.92026,18.42878,16.941202,15.449719,15.387249,15.324779,15.262308,15.199838,15.137367,15.816733,16.492195,17.17156,17.847023,18.526388,15.274021,12.025558,8.773191,5.5247293,2.2762666,6.5359693,10.799577,15.063184,19.326792,23.586494,20.435642,17.280884,14.130032,10.979179,7.824422,13.954333,20.084246,26.214157,32.344067,38.47398,37.326084,36.174286,35.026394,33.874596,32.7267,33.386543,34.046387,34.70623,35.366077,36.02592,29.46262,22.899319,16.33602,9.776623,3.213323,6.6687193,10.124115,13.579511,17.031002,20.486399,32.06295,43.6356,55.21215,66.788704,78.36135,66.21866,54.072067,41.925472,29.78278,17.636185,18.042242,18.448301,18.854359,19.256512,19.662569,16.117373,12.572175,9.026978,5.481781,1.9365835,8.8083315,15.676175,22.547922,29.415766,36.287514,31.820879,27.354242,22.883701,18.417065,13.950429,15.9221525,17.893875,19.865599,21.841227,23.81295,20.267752,16.722555,13.177358,9.63216,6.086963,8.484266,10.881569,13.2788725,15.676175,18.073479,16.976341,15.879204,14.782067,13.68493,12.587793,17.804073,23.01645,28.232733,33.449013,38.661392,34.628143,30.590992,26.557745,22.520592,18.487345,17.909492,17.331642,16.75379,16.175938,15.598087,15.945579,16.289165,16.636658,16.980246,17.323833,15.195933,13.0719385,10.944039,8.81614,6.688241,9.460366,12.232492,15.004618,17.776743,20.548868,19.971018,19.389261,18.81141,18.229654,17.651802,15.016331,12.384764,9.753197,7.1216297,4.4861584,6.211904,7.9376497,9.663396,11.389141,13.110983,11.791295,10.467703,9.14411,7.824422,6.5008297,5.8487945,5.196759,4.5408196,3.8887846,3.2367494,2.8345962,2.4324427,2.0302892,1.6281357,1.2259823,3.018103,4.8102236,6.602344,8.3944645,10.186585,13.431144,16.671797,19.916355,23.15701,26.401567,22.20824,18.014912,13.821584,9.628256,5.4388323,4.365122,3.2914112,2.2216048,1.1478943,0.07418364,0.96438736,1.8545911,2.7447948,3.6349986,4.5252023,4.2479897,3.970777,3.6935644,3.416352,3.1391394,2.7526035,2.366068,1.9834363,1.5969005,1.2142692,6.3407493,11.46723,16.59371,21.724094,26.850574,21.763138,16.679607,11.596075,6.5086384,1.4251068,1.6242313,1.8194515,2.018576,2.2137961,2.4129205,6.2938967,10.178777,14.059752,17.94073,21.82561,18.268698,14.711788,11.150972,7.5940623,4.037152,8.519405,13.001659,17.483913,21.966167,26.448421,21.298513,16.148607,10.998701,5.8487945,0.698888,0.61689556,0.5309987,0.44510186,0.359205,0.27330816,0.21864653,0.1639849,0.10932326,0.05466163,0.0,0.19912452,0.39824903,0.60127795,0.80040246,0.999527,1.1361811,1.2767396,1.4133936,1.5500476,1.6867018,2.0615244,2.436347,2.8111696,3.1859922,3.5608149,2.854118,2.1474214,1.4407244,0.7340276,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.07027924,0.14055848,0.21083772,0.28111696,0.3513962,0.28111696,0.21083772,0.14055848,0.07027924,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.12494087,0.19912452,0.27330816,0.3513962,0.42557985,0.339683,0.25378615,0.1717937,0.08589685,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.24207294,0.43338865,0.62860876,0.8199245,1.0112402,0.8238289,0.63641757,0.44900626,0.26159495,0.07418364,0.12103647,0.1717937,0.21864653,0.26549935,0.31235218,0.48414588,0.6520352,0.8238289,0.9917182,1.1635119,1.0463798,0.92924774,0.80821127,0.6910792,0.57394713,0.46462387,0.3553006,0.24597734,0.13665408,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.28111696,0.41386664,0.5466163,0.679366,0.81211567,0.78088045,0.75354964,0.7223144,0.6910792,0.6637484,0.7066968,0.75354964,0.79649806,0.8433509,0.8862993,0.79649806,0.7027924,0.60908675,0.5192855,0.42557985,0.4958591,0.5700427,0.6442264,0.7145056,0.78868926,0.98390937,1.183034,1.3782539,1.5773785,1.7765031,1.5227169,1.2689307,1.0190489,0.76526284,0.5114767,0.46071947,0.41386664,0.3631094,0.31235218,0.26159495,0.29673457,0.3318742,0.3670138,0.40215343,0.43729305,0.44900626,0.45681506,0.46852827,0.47633708,0.48805028,0.5583295,0.62860876,0.698888,0.76916724,0.8394465,0.92924774,1.0229534,1.116659,1.2064602,1.3001659,2.7213683,4.1464753,5.5676775,6.98888,8.413987,7.578445,6.746807,5.9151692,5.083532,4.251894,5.087436,5.9268827,6.7624245,7.601871,8.437413,9.526741,10.612165,11.701493,12.786918,13.8762455,13.950429,14.024612,14.098797,14.176885,14.251068,14.668839,15.086611,15.504381,15.918248,16.33602,16.48829,16.636658,16.788929,16.937298,17.085665,18.276506,19.463446,20.650383,21.837322,23.02426,24.710962,26.393759,28.080462,29.763258,31.44996,32.359688,33.269413,34.17914,35.088863,35.99859,34.760895,33.519295,32.281597,31.039997,29.798397,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.1756981,0.21083772,0.24988174,0.28892577,0.3240654,0.28892577,0.24988174,0.21083772,0.1756981,0.13665408,0.20302892,0.26940376,0.3318742,0.39824903,0.46071947,0.5075723,0.5544251,0.59737355,0.6442264,0.6871748,1.2494087,1.8077383,2.366068,2.9283018,3.4866312,3.7638438,4.037152,4.3143644,4.5876727,4.860981,5.8292727,6.79366,7.758047,8.722435,9.686822,8.324185,6.957645,5.591104,4.2284675,2.8619268,2.6159496,2.366068,2.1200905,1.8741131,1.6242313,1.5110037,1.3938715,1.2806439,1.1635119,1.0502841,1.3665408,1.678893,1.9951496,2.3114061,2.6237583,2.7916477,2.9556324,3.1196175,3.2836022,3.4514916,3.154757,2.8619268,2.5651922,2.2684577,1.9756275,2.1318035,2.2840753,2.4402514,2.5964274,2.7486992,2.736986,2.7252727,2.7135596,2.7018464,2.6862288,3.2875066,3.8887846,4.4861584,5.087436,5.688714,6.1767645,6.66091,7.1489606,7.6370106,8.125061,7.660437,7.195813,6.7311897,6.266566,5.801942,5.446641,5.095245,4.743849,4.388548,4.037152,4.0996222,4.1620927,4.224563,4.2870336,4.349504,4.552533,4.755562,4.958591,5.1616197,5.3607445,6.309514,7.2582836,8.203149,9.151918,10.100689,9.487698,8.874706,8.261715,7.648724,7.0357327,6.239235,5.4388323,4.6384296,3.8380275,3.0376248,2.998581,2.9634414,2.9243972,2.8892577,2.8502135,4.087909,5.3256044,6.5633,7.800996,9.0386915,9.616543,10.198298,10.77615,11.357906,11.935758,12.583888,13.228115,13.872341,14.516567,15.160794,16.320402,17.476105,18.635712,19.791414,20.951023,24.058928,27.16683,30.27083,33.378735,36.48664,33.19913,29.911625,26.624119,23.336613,20.049105,22.657246,25.265387,27.873528,30.481668,33.085903,34.33141,35.57301,36.81461,38.05621,39.301712,38.01326,36.72871,35.444164,34.159615,32.87507,32.00829,31.145416,30.278639,29.415766,28.548988,26.284435,24.015978,21.74752,19.479063,17.210606,17.175465,17.136421,17.101282,17.062239,17.023193,17.26917,17.511244,17.753317,17.99539,18.237463,14.938243,11.639023,8.335898,5.036679,1.737459,4.939069,8.136774,11.338385,14.53609,17.7377,15.781594,13.829392,11.873287,9.917182,7.9610763,13.798158,19.631334,25.468416,31.301594,37.138676,37.22457,37.314373,37.40027,37.486168,37.575966,38.05621,38.540356,39.0245,39.50474,39.988888,32.687656,25.386423,18.089096,10.787864,3.4866312,6.2353306,8.98403,11.728825,14.477524,17.226223,25.71049,34.198658,42.68683,51.175,59.66317,51.62401,43.580936,35.541775,27.50261,19.463446,20.498112,21.532778,22.567446,23.602112,24.636778,20.021774,15.406772,10.791768,6.1767645,1.5617609,9.600925,17.643993,25.683159,33.72232,41.761486,37.166004,32.56662,27.971138,23.371752,18.77627,19.646952,20.51373,21.38441,22.255093,23.125774,19.935879,16.745981,13.556085,10.366188,7.1762915,9.8195715,12.466757,15.110037,17.753317,20.400501,19.381453,18.3585,17.33945,16.320402,15.3013525,19.881216,24.46108,29.040943,33.620808,38.200672,34.628143,31.05952,27.490896,23.918367,20.349745,19.795319,19.240894,18.68647,18.12814,17.573715,16.827974,16.07833,15.332587,14.586847,13.837202,12.93138,12.029464,11.123642,10.217821,9.311999,10.608261,11.900618,13.196879,14.493141,15.789403,15.313066,14.840633,14.3682,13.895767,13.423335,12.533132,11.6468315,10.756628,9.866425,8.976221,9.651682,10.323239,10.998701,11.674163,12.349625,11.205634,10.061645,8.913751,7.7697606,6.6257706,6.008875,5.388075,4.7711797,4.154284,3.5373883,3.096191,2.6510892,2.2098918,1.7686942,1.3235924,2.959537,4.5954814,6.2314262,7.8634663,9.499411,12.447234,15.395058,18.342882,21.290705,24.23853,20.51373,16.792833,13.068034,9.347139,5.6262436,4.5173936,3.408543,2.3035975,1.1947471,0.08589685,0.92924774,1.7725986,2.6159496,3.4593005,4.298747,4.0215344,3.7404175,3.4593005,3.1781836,2.900971,2.5183394,2.135708,1.7530766,1.3704453,0.9878138,4.8687897,8.745861,12.626837,16.507812,20.388788,16.667892,12.946998,9.226103,5.5091114,1.7882162,2.069333,2.3543546,2.6354716,2.9165885,3.2016098,6.2158084,9.230007,12.244205,15.258404,18.276506,15.234978,12.193448,9.155824,6.114294,3.076669,6.426646,9.780528,13.134409,16.484386,19.838268,15.97291,12.111456,8.250002,4.388548,0.5231899,0.5309987,0.5349031,0.5388075,0.5466163,0.5505207,0.44119745,0.3318742,0.21864653,0.10932326,0.0,0.14836729,0.30063897,0.44900626,0.60127795,0.74964523,0.9136301,1.0737107,1.2376955,1.4016805,1.5617609,2.0263848,2.4871042,2.951728,3.4124475,3.873167,3.1118085,2.3465457,1.5812829,0.8160201,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.05075723,0.10541886,0.15617609,0.21083772,0.26159495,0.21083772,0.15617609,0.10541886,0.05075723,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.18741131,0.3357786,0.48805028,0.63641757,0.78868926,0.62860876,0.47243267,0.31625658,0.15617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.23426414,0.43338865,0.62860876,0.8277333,1.0268579,0.8511597,0.6754616,0.4997635,0.3240654,0.14836729,0.1717937,0.19131571,0.21083772,0.23035973,0.24988174,0.37872702,0.5036679,0.63251317,0.76135844,0.8862993,0.80430686,0.71841,0.63251317,0.5466163,0.46071947,0.37872702,0.29673457,0.21474212,0.13274968,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.23816854,0.3670138,0.4958591,0.62079996,0.74964523,0.7262188,0.7066968,0.6832704,0.659844,0.63641757,0.679366,0.71841,0.75745404,0.79649806,0.8394465,0.78868926,0.7418364,0.6949836,0.6481308,0.60127795,0.71841,0.8394465,0.96048295,1.0815194,1.1986516,1.4212024,1.639849,1.8584955,2.0810463,2.2996929,1.9717231,1.639849,1.3118792,0.98000497,0.6481308,0.61299115,0.57394713,0.5388075,0.4997635,0.46071947,0.5192855,0.57785153,0.63641757,0.6910792,0.74964523,0.6832704,0.61689556,0.5466163,0.48024148,0.41386664,0.46462387,0.5192855,0.5700427,0.62079996,0.6754616,0.77307165,0.8706817,0.96829176,1.0659018,1.1635119,2.2567444,3.3538816,4.447114,5.5442514,6.6374836,6.0479193,5.4583545,4.8687897,4.279225,3.6857557,4.388548,5.087436,5.786324,6.4891167,7.1880045,7.988407,8.78881,9.589212,10.38571,11.186112,11.373524,11.560935,11.748346,11.935758,12.123169,12.946998,13.770826,14.590752,15.41458,16.238409,16.636658,17.03881,17.437061,17.839214,18.237463,19.225277,20.21309,21.200905,22.188719,23.176533,24.570404,25.964275,27.358147,28.755922,30.149794,31.258644,32.36359,33.47244,34.58129,35.686237,34.18304,32.67594,31.172749,29.665648,28.162453,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.13665408,0.1639849,0.18741131,0.21083772,0.23816854,0.21083772,0.18741131,0.1639849,0.13665408,0.113227665,0.16008049,0.20693332,0.25378615,0.30063897,0.3513962,0.40605783,0.46071947,0.5153811,0.5700427,0.62470436,1.2415999,1.8545911,2.4714866,3.084478,3.7013733,4.1113358,4.5252023,4.939069,5.349031,5.7628975,6.1494336,6.532065,6.918601,7.3012323,7.687768,6.6140575,5.5442514,4.4705405,3.39683,2.3231194,2.1474214,1.9717231,1.7921207,1.6164225,1.43682,1.3274968,1.2181735,1.1088502,0.9956226,0.8862993,1.1361811,1.3821584,1.6281357,1.8780174,2.1239948,2.3738766,2.619854,2.8658314,3.1157131,3.3616903,3.0805733,2.803361,2.522244,2.241127,1.9639144,2.2216048,2.4792955,2.7330816,2.9907722,3.2484627,3.3265507,3.4007344,3.474918,3.5491016,3.6232853,4.138666,4.650143,5.1616197,5.6730967,6.1884775,6.649197,7.113821,7.57454,8.039165,8.499884,7.9532676,7.406651,6.8561306,6.309514,5.7628975,5.45445,5.142098,4.83365,4.521298,4.21285,4.263607,4.3143644,4.3612175,4.4119744,4.462732,4.9468775,5.4310236,5.919074,6.4032197,6.8873653,7.726812,8.566258,9.405705,10.249056,11.088503,10.6355915,10.186585,9.737579,9.288573,8.835662,7.9259367,7.012306,6.098676,5.1889505,4.2753205,4.224563,4.173806,4.126953,4.0761957,4.025439,5.212377,6.3993154,7.5862536,8.773191,9.964035,10.409137,10.8542385,11.29934,11.744442,12.185639,12.517513,12.849388,13.177358,13.509232,13.837202,14.754736,15.672271,16.589806,17.50734,18.424873,21.829514,25.234152,28.63879,32.04343,35.448067,32.250362,29.048752,25.851048,22.649437,19.451733,21.603058,23.758287,25.913517,28.068748,30.223978,31.395298,32.56662,33.734035,34.905357,36.076675,36.584248,37.095726,37.6033,38.114777,38.62625,37.739952,36.853653,35.971256,35.084957,34.198658,31.15713,28.111696,25.066263,22.020828,18.975395,18.963682,18.95197,18.936352,18.924637,18.912924,18.72161,18.526388,18.335073,18.143757,17.948538,14.59856,11.248583,7.898606,4.548629,1.1986516,3.338264,5.473972,7.6135845,9.749292,11.888905,11.131451,10.373997,9.616543,8.859089,8.101635,13.638077,19.178425,24.718771,30.259117,35.799465,37.12306,38.450554,39.774147,41.101643,42.425236,42.72978,43.03432,43.338863,43.64341,43.951855,35.912693,27.873528,19.838268,11.799104,3.7638438,5.801942,7.843944,9.882042,11.924045,13.962143,19.36193,24.761719,30.161507,35.561295,40.961082,37.025448,33.09371,29.158075,25.222439,21.2868,22.953981,24.617256,26.284435,27.947712,29.610987,23.926178,18.241367,12.556558,6.871748,1.1869383,10.397423,19.607908,28.818394,38.028877,47.239365,42.51113,37.7829,33.05467,28.326439,23.598207,23.367847,23.133583,22.903223,22.668959,22.4386,19.604004,16.769407,13.930907,11.096312,8.261715,11.154878,14.048039,16.941202,19.834364,22.723621,21.78266,20.8417,19.896833,18.955873,18.011007,21.958359,25.901804,29.849155,33.792603,37.73605,34.63205,31.528048,28.42405,25.316145,22.212145,21.681147,21.146242,20.615244,20.084246,19.549341,17.71037,15.871395,14.028518,12.189544,10.350571,10.666827,10.983084,11.303245,11.619501,11.935758,11.756155,11.572648,11.389141,11.205634,11.0260315,10.6590185,10.295909,9.928895,9.565785,9.198771,10.053836,10.904996,11.756155,12.611219,13.462379,13.087557,12.712734,12.337912,11.963089,11.588266,10.619974,9.651682,8.683391,7.719003,6.7507114,6.168956,5.5832953,5.001539,4.4197836,3.8380275,3.3538816,2.87364,2.3894942,1.9092526,1.4251068,2.900971,4.380739,5.8566036,7.336372,8.812236,11.4633255,14.118319,16.769407,19.4244,22.07549,18.823124,15.570756,12.318389,9.066022,5.813655,4.6696653,3.5256753,2.3855898,1.2415999,0.10151446,0.8941081,1.6906061,2.4831998,3.279698,4.0761957,3.7911747,3.5100577,3.2289407,2.9439192,2.6628022,2.2840753,1.901444,1.5227169,1.1439898,0.76135844,3.39683,6.028397,8.659965,11.291532,13.923099,11.568744,9.21439,6.860035,4.50568,2.1513257,2.5183394,2.8853533,3.252367,3.619381,3.9863946,6.133816,8.281238,10.4286585,12.576079,14.723501,12.201257,9.679013,7.1567693,4.6345253,2.1122816,4.3338866,6.5554914,8.781001,11.002605,13.224211,10.651209,8.074304,5.5013027,2.9243972,0.3513962,0.44510186,0.5388075,0.63641757,0.7301232,0.8238289,0.659844,0.4958591,0.3318742,0.1639849,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.6871748,0.8745861,1.0619974,1.2494087,1.43682,1.9873407,2.5378613,3.0883822,3.638903,4.1894236,3.3655949,2.541766,1.7218413,0.8980125,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.24988174,0.47633708,0.698888,0.92534333,1.1517987,0.92143893,0.6910792,0.46071947,0.23035973,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.22645533,0.42948425,0.63251317,0.8355421,1.038571,0.8745861,0.7106012,0.5505207,0.38653582,0.22645533,0.21864653,0.21083772,0.20302892,0.19522011,0.18741131,0.27330816,0.359205,0.44119745,0.5270943,0.61299115,0.5583295,0.5075723,0.45681506,0.40215343,0.3513962,0.29673457,0.23816854,0.1835069,0.12884527,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.19912452,0.32016098,0.44119745,0.5661383,0.6871748,0.6715572,0.6559396,0.6442264,0.62860876,0.61299115,0.6481308,0.6832704,0.71841,0.75354964,0.78868926,0.78478485,0.78088045,0.78088045,0.77697605,0.77307165,0.94096094,1.1088502,1.2767396,1.4446288,1.6125181,1.8545911,2.096664,2.338737,2.5808098,2.8267872,2.416825,2.0107672,1.6008049,1.1947471,0.78868926,0.76135844,0.737932,0.7106012,0.6871748,0.6637484,0.7418364,0.8238289,0.9019169,0.98390937,1.0619974,0.91753453,0.77307165,0.62860876,0.48414588,0.3357786,0.3709182,0.40605783,0.44119745,0.47633708,0.5114767,0.61689556,0.71841,0.8199245,0.92143893,1.0268579,1.7921207,2.5612879,3.3265507,4.095718,4.860981,4.513489,4.165997,3.8185053,3.4710135,3.1235218,3.6857557,4.251894,4.814128,5.376362,5.938596,6.4500723,6.9615493,7.473026,7.988407,8.499884,8.800523,9.101162,9.4018,9.698535,9.999174,11.229061,12.455043,13.6810255,14.9109125,16.136894,16.788929,17.437061,18.089096,18.737226,19.389261,20.174046,20.962736,21.751425,22.53621,23.3249,24.429846,25.53479,26.639736,27.744682,28.849628,30.153698,31.461674,32.765743,34.069813,35.373886,33.60519,31.836496,30.063898,28.295202,26.526508,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.10151446,0.113227665,0.12494087,0.13665408,0.14836729,0.13665408,0.12494087,0.113227665,0.10151446,0.08589685,0.11713207,0.14836729,0.1756981,0.20693332,0.23816854,0.30063897,0.3670138,0.43338865,0.4958591,0.5622339,1.2337911,1.901444,2.5730011,3.240654,3.912211,4.462732,5.0132523,5.563773,6.114294,6.66091,6.46569,6.2743745,6.0791545,5.883934,5.688714,4.9078336,4.126953,3.3460727,2.5690966,1.7882162,1.678893,1.5734742,1.4641509,1.358732,1.2494087,1.1439898,1.038571,0.93315214,0.8316377,0.7262188,0.9058213,1.0854238,1.2650263,1.4446288,1.6242313,1.9561055,2.2840753,2.6159496,2.9439192,3.2757936,3.0102942,2.7447948,2.4792955,2.2137961,1.9482968,2.3114061,2.6706111,3.0298162,3.3890212,3.7482262,3.912211,4.0761957,4.2362766,4.4002614,4.564246,4.985922,5.4115014,5.8370814,6.262661,6.688241,7.125534,7.562827,8.00012,8.437413,8.874706,8.246098,7.6135845,6.984976,6.356367,5.7238536,5.4583545,5.1889505,4.9234514,4.6540475,4.388548,4.423688,4.462732,4.5017757,4.5369153,4.575959,5.3412223,6.1103897,6.8756523,7.6448197,8.413987,9.14411,9.878138,10.608261,11.342289,12.076316,11.787391,11.498465,11.213444,10.924518,10.6355915,9.612638,8.58578,7.562827,6.5359693,5.5130157,5.4505453,5.388075,5.3256044,5.263134,5.2006636,6.336845,7.47693,8.6131115,9.749292,10.889378,11.197825,11.506273,11.818625,12.127073,12.439425,12.4511385,12.466757,12.482374,12.497992,12.513609,13.189071,13.868437,14.543899,15.223265,15.8987255,19.604004,23.305378,27.00675,30.708124,34.413403,31.301594,28.18588,25.074072,21.962263,18.850454,20.552773,22.255093,23.957413,25.65973,27.362051,28.459188,29.556326,30.653461,31.750599,32.85164,35.15524,37.458836,39.76634,42.069935,44.37353,43.471615,42.565792,41.659973,40.75415,39.848328,36.02592,32.20351,28.3811,24.558691,20.73628,20.751898,20.76361,20.775324,20.787037,20.79875,20.174046,19.545437,18.916828,18.28822,17.663515,14.262781,10.862047,7.461313,4.0605783,0.6637484,1.737459,2.8111696,3.8887846,4.9624953,6.036206,6.477403,6.918601,7.355894,7.7970915,8.238289,13.481901,18.725513,23.97303,29.216642,34.464157,37.025448,39.586735,42.151928,44.713215,47.2745,47.403347,47.52829,47.657135,47.78598,47.91092,39.13773,30.364536,21.58744,12.814248,4.037152,5.368553,6.703859,8.03526,9.366661,10.698062,13.013372,15.324779,17.636185,19.951496,22.262901,22.430792,22.602585,22.770473,22.942268,23.114061,25.405945,27.701735,29.997522,32.293312,34.5891,27.834484,21.075964,14.321347,7.5667315,0.81211567,11.193921,21.571823,31.953629,42.331528,52.713333,47.85626,42.999184,38.138203,33.281124,28.42405,27.088743,25.753437,24.41813,23.086731,21.751425,19.268225,16.788929,14.309634,11.8303385,9.351044,12.490183,15.629322,18.768461,21.911505,25.050644,24.183868,23.320995,22.454218,21.591345,20.724567,24.0355,27.346434,30.653461,33.964394,37.27533,34.635952,31.996576,29.353296,26.71392,24.074545,23.566973,23.055496,22.544018,22.036446,21.52497,18.592764,15.660558,12.728352,9.796145,6.8639393,8.402273,9.940608,11.482847,13.021181,14.56342,12.90405,11.240774,9.581403,7.9220324,6.262661,6.0049706,5.74728,5.4895897,5.2318993,4.9742084,7.570636,10.163159,12.759586,15.356014,17.948538,16.52343,15.098324,13.673217,12.24811,10.826907,10.034314,9.245625,8.453031,7.6643414,6.8756523,6.329036,5.7785153,5.2318993,4.6852827,4.138666,3.6154766,3.0922866,2.5690966,2.0459068,1.5266213,2.8463092,4.165997,5.4856853,6.805373,8.125061,10.48332,12.841579,15.195933,17.554192,19.91245,17.128613,14.348679,11.564839,8.781001,6.001066,4.8219366,3.6467118,2.4675822,1.2884527,0.113227665,0.8589685,1.6086137,2.3543546,3.1039999,3.8497405,3.5647192,3.279698,2.9946766,2.7096553,2.4246337,2.0459068,1.6710842,1.2923572,0.9136301,0.5388075,1.9209659,3.3070288,4.6930914,6.0791545,7.461313,6.473499,5.481781,4.493967,3.5022488,2.514435,2.9634414,3.416352,3.8692627,4.322173,4.775084,6.055728,7.336372,8.6131115,9.893755,11.174399,9.171441,7.164578,5.1616197,3.154757,1.1517987,2.241127,3.3343596,4.4275923,5.520825,6.6140575,5.3256044,4.037152,2.7486992,1.4641509,0.1756981,0.359205,0.5466163,0.7301232,0.9136301,1.1010414,0.8784905,0.659844,0.44119745,0.21864653,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.46071947,0.6754616,0.8862993,1.1010414,1.3118792,1.9482968,2.5886188,3.2250361,3.8614538,4.5017757,3.619381,2.7408905,1.8584955,0.98000497,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.31235218,0.61299115,0.9136301,1.2142692,1.5110037,1.2103647,0.9058213,0.60518235,0.30063897,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.21864653,0.42557985,0.63641757,0.8433509,1.0502841,0.9019169,0.74964523,0.60127795,0.44900626,0.30063897,0.26549935,0.23035973,0.19522011,0.16008049,0.12494087,0.1678893,0.21083772,0.25378615,0.29673457,0.3357786,0.31625658,0.29673457,0.27721256,0.25769055,0.23816854,0.21083772,0.1835069,0.15617609,0.12884527,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.15617609,0.27330816,0.39044023,0.5075723,0.62470436,0.61689556,0.60908675,0.60127795,0.59346914,0.58566034,0.61689556,0.6481308,0.679366,0.7066968,0.737932,0.78088045,0.8238289,0.8667773,0.9058213,0.94876975,1.1635119,1.3782539,1.5969005,1.8116426,2.0263848,2.2918842,2.5534792,2.8189783,3.084478,3.349977,2.8658314,2.3816853,1.893635,1.4094892,0.92534333,0.9136301,0.9019169,0.8862993,0.8745861,0.8628729,0.96438736,1.0659018,1.1713207,1.2728351,1.3743496,1.1517987,0.92924774,0.7066968,0.48414588,0.26159495,0.28111696,0.29673457,0.31625658,0.3318742,0.3513962,0.45681506,0.5661383,0.6715572,0.78088045,0.8862993,1.3274968,1.7686942,2.2059872,2.6471848,3.0883822,2.9829633,2.8775444,2.7721257,2.6667068,2.5612879,2.9868677,3.4124475,3.8380275,4.263607,4.689187,4.911738,5.138193,5.3607445,5.5871997,5.813655,6.223617,6.6374836,7.0513506,7.461313,7.8751793,9.507219,11.139259,12.771299,14.40334,16.039284,16.937298,17.839214,18.737226,19.639143,20.537155,21.12672,21.712381,22.301945,22.887606,23.473267,24.289286,25.105307,25.921326,26.733442,27.549461,29.052658,30.555853,32.059048,33.55834,35.06153,33.02734,30.993145,28.958952,26.920853,24.88666,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.19912452,0.27330816,0.3513962,0.42557985,0.4997635,1.2259823,1.9482968,2.6745155,3.4007344,4.123049,4.814128,5.5013027,6.1884775,6.8756523,7.562827,6.785851,6.012779,5.2358036,4.462732,3.6857557,3.2016098,2.7135596,2.2255092,1.737459,1.2494087,1.2142692,1.175225,1.1361811,1.1010414,1.0619974,0.96438736,0.8628729,0.76135844,0.6637484,0.5622339,0.6754616,0.78868926,0.9019169,1.0112402,1.1244678,1.5383345,1.9482968,2.3621633,2.77603,3.1859922,2.9361105,2.6862288,2.436347,2.1864653,1.9365835,2.4012074,2.8619268,3.3265507,3.78727,4.251894,4.5017757,4.7516575,5.001539,5.251421,5.5013027,5.8370814,6.1767645,6.5125427,6.8483214,7.1880045,7.601871,8.011833,8.4257,8.835662,9.249529,8.538928,7.824422,7.113821,6.3993154,5.688714,5.462259,5.2358036,5.0132523,4.786797,4.564246,4.5876727,4.6110992,4.6384296,4.661856,4.689187,5.735567,6.785851,7.8361354,8.886419,9.936704,10.561408,11.186112,11.810817,12.439425,13.06413,12.939189,12.814248,12.689307,12.564366,12.439425,11.29934,10.163159,9.023073,7.8868923,6.7507114,6.676528,6.5984397,6.524256,6.4500723,6.375889,7.461313,8.550641,9.636065,10.725393,11.810817,11.986515,12.162213,12.337912,12.513609,12.689307,12.388668,12.08803,11.787391,11.486752,11.186112,11.623405,12.0606985,12.501896,12.939189,13.376482,17.37459,21.376602,25.37471,29.376722,33.374832,30.348919,27.326912,24.300999,21.275087,18.249176,19.498585,20.751898,22.001307,23.250715,24.500124,25.523077,26.549934,27.576794,28.599747,29.626604,33.726227,37.825848,41.925472,46.025093,50.124718,49.19937,48.27403,47.348686,46.423344,45.501904,40.898613,36.29923,31.699842,27.100456,22.50107,22.53621,22.575254,22.614298,22.649437,22.688482,21.626484,20.560583,19.498585,18.436588,17.37459,13.927003,10.475512,7.0240197,3.5764325,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,1.8233559,3.4632049,5.099149,6.7389984,8.374943,13.325725,18.276506,23.223385,28.174168,33.12495,36.92393,40.726818,44.525803,48.324787,52.12377,52.076916,52.02616,51.975403,51.924644,51.87389,42.362766,32.85164,23.336613,13.825488,4.3143644,4.939069,5.563773,6.1884775,6.813182,7.437886,6.66091,5.8878384,5.1108627,4.337791,3.5608149,7.8361354,12.111456,16.386776,20.662096,24.937418,27.861814,30.786211,33.71451,36.638912,39.56331,31.738886,23.914463,16.086138,8.261715,0.43729305,11.986515,23.535736,35.088863,46.638084,58.187305,53.201385,48.21156,43.225636,38.235813,33.24989,30.813543,28.373291,25.936945,23.500597,21.06425,18.936352,16.812357,14.688361,12.564366,10.436467,13.825488,17.210606,20.599627,23.988647,27.373764,26.58898,25.80029,25.0116,24.226816,23.438128,26.112642,28.787157,31.461674,34.13619,36.810703,34.635952,32.4612,30.286448,28.111696,25.936945,25.448895,24.960844,24.476698,23.988647,23.500597,19.475159,15.449719,11.424281,7.3988423,3.3734035,6.13772,8.898132,11.66245,14.426766,17.18718,14.051944,10.912805,7.773665,4.6384296,1.4992905,1.3509232,1.1986516,1.0502841,0.9019169,0.74964523,5.087436,9.425227,13.763018,18.10081,22.4386,19.96321,17.487818,15.012426,12.537036,10.061645,9.448653,8.835662,8.226576,7.6135845,7.000593,6.4891167,5.9737353,5.462259,4.950782,4.4393053,3.873167,3.310933,2.7486992,2.1864653,1.6242313,2.787743,3.951255,5.1108627,6.2743745,7.437886,9.499411,11.560935,13.626364,15.687888,17.749413,15.438006,13.1266,10.81129,8.499884,6.1884775,4.9742084,3.7638438,2.5495746,1.33921,0.12494087,0.8238289,1.5266213,2.2255092,2.9243972,3.6232853,3.338264,3.049338,2.7643168,2.475391,2.1864653,1.8116426,1.43682,1.0619974,0.6871748,0.31235218,0.44900626,0.58566034,0.7262188,0.8628729,0.999527,1.3743496,1.7491722,2.1239948,2.4988174,2.87364,3.4124475,3.951255,4.4861584,5.024966,5.563773,5.9737353,6.387602,6.801469,7.211431,7.6252975,6.13772,4.650143,3.1625657,1.6749885,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.27330816,0.5505207,0.8238289,1.1010414,1.3743496,1.1010414,0.8238289,0.5505207,0.27330816,0.0,0.0,0.0,0.0,0.0,0.0,0.23816854,0.47633708,0.7106012,0.94876975,1.1869383,1.9131571,2.639376,3.3616903,4.087909,4.814128,3.873167,2.9361105,1.999054,1.0619974,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.37482262,0.74964523,1.1244678,1.4992905,1.8741131,1.4992905,1.1244678,0.74964523,0.37482262,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21083772,0.42557985,0.63641757,0.8511597,1.0619974,0.92534333,0.78868926,0.6481308,0.5114767,0.37482262,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.113227665,0.22645533,0.3357786,0.44900626,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.58566034,0.61299115,0.63641757,0.6637484,0.6871748,0.77307165,0.8628729,0.94876975,1.038571,1.1244678,1.3860629,1.6515622,1.9131571,2.174752,2.436347,2.7252727,3.0141985,3.2992198,3.5881457,3.873167,3.310933,2.7486992,2.1864653,1.6242313,1.0619974,1.0619974,1.0619974,1.0619974,1.0619974,1.0619974,1.1869383,1.3118792,1.43682,1.5617609,1.6867018,1.3860629,1.0893283,0.78868926,0.48805028,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.30063897,0.41386664,0.5231899,0.63641757,0.74964523,0.8628729,0.97610056,1.0893283,1.1986516,1.3118792,1.4485333,1.5890918,1.7257458,1.8623998,1.999054,2.2879796,2.5769055,2.8619268,3.1508527,3.435874,3.3734035,3.310933,3.2484627,3.1859922,3.1235218,3.6506162,4.173806,4.7009,5.22409,5.7511845,7.7892823,9.823476,11.861574,13.899672,15.93777,17.085665,18.237463,19.389261,20.537155,21.688955,22.07549,22.462027,22.848562,23.239002,23.625538,24.148727,24.675823,25.199013,25.726107,26.249296,27.951616,29.65003,31.348446,33.050766,34.74918,32.449486,30.149794,27.850101,25.550407,23.250715,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.058566034,0.07027924,0.078088045,0.08980125,0.10151446,0.16008049,0.21864653,0.28111696,0.339683,0.39824903,1.1244678,1.8506867,2.5769055,3.2992198,4.025439,4.8687897,5.716045,6.559396,7.406651,8.250002,7.523783,6.79366,6.067441,5.3412223,4.6110992,4.025439,3.435874,2.8502135,2.260649,1.6749885,1.5695697,1.4641509,1.358732,1.2533131,1.1517987,1.077615,1.0034313,0.93315214,0.8589685,0.78868926,0.8433509,0.9019169,0.96048295,1.0190489,1.0737107,1.5227169,1.9717231,2.416825,2.8658314,3.310933,3.2289407,3.1469483,3.0649557,2.9829633,2.900971,3.2562714,3.611572,3.9668727,4.318269,4.6735697,4.7985106,4.919547,5.040583,5.165524,5.2865605,5.6262436,5.9620223,6.3017054,6.6374836,6.9732623,7.2036223,7.4300776,7.656533,7.8868923,8.113348,7.726812,7.336372,6.949836,6.5633,6.1767645,6.0205884,5.8644123,5.708236,5.5559645,5.3997884,5.212377,5.024966,4.8375545,4.650143,4.462732,5.716045,6.969358,8.218767,9.47208,10.725393,11.2642,11.806912,12.34572,12.884527,13.423335,13.212498,13.001659,12.786918,12.576079,12.361338,11.631214,10.897186,10.163159,9.433036,8.699008,8.663869,8.624825,8.58578,8.550641,8.511597,9.0035515,9.499411,9.991365,10.48332,10.975275,11.131451,11.291532,11.447707,11.603884,11.763964,11.896713,12.033368,12.166118,12.302772,12.439425,13.618555,14.801589,15.984623,17.167656,18.35069,21.36489,24.379087,27.393286,30.411388,33.425587,31.133703,28.845724,26.55384,24.26586,21.973976,22.356607,22.735334,23.114061,23.496693,23.87542,24.109684,24.343948,24.578213,24.816381,25.050644,28.080462,31.110277,34.140095,37.16991,40.199726,39.524265,38.8488,38.17334,37.501785,36.82632,33.792603,30.75888,27.729065,24.695345,21.661623,21.981785,22.301945,22.622107,22.942268,23.262428,22.048159,20.83389,19.615717,18.401447,17.18718,14.789876,12.392572,9.99527,7.5979667,5.2006636,5.02887,4.853172,4.6813784,4.5095844,4.337791,5.0054436,5.6730967,6.3407493,7.008402,7.676055,11.978706,16.281357,20.58401,24.88666,29.189312,32.84383,36.50226,40.160683,43.819107,47.473625,47.169083,46.86454,46.559998,46.255455,45.95091,38.149914,30.348919,22.547922,14.750832,6.949836,8.367134,9.784432,11.20173,12.619028,14.036326,12.103647,10.167064,8.23048,6.297801,4.3612175,7.703386,11.045554,14.391626,17.733795,21.075964,24.441559,27.80325,31.168842,34.53444,37.900032,30.395771,22.89151,15.383345,7.8790836,0.37482262,10.42085,20.462973,30.508999,40.555027,50.60105,46.442863,42.284676,38.126488,33.9683,29.814016,27.221493,24.62897,22.036446,19.443924,16.8514,15.84016,14.828919,13.821584,12.810344,11.799104,14.56342,17.323833,20.08815,22.848562,25.612879,25.179491,24.746101,24.316618,23.883228,23.44984,25.058455,26.67097,28.279585,29.888199,31.500717,30.75888,30.01314,29.271303,28.529467,27.78763,26.955994,26.124355,25.288813,24.457176,23.625538,20.263847,16.906061,13.544372,10.186585,6.824895,8.796618,10.764437,12.73616,14.703979,16.675701,13.622459,10.569217,7.5159745,4.466636,1.4133936,2.8306916,4.2479897,5.6652875,7.082586,8.499884,10.584834,12.6697855,14.754736,16.839687,18.924637,16.843592,14.766449,12.685403,10.604357,8.52331,7.9610763,7.3988423,6.8366084,6.2743745,5.7121406,5.309987,4.9078336,4.50568,4.1035266,3.7013733,3.2289407,2.7604125,2.2918842,1.8194515,1.3509232,2.2918842,3.2289407,4.169902,5.1108627,6.0518236,7.832231,9.616543,11.39695,13.181262,14.96167,13.009468,11.057267,9.105066,7.152865,5.2006636,4.1894236,3.1781836,2.1708477,1.1596074,0.14836729,0.79649806,1.4446288,2.0927596,2.7408905,3.3890212,3.06886,2.7486992,2.4285383,2.1083772,1.7882162,1.6749885,1.5617609,1.4485333,1.33921,1.2259823,1.1517987,1.0737107,0.999527,0.92534333,0.8511597,1.1517987,1.4485333,1.7491722,2.0498111,2.35045,2.87364,3.4007344,3.9239242,4.4510183,4.9742084,5.2006636,5.4310236,5.657479,5.883934,6.114294,5.009348,3.9083066,2.803361,1.7023194,0.60127795,0.5544251,0.5114767,0.46462387,0.42167544,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.21864653,0.44119745,0.659844,0.8784905,1.1010414,0.8784905,0.659844,0.44119745,0.21864653,0.0,0.0,0.0,0.0,0.0,0.0,0.19131571,0.37872702,0.5700427,0.76135844,0.94876975,2.4910088,4.0332475,5.579391,7.1216297,8.663869,6.949836,5.2358036,3.5256753,1.8116426,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.16008049,0.19522011,0.23035973,0.26549935,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.30063897,0.60127795,0.9019169,1.1986516,1.4992905,1.2103647,0.92143893,0.62860876,0.339683,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1835069,0.3631094,0.5466163,0.7301232,0.9136301,0.8941081,0.8706817,0.8511597,0.8316377,0.81211567,0.7340276,0.6559396,0.58175594,0.5036679,0.42557985,0.3631094,0.30454338,0.24597734,0.1835069,0.12494087,0.12103647,0.12103647,0.11713207,0.113227665,0.113227665,0.11713207,0.12103647,0.12884527,0.13274968,0.13665408,0.10932326,0.08199245,0.05466163,0.027330816,0.0,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,0.60908675,0.58956474,0.57394713,0.5544251,0.5388075,0.5661383,0.59346914,0.62079996,0.6481308,0.6754616,0.80821127,0.94486535,1.0815194,1.2142692,1.3509232,1.5617609,1.7686942,1.979532,2.1903696,2.4012074,2.5612879,2.7213683,2.8814487,3.0415294,3.2016098,2.7838387,2.366068,1.9482968,1.5305257,1.1127546,1.2025559,1.2923572,1.3821584,1.4719596,1.5617609,1.6632754,1.7608855,1.8623998,1.9639144,2.0615244,1.7257458,1.3860629,1.0502841,0.7106012,0.37482262,0.3553006,0.3357786,0.31625658,0.29673457,0.27330816,0.3435874,0.40996224,0.47633708,0.5466163,0.61299115,0.7066968,0.79649806,0.8902037,0.98390937,1.0737107,1.1908426,1.3040704,1.4212024,1.53443,1.6515622,1.893635,2.1396124,2.3855898,2.631567,2.87364,2.9087796,2.9400148,2.97125,3.0063896,3.0376248,3.4983444,3.9629683,4.423688,4.8883114,5.349031,7.125534,8.902037,10.674636,12.4511385,14.223738,15.328683,16.43363,17.538574,18.64352,19.748466,20.076437,20.400501,20.724567,21.048632,21.376602,21.895887,22.419077,22.942268,23.465458,23.988647,25.620687,27.252728,28.884768,30.516808,32.14885,30.520712,28.89648,27.268345,25.64021,24.012074,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.046852827,0.05075723,0.058566034,0.06637484,0.07418364,0.12103647,0.1639849,0.21083772,0.25378615,0.30063897,1.0268579,1.7491722,2.475391,3.2016098,3.9239242,4.927356,5.930787,6.9342184,7.9337454,8.937177,8.257811,7.578445,6.899079,6.2158084,5.5364423,4.8492675,4.1620927,3.474918,2.787743,2.1005683,1.9287747,1.7530766,1.5812829,1.4094892,1.2376955,1.1908426,1.1478943,1.1010414,1.0580931,1.0112402,1.0151446,1.0190489,1.0190489,1.0229534,1.0268579,1.5070993,1.9912452,2.4714866,2.9556324,3.435874,3.521771,3.6076677,3.6935644,3.775557,3.8614538,4.1113358,4.357313,4.60329,4.853172,5.099149,5.095245,5.0913405,5.083532,5.0796275,5.0757227,5.4115014,5.7511845,6.086963,6.426646,6.7624245,6.805373,6.8483214,6.89127,6.9342184,6.9732623,6.910792,6.8483214,6.785851,6.7233806,6.66091,6.578918,6.493021,6.407124,6.321227,6.239235,5.8370814,5.4388323,5.036679,4.6384296,4.2362766,5.6926184,7.1489606,8.601398,10.05774,11.514082,11.966993,12.423808,12.8767185,13.333533,13.786445,13.4858055,13.189071,12.888432,12.587793,12.287154,11.959184,11.631214,11.303245,10.979179,10.651209,10.651209,10.651209,10.651209,10.651209,10.651209,10.545791,10.444276,10.342762,10.241247,10.135828,10.276386,10.416945,10.557504,10.698062,10.838621,11.408664,11.978706,12.548749,13.118792,13.688834,15.613705,17.542479,19.471254,21.396124,23.3249,25.355188,27.385477,29.415766,31.446056,33.476345,31.918488,30.364536,28.810585,27.256632,25.698776,25.210726,24.718771,24.23072,23.738766,23.250715,22.696291,22.141865,21.583536,21.02911,20.474686,22.434696,24.394705,26.354715,28.314726,30.274734,29.849155,29.423576,28.997995,28.57632,28.15074,26.68659,25.218534,23.754383,22.290232,20.826082,21.42736,22.028637,22.63382,23.235098,23.836376,22.469835,21.103294,19.736753,18.366308,16.999767,15.656653,14.309634,12.96652,11.619501,10.276386,9.917182,9.561881,9.202676,8.843472,8.488171,8.183627,7.882988,7.578445,7.277806,6.9732623,10.631687,14.286208,17.94073,21.59525,25.24977,28.763731,32.281597,35.79556,39.30952,42.823483,42.265156,41.706825,41.144592,40.58626,40.02403,33.937065,27.850101,21.763138,15.676175,9.589212,11.799104,14.008995,16.218887,18.42878,20.63867,17.542479,14.446288,11.354002,8.257811,5.1616197,7.570636,9.983557,12.392572,14.801589,17.210606,21.017397,24.82419,28.627077,32.43387,36.23676,29.052658,21.868557,14.6805525,7.4964523,0.31235218,8.85128,17.394112,25.93304,34.471966,43.010895,39.684345,36.357796,33.031242,29.700788,26.374237,23.629442,20.880743,18.132044,15.383345,12.63855,12.743969,12.849388,12.950902,13.056321,13.16174,15.3013525,17.437061,19.576674,21.712381,23.84809,23.773905,23.695818,23.61773,23.53964,23.461554,24.00817,24.55088,25.097498,25.644114,26.186827,26.877905,27.568985,28.256159,28.947239,29.638317,28.459188,27.283962,26.104834,24.925705,23.750479,21.056442,18.3585,15.664462,12.970425,10.276386,11.4516115,12.630741,13.805966,14.985096,16.164225,13.196879,10.229534,7.2582836,4.290938,1.3235924,4.31046,7.2934237,10.280292,13.263254,16.250122,16.082233,15.914344,15.746454,15.578565,15.410676,13.727879,12.041177,10.358379,8.671678,6.98888,6.473499,5.9620223,5.4505453,4.939069,4.423688,4.1308575,3.8419318,3.5491016,3.2562714,2.9634414,2.5847144,2.2059872,1.8311646,1.4524376,1.0737107,1.7921207,2.5105307,3.2289407,3.9434462,4.661856,6.165051,7.6682463,9.171441,10.670732,12.173926,10.58093,8.991838,7.3988423,5.805846,4.21285,3.4046388,2.5964274,1.7882162,0.98390937,0.1756981,0.76916724,1.3665408,1.9600099,2.5534792,3.1508527,2.795552,2.4441557,2.0927596,1.7413634,1.3860629,1.5383345,1.6867018,1.8389735,1.9873407,2.135708,1.8506867,1.5617609,1.2767396,0.9878138,0.698888,0.92534333,1.1517987,1.3743496,1.6008049,1.8233559,2.338737,2.8502135,3.3616903,3.873167,4.388548,4.4314966,4.4705405,4.513489,4.5564375,4.5993857,3.8809757,3.1664703,2.4480603,1.7296503,1.0112402,0.96048295,0.9058213,0.8550641,0.80430686,0.74964523,0.60127795,0.44900626,0.30063897,0.14836729,0.0,0.1639849,0.3318742,0.4958591,0.659844,0.8238289,0.659844,0.4958591,0.3318742,0.1639849,0.0,0.0,0.0,0.0,0.0,0.0,0.14055848,0.28502136,0.42557985,0.5700427,0.7106012,3.0727646,5.4310236,7.793187,10.151445,12.513609,10.0265045,7.5394006,5.0483923,2.5612879,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.3513962,0.3240654,0.30063897,0.27330816,0.24988174,0.32016098,0.39044023,0.46071947,0.5309987,0.60127795,0.48024148,0.359205,0.23816854,0.12103647,0.0,0.22645533,0.44900626,0.6754616,0.9019169,1.1244678,0.92143893,0.7145056,0.5114767,0.30454338,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15227169,0.30454338,0.45681506,0.60908675,0.76135844,0.8589685,0.95657855,1.0541886,1.1517987,1.2494087,1.1557031,1.0659018,0.97219616,0.8784905,0.78868926,0.6676528,0.5466163,0.42557985,0.30844778,0.18741131,0.1717937,0.15227169,0.13665408,0.11713207,0.10151446,0.10932326,0.12103647,0.12884527,0.14055848,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.13665408,0.27330816,0.41386664,0.5505207,0.6871748,0.6520352,0.61689556,0.58175594,0.5466163,0.5114767,0.5427119,0.57394713,0.60127795,0.63251317,0.6637484,0.8433509,1.0268579,1.2103647,1.3938715,1.5734742,1.7335546,1.8897307,2.0459068,2.2059872,2.3621633,2.3933985,2.4285383,2.4597735,2.4910088,2.5261483,2.25284,1.979532,1.7062237,1.43682,1.1635119,1.3431144,1.5227169,1.7023194,1.8819219,2.0615244,2.135708,2.2137961,2.2879796,2.3621633,2.436347,2.0615244,1.6867018,1.3118792,0.93705654,0.5622339,0.5231899,0.48414588,0.44119745,0.40215343,0.3631094,0.38653582,0.40605783,0.42948425,0.45291066,0.47633708,0.5466163,0.62079996,0.6910792,0.76526284,0.8394465,0.92924774,1.0229534,1.116659,1.2064602,1.3001659,1.5031948,1.7062237,1.9092526,2.1083772,2.3114061,2.4402514,2.5690966,2.6940374,2.822883,2.951728,3.349977,3.7482262,4.1503797,4.548629,4.950782,6.461786,7.9766936,9.487698,10.998701,12.513609,13.571702,14.633699,15.6917925,16.75379,17.811884,18.073479,18.338978,18.600573,18.862167,19.123762,19.646952,20.166237,20.685524,21.20481,21.724094,23.289759,24.855425,26.42109,27.986755,29.548515,28.595842,27.639263,26.68659,25.730011,24.773432,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.031235218,0.03513962,0.039044023,0.046852827,0.05075723,0.078088045,0.10932326,0.14055848,0.1717937,0.19912452,0.92534333,1.6515622,2.3738766,3.1000953,3.8263142,4.985922,6.1455293,7.3051367,8.464745,9.6243515,8.991838,8.359325,7.726812,7.094299,6.461786,5.6730967,4.8883114,4.0996222,3.310933,2.5261483,2.2840753,2.0459068,1.8038338,1.5656652,1.3235924,1.3079748,1.2884527,1.2728351,1.2533131,1.2376955,1.1869383,1.1322767,1.0815194,1.0268579,0.97610056,1.4914817,2.0107672,2.5261483,3.0454338,3.5608149,3.814601,4.068387,4.318269,4.572055,4.825841,4.9663997,5.1069584,5.2436123,5.3841705,5.5247293,5.3919797,5.2592297,5.12648,4.9937305,4.860981,5.2006636,5.5364423,5.8761253,6.211904,6.551587,6.407124,6.266566,6.1221027,5.9815445,5.8370814,6.098676,6.364176,6.6257706,6.8873653,7.1489606,7.1333427,7.1216297,7.1060123,7.0903945,7.0747766,6.461786,5.8487945,5.2358036,4.6267166,4.0137253,5.6691923,7.328563,8.98403,10.6434,12.298867,12.6697855,13.040704,13.411622,13.778636,14.149553,13.763018,13.376482,12.986042,12.599506,12.212971,12.291059,12.369146,12.44333,12.521418,12.599506,12.63855,12.67369,12.712734,12.751778,12.786918,12.091934,11.393045,10.694158,9.999174,9.300286,9.421323,9.546264,9.6673,9.788337,9.913278,10.916709,11.924045,12.927476,13.930907,14.938243,17.608854,20.28337,22.953981,25.628496,28.299107,29.345488,30.391867,31.434343,32.48072,33.523197,32.703274,31.883348,31.063425,30.2435,29.423576,28.064844,26.706112,25.343475,23.984743,22.62601,21.278992,19.935879,18.58886,17.245745,15.8987255,16.788929,17.679134,18.569338,19.459541,20.349745,20.174046,19.998348,19.826555,19.650856,19.475159,19.576674,19.678188,19.783606,19.88512,19.986635,20.872934,21.759233,22.641628,23.527927,24.414227,22.89151,21.372698,19.853886,18.33117,16.812357,16.519526,16.226696,15.933866,15.641035,15.348206,14.809398,14.2666855,13.723974,13.181262,12.63855,11.365715,10.09288,8.8200445,7.5472097,6.2743745,9.280765,12.291059,15.297448,18.303837,21.314133,24.683632,28.057035,31.430439,34.80384,38.17334,37.361225,36.545204,35.729183,34.913166,34.101048,29.724215,25.351284,20.97445,16.601519,12.224684,15.227169,18.229654,21.23214,24.234625,27.23711,22.981312,18.729418,14.473619,10.217821,5.9620223,7.4417906,8.917655,10.393518,11.873287,13.349152,17.593237,21.841227,26.085312,30.329397,34.573483,27.709543,20.845604,13.981665,7.113821,0.24988174,7.2856145,14.321347,21.353176,28.388908,35.42464,32.925823,30.430912,27.932095,25.433277,22.938364,20.033487,17.132517,14.231546,11.326671,8.4257,9.643873,10.865952,12.084125,13.306203,14.524376,16.039284,17.550287,19.061293,20.5762,22.087204,22.364416,22.641628,22.91884,23.196054,23.473267,22.953981,22.434696,21.91541,21.396124,20.872934,22.99693,25.120924,27.241014,29.36501,31.489004,29.966288,28.443571,26.920853,25.398136,23.87542,21.84513,19.814842,17.784552,15.754263,13.723974,14.11051,14.493141,14.879677,15.266212,15.648844,12.767395,9.885946,7.000593,4.1191444,1.2376955,5.7902284,10.342762,14.895294,19.447828,24.00036,21.579632,19.158901,16.738173,14.321347,11.900618,10.608261,9.319808,8.031356,6.7389984,5.4505453,4.985922,4.5252023,4.0605783,3.5998588,3.1391394,2.9556324,2.7721257,2.5886188,2.4090161,2.2255092,1.9404879,1.6554666,1.3704453,1.0854238,0.80040246,1.2962615,1.7882162,2.2840753,2.7799344,3.2757936,4.4978714,5.7199492,6.942027,8.164105,9.386183,8.156297,6.9225054,5.688714,4.4588275,3.2250361,2.619854,2.0146716,1.4094892,0.80430686,0.19912452,0.7418364,1.2845483,1.8272603,2.3699722,2.912684,2.5261483,2.1435168,1.756981,1.3743496,0.9878138,1.4016805,1.8116426,2.2255092,2.639376,3.049338,2.5495746,2.0498111,1.5500476,1.0502841,0.5505207,0.698888,0.8511597,0.999527,1.1517987,1.3001659,1.7999294,2.2996929,2.7994564,3.2992198,3.7989833,3.6584249,3.513962,3.3734035,3.2289407,3.0883822,2.7565079,2.4207294,2.0888553,1.756981,1.4251068,1.3665408,1.3040704,1.2455044,1.1869383,1.1244678,0.9019169,0.6754616,0.44900626,0.22645533,0.0,0.10932326,0.21864653,0.3318742,0.44119745,0.5505207,0.44119745,0.3318742,0.21864653,0.10932326,0.0,0.0,0.0,0.0,0.0,0.0,0.093705654,0.19131571,0.28502136,0.37872702,0.47633708,3.6545205,6.8287997,10.006983,13.185166,16.36335,13.09927,9.839094,6.575013,3.310933,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.113227665,0.22645533,0.3357786,0.44900626,0.5622339,0.5231899,0.48805028,0.44900626,0.41386664,0.37482262,0.48024148,0.58566034,0.6910792,0.79649806,0.9019169,0.71841,0.5388075,0.359205,0.1796025,0.0,0.14836729,0.30063897,0.44900626,0.60127795,0.74964523,0.62860876,0.5114767,0.39044023,0.26940376,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12103647,0.24597734,0.3670138,0.48805028,0.61299115,0.8277333,1.0424755,1.2572175,1.4719596,1.6867018,1.5812829,1.4719596,1.3665408,1.2572175,1.1517987,0.96829176,0.78868926,0.60908675,0.42948425,0.24988174,0.21864653,0.1835069,0.15227169,0.12103647,0.08589685,0.10151446,0.11713207,0.13274968,0.14836729,0.1639849,0.12884527,0.09761006,0.06637484,0.031235218,0.0,0.14836729,0.30063897,0.44900626,0.60127795,0.74964523,0.698888,0.6442264,0.59346914,0.5388075,0.48805028,0.5192855,0.5544251,0.58566034,0.61689556,0.6481308,0.8784905,1.1088502,1.33921,1.5695697,1.7999294,1.9053483,2.0107672,2.1161861,2.2216048,2.3231194,2.2294137,2.135708,2.0380979,1.9443923,1.8506867,1.7218413,1.5969005,1.4680552,1.33921,1.2142692,1.4836729,1.7530766,2.0224805,2.2918842,2.5612879,2.612045,2.6628022,2.7135596,2.7643168,2.8111696,2.4012074,1.9873407,1.5734742,1.1635119,0.74964523,0.6910792,0.62860876,0.5700427,0.5114767,0.44900626,0.42557985,0.40605783,0.38263142,0.359205,0.3357786,0.39044023,0.44119745,0.4958591,0.5466163,0.60127795,0.6715572,0.7418364,0.80821127,0.8784905,0.94876975,1.1088502,1.2689307,1.4290112,1.5890918,1.7491722,1.9717231,2.194274,2.416825,2.639376,2.8619268,3.2016098,3.5373883,3.873167,4.21285,4.548629,5.801942,7.0513506,8.300759,9.550168,10.799577,11.814721,12.829865,13.845011,14.860155,15.875299,16.074425,16.273548,16.476578,16.675701,16.874826,17.394112,17.909492,18.42878,18.94416,19.463446,20.958832,22.458122,23.953508,25.452799,26.948185,26.667067,26.38595,26.10093,25.819813,25.538694,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.015617609,0.015617609,0.019522011,0.023426414,0.023426414,0.039044023,0.05466163,0.07027924,0.08589685,0.10151446,0.8238289,1.5500476,2.2762666,2.998581,3.7247996,5.040583,6.3602715,7.676055,8.995743,10.311526,9.725866,9.14411,8.55845,7.9727893,7.387129,6.5008297,5.610626,4.7243266,3.8380275,2.951728,2.6432803,2.3348327,2.0263848,1.7218413,1.4133936,1.4212024,1.4329157,1.4407244,1.4524376,1.4641509,1.3548276,1.2494087,1.1400855,1.0307622,0.92534333,1.475864,2.0302892,2.5808098,3.135235,3.6857557,4.1074314,4.5291066,4.9468775,5.368553,5.786324,5.8214636,5.852699,5.883934,5.919074,5.950309,5.688714,5.4310236,5.169429,4.911738,4.650143,4.985922,5.3256044,5.661383,6.001066,6.336845,6.008875,5.6809053,5.35684,5.02887,4.7009,5.2865605,5.8761253,6.461786,7.0513506,7.6370106,7.6916723,7.746334,7.800996,7.8556576,7.914223,7.08649,6.262661,5.4388323,4.6110992,3.78727,5.645766,7.5081654,9.366661,11.229061,13.087557,13.372578,13.657599,13.94262,14.227642,14.512663,14.036326,13.563893,13.087557,12.611219,12.138786,12.619028,13.103174,13.583415,14.067561,14.551707,14.625891,14.700074,14.774258,14.848442,14.92653,13.634172,12.341816,11.045554,9.753197,8.460839,8.566258,8.671678,8.777096,8.882515,8.987934,10.4286585,11.869383,13.306203,14.746927,16.187653,19.604004,23.02426,26.440613,29.856964,33.273315,33.335785,33.394352,33.45682,33.51539,33.573956,33.491962,33.406067,33.320168,33.234272,33.148376,30.91896,28.689548,26.460135,24.23072,22.001307,19.865599,17.72989,15.594183,13.458474,11.326671,11.143164,10.963562,10.783959,10.604357,10.424754,10.498938,10.573121,10.651209,10.725393,10.799577,12.470661,14.141745,15.808925,17.48001,19.151093,20.31851,21.485926,22.653341,23.820759,24.988174,23.313187,21.642101,19.971018,18.296028,16.624945,17.386303,18.143757,18.905115,19.666473,20.423927,19.69771,18.97149,18.241367,17.515148,16.788929,14.543899,12.302772,10.061645,7.816613,5.575486,7.9337454,10.295909,12.654168,15.016331,17.37459,20.60353,23.836376,27.065317,30.294256,33.523197,32.453392,31.383585,30.31378,29.243973,28.174168,25.511364,22.848562,20.18576,17.526861,14.864059,18.659138,22.454218,26.249296,30.044374,33.839455,28.42405,23.008642,17.593237,12.177831,6.7624245,7.309041,7.8517528,8.398369,8.941081,9.487698,14.17298,18.858263,23.543545,28.228828,32.914112,26.366428,19.82265,13.2788725,6.7311897,0.18741131,5.716045,11.248583,16.777216,22.305851,27.838388,26.171207,24.504028,22.832945,21.165764,19.498585,16.441439,13.384291,10.327144,7.269997,4.21285,6.547683,8.882515,11.217348,13.55218,15.8870125,16.773312,17.663515,18.549814,19.436115,20.326319,20.958832,21.591345,22.223858,22.85637,23.488884,21.903696,20.31851,18.733322,17.148134,15.562947,19.115953,22.672863,26.22587,29.78278,33.335785,31.469482,29.603178,27.736874,25.866665,24.00036,22.63382,21.271183,19.904642,18.538101,17.175465,16.769407,16.359446,15.953387,15.543426,15.137367,12.341816,9.542359,6.746807,3.9473507,1.1517987,7.269997,13.388195,19.510298,25.628496,31.750599,27.07703,22.40346,17.733795,13.0602255,8.386656,7.492548,6.5984397,5.704332,4.806319,3.912211,3.4983444,3.0883822,2.6745155,2.260649,1.8506867,1.7765031,1.7062237,1.6320401,1.5617609,1.4875772,1.2962615,1.1010414,0.9097257,0.71841,0.5231899,0.79649806,1.0698062,1.3431144,1.6164225,1.8858263,2.8306916,3.7716527,4.716518,5.657479,6.5984397,5.727758,4.853172,3.9824903,3.1118085,2.2372224,1.8350691,1.4329157,1.0307622,0.62860876,0.22645533,0.7145056,1.2064602,1.6945106,2.1864653,2.6745155,2.2567444,1.8389735,1.4212024,1.0034313,0.58566034,1.261122,1.9365835,2.612045,3.2875066,3.9629683,3.2484627,2.5378613,1.8233559,1.1127546,0.39824903,0.47633708,0.5505207,0.62470436,0.698888,0.77307165,1.261122,1.7491722,2.2372224,2.7252727,3.213323,2.8853533,2.5573835,2.2294137,1.901444,1.5734742,1.6281357,1.678893,1.7335546,1.7843118,1.8389735,1.7686942,1.7023194,1.6359446,1.5656652,1.4992905,1.1986516,0.9019169,0.60127795,0.30063897,0.0,0.05466163,0.10932326,0.1639849,0.21864653,0.27330816,0.21864653,0.1639849,0.10932326,0.05466163,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.093705654,0.14055848,0.19131571,0.23816854,4.2323723,8.226576,12.220779,16.218887,20.21309,16.175938,12.138786,8.101635,4.0605783,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14836729,0.30063897,0.44900626,0.60127795,0.74964523,0.698888,0.6481308,0.60127795,0.5505207,0.4997635,0.64032197,0.78088045,0.92143893,1.0580931,1.1986516,0.96048295,0.71841,0.48024148,0.23816854,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.339683,0.30454338,0.26940376,0.23426414,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.093705654,0.1835069,0.27721256,0.3709182,0.46071947,0.79649806,1.1283722,1.4602464,1.7921207,2.1239948,2.0029583,1.8819219,1.756981,1.6359446,1.5110037,1.2728351,1.0307622,0.79259366,0.5544251,0.31235218,0.26549935,0.21864653,0.1717937,0.12103647,0.07418364,0.093705654,0.113227665,0.13665408,0.15617609,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.1639849,0.3240654,0.48805028,0.6481308,0.81211567,0.7418364,0.6715572,0.60127795,0.5309987,0.46071947,0.4958591,0.5309987,0.5661383,0.60127795,0.63641757,0.9136301,1.1908426,1.4719596,1.7491722,2.0263848,2.077142,2.1318035,2.182561,2.233318,2.2879796,2.0654287,1.8428779,1.620327,1.397776,1.175225,1.1908426,1.2103647,1.2259823,1.2455044,1.261122,1.6242313,1.9834363,2.3426414,2.7018464,3.0610514,3.0883822,3.1118085,3.1391394,3.1625657,3.1859922,2.736986,2.2879796,1.8389735,1.3860629,0.93705654,0.8589685,0.77697605,0.698888,0.61689556,0.5388075,0.46852827,0.40215343,0.3357786,0.26940376,0.19912452,0.23426414,0.26549935,0.29673457,0.3318742,0.3631094,0.40996224,0.45681506,0.5036679,0.5544251,0.60127795,0.71841,0.8355421,0.95267415,1.0698062,1.1869383,1.5031948,1.8233559,2.1396124,2.455869,2.77603,3.049338,3.3265507,3.5998588,3.873167,4.1503797,5.138193,6.126007,7.113821,8.101635,9.085544,10.05774,11.0260315,11.998228,12.96652,13.938716,14.07537,14.212025,14.348679,14.489237,14.625891,15.141272,15.656653,16.168129,16.683512,17.198893,18.631807,20.06082,21.48983,22.91884,24.351757,24.738293,25.128733,25.519173,25.909613,26.300053,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7262188,1.4485333,2.174752,2.900971,3.6232853,5.099149,6.575013,8.050878,9.526741,10.998701,10.4637985,9.924991,9.386183,8.85128,8.312472,7.3246584,6.336845,5.349031,4.3612175,3.3734035,2.998581,2.6237583,2.2489357,1.8741131,1.4992905,1.5383345,1.5734742,1.6125181,1.6515622,1.6867018,1.5266213,1.3626363,1.1986516,1.038571,0.8745861,1.4641509,2.0498111,2.639376,3.2250361,3.8106966,4.4002614,4.985922,5.575486,6.1611466,6.7507114,6.676528,6.5984397,6.524256,6.4500723,6.375889,5.989353,5.5989127,5.212377,4.825841,4.4393053,4.775084,5.1108627,5.4505453,5.786324,6.126007,5.610626,5.099149,4.5876727,4.0761957,3.5608149,4.474445,5.388075,6.3017054,7.211431,8.125061,8.250002,8.374943,8.499884,8.624825,8.749765,7.7111945,6.676528,5.6379566,4.5993857,3.5608149,5.6262436,7.687768,9.749292,11.810817,13.8762455,14.07537,14.274494,14.473619,14.676648,14.875772,14.313539,13.751305,13.189071,12.626837,12.0606985,12.950902,13.837202,14.723501,15.613705,16.500004,16.613232,16.72646,16.835783,16.94901,17.062239,15.176412,13.286681,11.400854,9.511124,7.6252975,7.7111945,7.800996,7.8868923,7.9766936,8.062591,9.936704,11.810817,13.688834,15.562947,17.437061,21.599154,25.761246,29.92334,34.089336,38.25143,37.326084,36.40074,35.4754,34.550056,33.624714,34.27675,34.924877,35.576912,36.225044,36.873177,33.776985,30.67689,27.576794,24.476698,21.376602,18.448301,15.523903,12.599506,9.675109,6.7507114,5.5013027,4.251894,2.998581,1.7491722,0.4997635,0.8238289,1.1517987,1.475864,1.7999294,2.1239948,5.3607445,8.601398,11.838148,15.074897,18.311647,19.764084,21.212618,22.66115,24.113588,25.562122,23.738766,21.911505,20.08815,18.26089,16.437534,18.249176,20.06082,21.876366,23.68801,25.499651,24.586021,23.676296,22.762665,21.849035,20.93931,17.725986,14.512663,11.29934,8.086017,4.8765984,6.5867267,8.300759,10.010887,11.72492,13.438952,16.52343,19.611813,22.700195,25.788576,28.873055,27.549461,26.22587,24.898373,23.574781,22.251188,21.298513,20.349745,19.400974,18.448301,17.49953,22.087204,26.674877,31.262548,35.85022,40.437893,33.86288,27.287867,20.712854,14.13784,7.562827,7.1762915,6.785851,6.3993154,6.012779,5.6262436,10.748819,15.875299,21.00178,26.124355,31.250835,25.023314,18.799696,12.576079,6.348558,0.12494087,4.1503797,8.175818,12.201257,16.226696,20.24823,19.412687,18.573242,17.7377,16.898252,16.062712,12.849388,9.636065,6.426646,3.213323,0.0,3.4514916,6.899079,10.350571,13.798158,17.24965,17.511244,17.776743,18.038338,18.299932,18.56153,19.549341,20.537155,21.52497,22.512783,23.500597,20.849508,18.19842,15.551234,12.900145,10.249056,15.238882,20.224804,25.210726,30.200552,35.186474,32.97658,30.762785,28.548988,26.339098,24.125301,23.426414,22.723621,22.024733,21.325846,20.623053,19.4244,18.22575,17.023193,15.824542,14.625891,11.912332,9.198771,6.4891167,3.775557,1.0619974,8.749765,16.437534,24.125301,31.81307,39.50084,32.57443,25.651922,18.725513,11.799104,4.8765984,4.376835,3.873167,3.3734035,2.87364,2.3738766,2.0107672,1.6515622,1.2884527,0.92534333,0.5622339,0.60127795,0.63641757,0.6754616,0.7106012,0.74964523,0.6481308,0.5505207,0.44900626,0.3513962,0.24988174,0.30063897,0.3513962,0.39824903,0.44900626,0.4997635,1.1635119,1.8233559,2.4871042,3.1508527,3.8106966,3.2992198,2.787743,2.2762666,1.7608855,1.2494087,1.0502841,0.8511597,0.6481308,0.44900626,0.24988174,0.6871748,1.1244678,1.5617609,1.999054,2.436347,1.9873407,1.5383345,1.0893283,0.63641757,0.18741131,1.1244678,2.0615244,2.998581,3.9356375,4.8765984,3.951255,3.0259118,2.1005683,1.175225,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.7262188,1.1986516,1.6749885,2.1513257,2.6237583,2.1122816,1.6008049,1.0893283,0.57394713,0.062470436,0.4997635,0.93705654,1.3743496,1.8116426,2.2489357,2.174752,2.1005683,2.0263848,1.9482968,1.8741131,1.4992905,1.1244678,0.74964523,0.37482262,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,4.814128,9.6243515,14.438479,19.248703,24.062832,19.248703,14.438479,9.6243515,4.814128,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18741131,0.37482262,0.5622339,0.74964523,0.93705654,0.8745861,0.81211567,0.74964523,0.6871748,0.62470436,0.80040246,0.97610056,1.1517987,1.3235924,1.4992905,1.1986516,0.9019169,0.60127795,0.30063897,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.76135844,1.2142692,1.6632754,2.1122816,2.5612879,2.4246337,2.2879796,2.1513257,2.0107672,1.8741131,1.5734742,1.2767396,0.97610056,0.6754616,0.37482262,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.1756981,0.3513962,0.5231899,0.698888,0.8745861,0.78868926,0.698888,0.61299115,0.5231899,0.43729305,0.47633708,0.5114767,0.5505207,0.58566034,0.62470436,0.94876975,1.2767396,1.6008049,1.9248703,2.2489357,2.2489357,2.2489357,2.2489357,2.2489357,2.2489357,1.901444,1.5500476,1.1986516,0.8511597,0.4997635,0.6637484,0.8238289,0.9878138,1.1517987,1.3118792,1.7608855,2.2137961,2.6628022,3.1118085,3.5608149,3.5608149,3.5608149,3.5608149,3.5608149,3.5608149,3.076669,2.5886188,2.1005683,1.6125181,1.1244678,1.0268579,0.92534333,0.8238289,0.7262188,0.62470436,0.5114767,0.39824903,0.28892577,0.1756981,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.14836729,0.1756981,0.19912452,0.22645533,0.24988174,0.3240654,0.39824903,0.47633708,0.5505207,0.62470436,1.038571,1.4485333,1.8623998,2.2762666,2.6862288,2.900971,3.1118085,3.3265507,3.5373883,3.7482262,4.474445,5.2006636,5.9268827,6.649197,7.375416,8.300759,9.226103,10.151445,11.076789,11.998228,12.076316,12.150499,12.224684,12.298867,12.373051,12.888432,13.399908,13.911386,14.426766,14.938243,16.300879,17.663515,19.026152,20.388788,21.751425,22.813423,23.87542,24.937418,25.999414,27.061413,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.60127795,1.1986516,1.7999294,2.4012074,2.998581,4.454923,5.911265,7.363703,8.8200445,10.276386,10.03041,9.784432,9.538455,9.296382,9.050405,7.9259367,6.805373,5.6809053,4.560342,3.435874,3.1157131,2.7994564,2.4792955,2.1591344,1.8389735,1.9443923,2.0459068,2.1513257,2.2567444,2.3621633,2.1669433,1.9717231,1.7765031,1.5812829,1.3860629,2.018576,2.6471848,3.2757936,3.9083066,4.5369153,5.298274,6.055728,6.817086,7.578445,8.335898,8.1992445,8.062591,7.9259367,7.7892823,7.648724,7.2036223,6.754616,6.3056097,5.860508,5.4115014,5.5091114,5.602817,5.6965227,5.794133,5.8878384,5.376362,4.8687897,4.357313,3.8458362,3.338264,4.2362766,5.134289,6.028397,6.9264097,7.824422,8.121157,8.421796,8.718531,9.0152645,9.311999,8.335898,7.363703,6.387602,5.4115014,4.4393053,5.9932575,7.5472097,9.101162,10.6590185,12.212971,12.240301,12.267632,12.294963,12.322293,12.349625,11.877192,11.404759,10.932326,10.459893,9.987461,10.936231,11.881096,12.829865,13.778636,14.723501,15.145176,15.566852,15.984623,16.406298,16.82407,15.516094,14.204215,12.89624,11.584361,10.276386,10.901091,11.525795,12.150499,12.775204,13.399908,15.008522,16.62104,18.229654,19.838268,21.450787,24.211199,26.971611,29.732023,32.488533,35.248943,34.007343,32.765743,31.524143,30.278639,29.037039,29.681267,30.321589,30.965815,31.606136,32.250362,32.164467,32.074665,31.988768,31.898966,31.81307,29.376722,26.936472,24.500124,22.063778,19.623526,17.780647,15.933866,14.090988,12.244205,10.401327,10.303718,10.2100115,10.116306,10.018696,9.924991,11.084598,12.244205,13.403813,14.56342,15.726933,16.765503,17.804073,18.84655,19.88512,20.92369,20.181856,19.44002,18.698183,17.956347,17.210606,17.850927,18.487345,19.123762,19.764084,20.400501,19.705519,19.010534,18.315552,17.620567,16.925583,14.379913,11.834243,9.288573,6.746807,4.2011366,6.1103897,8.019642,9.928895,11.838148,13.751305,15.621513,17.495626,19.365835,21.239948,23.114061,22.05597,21.00178,19.947592,18.893402,17.839214,17.077856,16.316498,15.559043,14.797685,14.036326,17.917301,21.798277,25.679255,29.556326,33.4373,27.99066,22.544018,17.093473,11.6468315,6.2001905,6.493021,6.785851,7.0786815,7.3715115,7.6643414,11.490656,15.31697,19.143284,22.973503,26.799816,22.700195,18.600573,14.50095,10.401327,6.3017054,12.142691,17.983677,23.828568,29.669552,35.51054,32.285503,29.056562,25.831526,22.602585,19.373644,17.464392,15.555139,13.645885,11.736633,9.823476,11.4398985,13.056321,14.668839,16.285261,17.901684,19.322887,20.74409,22.169195,23.590399,25.0116,24.995983,24.976461,24.960844,24.941322,24.925705,23.668486,22.415173,21.157955,19.904642,18.651329,22.036446,25.421562,28.80668,32.191795,35.576912,32.601757,29.630508,26.659258,23.684105,20.712854,20.693333,20.677715,20.658192,20.642574,20.623053,19.92807,19.229181,18.534197,17.83531,17.136421,13.919194,10.701966,7.4847393,4.267512,1.0502841,8.8083315,16.56638,24.324427,32.078568,39.836617,35.100574,30.360632,25.624592,20.888552,16.148607,14.50095,12.849388,11.20173,9.550168,7.898606,6.4110284,4.9234514,3.435874,1.9482968,0.46071947,1.2415999,2.0224805,2.803361,3.5842414,4.3612175,3.5686235,2.77603,1.9834363,1.1908426,0.39824903,0.40215343,0.40605783,0.40605783,0.40996224,0.41386664,0.95657855,1.4992905,2.0380979,2.5808098,3.1235218,2.7057507,2.2918842,1.8741131,1.456342,1.038571,1.0112402,0.9878138,0.96438736,0.93705654,0.9136301,1.1361811,1.3626363,1.5890918,1.8116426,2.0380979,1.6671798,1.2962615,0.92924774,0.5583295,0.18741131,0.93315214,1.6827974,2.4285383,3.1781836,3.9239242,3.1898966,2.455869,1.7218413,0.98390937,0.24988174,0.3553006,0.46071947,0.5661383,0.6715572,0.77307165,1.0502841,1.3235924,1.6008049,1.8741131,2.1513257,1.7530766,1.358732,0.96438736,0.5700427,0.1756981,0.5309987,0.8862993,1.2415999,1.5969005,1.9482968,1.8584955,1.7686942,1.678893,1.5890918,1.4992905,1.1986516,0.9019169,0.60127795,0.30063897,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.08980125,0.1796025,0.26940376,0.359205,0.44900626,4.2089458,7.968885,11.728825,15.488764,19.248703,15.398962,11.549222,7.699481,3.8497405,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14836729,0.30063897,0.44900626,0.60127795,0.74964523,1.456342,2.1630387,2.87364,3.5803368,4.2870336,3.873167,3.4632049,3.049338,2.639376,2.2255092,1.8038338,1.3782539,0.95657855,0.5349031,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.26940376,0.5388075,0.80821127,1.0815194,1.3509232,1.0815194,0.80821127,0.5388075,0.26940376,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.031235218,0.039044023,0.046852827,0.05466163,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05466163,0.10932326,0.1639849,0.21864653,0.27330816,0.6442264,1.0151446,1.3860629,1.7530766,2.1239948,2.0615244,1.999054,1.9365835,1.8741131,1.8116426,1.5656652,1.3157835,1.0698062,0.8238289,0.57394713,0.5192855,0.46462387,0.40996224,0.3553006,0.30063897,0.27721256,0.25378615,0.23426414,0.21083772,0.18741131,0.16008049,0.13274968,0.10541886,0.078088045,0.05075723,0.19912452,0.3435874,0.49195468,0.64032197,0.78868926,0.71841,0.6481308,0.57785153,0.5075723,0.43729305,0.57394713,0.7106012,0.8511597,0.9878138,1.1244678,1.3626363,1.6008049,1.8389735,2.0732377,2.3114061,2.2918842,2.2684577,2.2450314,2.2216048,2.1981785,1.8741131,1.5500476,1.2259823,0.9019169,0.57394713,0.77307165,0.96829176,1.1674163,1.3665408,1.5617609,2.0380979,2.5183394,2.9946766,3.4710135,3.951255,3.9473507,3.9434462,3.9434462,3.9395418,3.9356375,3.4514916,2.9673457,2.4831998,1.999054,1.5110037,1.3860629,1.261122,1.1361811,1.0112402,0.8862993,0.79259366,0.698888,0.60127795,0.5075723,0.41386664,0.38263142,0.3513962,0.3240654,0.29283017,0.26159495,0.25769055,0.25378615,0.24597734,0.24207294,0.23816854,0.29283017,0.3474918,0.40215343,0.45681506,0.5114767,0.8433509,1.1791295,1.5110037,1.8428779,2.174752,2.3543546,2.5300527,2.7057507,2.8853533,3.0610514,3.7130866,4.3612175,5.0132523,5.661383,6.3134184,7.1021075,7.890797,8.683391,9.47208,10.260769,10.604357,10.947944,11.291532,11.631214,11.974802,12.564366,13.153932,13.743496,14.33306,14.92653,16.199366,17.468296,18.74113,20.013966,21.2868,22.294136,23.301472,24.30881,25.316145,26.32348,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.47633708,0.94876975,1.4251068,1.901444,2.3738766,3.8106966,5.2436123,6.6804323,8.113348,9.550168,9.597021,9.643873,9.690726,9.741484,9.788337,8.531119,7.2739015,6.016684,4.755562,3.4983444,3.2367494,2.97125,2.7057507,2.4402514,2.174752,2.3465457,2.5183394,2.6940374,2.8658314,3.0376248,2.8111696,2.5808098,2.3543546,2.1278992,1.901444,2.5730011,3.2445583,3.9161155,4.591577,5.263134,6.196286,7.125534,8.058686,8.991838,9.924991,9.725866,9.526741,9.323712,9.124588,8.925464,8.4178915,7.910319,7.4027467,6.8951745,6.387602,6.239235,6.0908675,5.9464045,5.7980375,5.64967,5.142098,4.6345253,4.126953,3.619381,3.1118085,3.9942036,4.8765984,5.758993,6.6413884,7.523783,7.996216,8.464745,8.933272,9.405705,9.874233,8.960603,8.050878,7.137247,6.223617,5.3138914,6.3602715,7.406651,8.456935,9.503315,10.549695,10.405232,10.260769,10.116306,9.971844,9.823476,9.440845,9.058213,8.675582,8.296855,7.914223,8.921559,9.928895,10.936231,11.943566,12.950902,13.677121,14.40334,15.133463,15.859682,16.585901,15.855778,15.12175,14.391626,13.657599,12.923572,14.087084,15.250595,16.414106,17.573715,18.737226,20.084246,21.42736,22.774378,24.117493,25.460608,26.81934,28.178072,29.536802,30.89163,32.250362,30.688602,29.130745,27.568985,26.011127,24.449368,25.085785,25.718298,26.354715,26.991133,27.623646,30.548042,33.476345,36.40074,39.325138,42.24954,40.30124,38.349037,36.40074,34.44854,32.500244,30.059994,27.619741,25.179491,22.739239,20.298986,19.783606,19.268225,18.756748,18.241367,17.725986,16.808453,15.890917,14.973383,14.055848,13.138313,13.766922,14.395531,15.028045,15.656653,16.289165,16.628849,16.968533,17.308216,17.647898,17.987581,17.448774,16.91387,16.375063,15.836256,15.3013525,14.821111,14.344774,13.868437,13.388195,12.911859,11.033841,9.155824,7.28171,5.4036927,3.5256753,5.6340523,7.7385254,9.846903,11.955279,14.063657,14.719597,15.375536,16.03538,16.69132,17.351164,16.56638,15.781594,14.996809,14.208119,13.423335,12.853292,12.28325,11.713207,11.143164,10.573121,13.7474,16.921679,20.092054,23.266333,26.436708,22.118439,17.796265,13.477997,9.155824,4.8375545,5.8097506,6.7819467,7.7541428,8.726339,9.698535,12.228588,14.75864,17.288692,19.818747,22.348799,20.37317,18.401447,16.42582,14.450192,12.4745655,20.135002,27.795439,35.455875,43.116314,50.776752,45.158318,39.539883,33.921448,28.303013,22.688482,22.079395,21.474213,20.865126,20.256039,19.650856,19.428307,19.20966,18.991013,18.768461,18.549814,21.130625,23.71534,26.296148,28.880863,31.461674,30.43872,29.415766,28.396717,27.373764,26.350811,26.49137,26.631927,26.768581,26.90914,27.049698,28.834011,30.614418,32.39873,34.17914,35.963448,32.23084,28.498232,24.765623,21.033014,17.300406,17.964155,18.631807,19.295555,19.959305,20.623053,20.431738,20.236517,20.041296,19.846077,19.650856,15.926057,12.205161,8.484266,4.759466,1.038571,8.862993,16.69132,24.519646,32.347973,40.1763,37.626724,35.073246,32.52367,29.974096,27.424522,24.625065,21.82561,19.026152,16.226696,13.423335,10.81129,8.1992445,5.5871997,2.9751544,0.3631094,1.8858263,3.408543,4.93126,6.453977,7.9766936,6.4891167,5.0054436,3.521771,2.0341935,0.5505207,0.5036679,0.46071947,0.41386664,0.3709182,0.3240654,0.74574083,1.1713207,1.5929961,2.0146716,2.436347,2.1161861,1.7921207,1.4680552,1.1478943,0.8238289,0.97610056,1.1244678,1.2767396,1.4251068,1.5734742,1.5890918,1.6008049,1.6125181,1.6242313,1.6359446,1.3470187,1.0580931,0.76916724,0.47633708,0.18741131,0.74574083,1.3040704,1.8584955,2.416825,2.9751544,2.4285383,1.8858263,1.33921,0.79649806,0.24988174,0.46071947,0.6715572,0.8784905,1.0893283,1.3001659,1.3743496,1.4485333,1.5266213,1.6008049,1.6749885,1.397776,1.1205635,0.8433509,0.5661383,0.28892577,0.5583295,0.8316377,1.1049459,1.3782539,1.6515622,1.5461433,1.4407244,1.3353056,1.2298868,1.1244678,0.9019169,0.6754616,0.44900626,0.22645533,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.1796025,0.359205,0.5388075,0.71841,0.9019169,3.6076677,6.3134184,9.023073,11.728825,14.438479,11.549222,8.663869,5.774611,2.8892577,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.113227665,0.22645533,0.3357786,0.44900626,0.5622339,2.0420024,3.5178664,4.9937305,6.473499,7.9493628,6.949836,5.950309,4.950782,3.951255,2.951728,2.4051118,1.8584955,1.3157835,0.76916724,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.49195468,0.98000497,1.4719596,1.9600099,2.4480603,1.9600099,1.4719596,0.98000497,0.48805028,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05466163,0.058566034,0.058566034,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.093705654,0.14055848,0.19131571,0.23816854,0.5270943,0.8160201,1.1088502,1.397776,1.6867018,1.698415,1.7140326,1.7257458,1.737459,1.7491722,1.5539521,1.358732,1.1635119,0.96829176,0.77307165,0.7262188,0.679366,0.63251317,0.58566034,0.5388075,0.46852827,0.39824903,0.3279698,0.25769055,0.18741131,0.1717937,0.15227169,0.13665408,0.11713207,0.10151446,0.21864653,0.339683,0.46071947,0.58175594,0.698888,0.6481308,0.59346914,0.5427119,0.49195468,0.43729305,0.6754616,0.9136301,1.1517987,1.3860629,1.6242313,1.7765031,1.9248703,2.0732377,2.2255092,2.3738766,2.330928,2.2840753,2.241127,2.194274,2.1513257,1.8506867,1.5500476,1.2494087,0.94876975,0.6481308,0.8823949,1.116659,1.3470187,1.5812829,1.8116426,2.3192148,2.822883,3.3265507,3.8341231,4.337791,4.3338866,4.3260775,4.322173,4.318269,4.3143644,3.8302186,3.3460727,2.8658314,2.3816853,1.901444,1.7491722,1.6008049,1.4485333,1.3001659,1.1517987,1.0737107,0.9956226,0.91753453,0.8394465,0.76135844,0.6910792,0.61689556,0.5466163,0.47243267,0.39824903,0.3631094,0.3318742,0.29673457,0.26159495,0.22645533,0.26159495,0.29673457,0.3318742,0.3631094,0.39824903,0.6520352,0.9058213,1.1557031,1.4094892,1.6632754,1.8038338,1.9482968,2.0888553,2.233318,2.3738766,2.951728,3.5256753,4.0996222,4.6735697,5.251421,5.903456,6.559396,7.2153354,7.871275,8.52331,9.136301,9.745388,10.354475,10.963562,11.576552,12.244205,12.911859,13.575606,14.243259,14.9109125,16.093946,17.27698,18.460014,19.643047,20.826082,21.778755,22.73143,23.684105,24.636778,25.585548,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3513962,0.698888,1.0502841,1.4016805,1.7491722,3.1664703,4.579864,5.9932575,7.4105554,8.823949,9.163632,9.503315,9.846903,10.186585,10.526268,9.132397,7.7385254,6.348558,4.9546866,3.5608149,3.3538816,3.1430438,2.9322062,2.7213683,2.514435,2.7526035,2.9907722,3.232845,3.4710135,3.7130866,3.4514916,3.193801,2.9322062,2.6706111,2.4129205,3.1274261,3.8419318,4.5564375,5.270943,5.989353,7.094299,8.1992445,9.304191,10.409137,11.514082,11.248583,10.986988,10.725393,10.4637985,10.198298,9.63216,9.066022,8.495979,7.929841,7.363703,6.9732623,6.5828223,6.192382,5.801942,5.4115014,4.9078336,4.4041657,3.8965936,3.3929255,2.8892577,3.7560349,4.6228123,5.4895897,6.356367,7.223144,7.8673706,8.511597,9.151918,9.796145,10.436467,9.589212,8.738052,7.8868923,7.0357327,6.1884775,6.727285,7.266093,7.8088045,8.347612,8.886419,8.570163,8.253906,7.9337454,7.617489,7.3012323,7.008402,6.715572,6.422742,6.1299114,5.8370814,6.902983,7.9727893,9.0386915,10.108498,11.174399,12.209065,13.243732,14.278399,15.313066,16.351637,16.195461,16.039284,15.883108,15.730837,15.57466,17.27698,18.975395,20.67381,22.37613,24.074545,25.156063,26.233679,27.315199,28.396717,29.474333,29.431385,29.384531,29.341583,29.29473,29.251781,27.373764,25.495747,23.61773,21.739712,19.861694,20.490303,21.118912,21.743616,22.372225,23.000834,28.935526,34.874123,40.812717,46.751312,52.686005,51.225758,49.76161,48.30136,46.837208,45.376965,42.339336,39.30562,36.271896,33.234272,30.200552,29.263494,28.330343,27.393286,26.460135,25.526981,22.5284,19.533724,16.539047,13.544372,10.549695,10.768341,10.990892,11.209538,11.428185,11.650736,13.0719385,14.493141,15.918248,17.33945,18.760653,17.050524,15.336493,13.626364,11.912332,10.198298,9.940608,9.679013,9.421323,9.159728,8.898132,7.6916723,6.481308,5.270943,4.0605783,2.8502135,5.153811,7.461313,9.76491,12.068507,14.376009,13.817679,13.25935,12.70102,12.146595,11.588266,11.072885,10.557504,10.042123,9.526741,9.01136,8.632633,8.253906,7.871275,7.492548,7.113821,9.577498,12.041177,14.508759,16.972437,19.436115,16.246218,13.052417,9.858616,6.6687193,3.474918,5.12648,6.7780423,8.433509,10.085071,11.736633,12.970425,14.204215,15.434102,16.667892,17.901684,18.05005,18.19842,18.35069,18.499058,18.651329,28.127314,37.6033,47.083187,56.55917,66.03906,58.03113,50.0232,42.015274,34.007343,25.999414,26.694399,27.389381,28.084366,28.779348,29.474333,27.420616,25.366901,23.309282,21.255566,19.20185,22.942268,26.68659,30.427008,34.17133,37.911747,35.88536,33.85898,31.828688,29.802303,27.775917,29.310349,30.844778,32.379208,33.91364,35.451973,35.631577,35.811176,35.99078,36.170383,36.349983,31.856018,27.365955,22.871988,18.378021,13.887959,15.234978,16.581997,17.929016,19.276033,20.623053,20.931501,21.239948,21.548395,21.856844,22.161386,17.936825,13.708356,9.479889,5.251421,1.0268579,8.921559,16.820166,24.718771,32.613472,40.512077,40.148968,39.78586,39.426655,39.063545,38.700436,34.74918,30.80183,26.850574,22.899319,18.95197,15.211552,11.475039,7.7385254,3.998108,0.26159495,2.5261483,4.7907014,7.0591593,9.323712,11.588266,9.40961,7.230953,5.056201,2.8775444,0.698888,0.60908675,0.5153811,0.42167544,0.3318742,0.23816854,0.5388075,0.8433509,1.1439898,1.4485333,1.7491722,1.5227169,1.2962615,1.0659018,0.8394465,0.61299115,0.93705654,1.261122,1.5890918,1.9131571,2.2372224,2.0380979,1.8389735,1.6359446,1.43682,1.2376955,1.0268579,0.8160201,0.60908675,0.39824903,0.18741131,0.5544251,0.92143893,1.2884527,1.6593709,2.0263848,1.6710842,1.3157835,0.96048295,0.60518235,0.24988174,0.5661383,0.8784905,1.1947471,1.5110037,1.8233559,1.698415,1.5734742,1.4485333,1.3235924,1.1986516,1.038571,0.8784905,0.71841,0.5583295,0.39824903,0.58956474,0.78088045,0.96829176,1.1596074,1.3509232,1.2298868,1.1088502,0.9917182,0.8706817,0.74964523,0.60127795,0.44900626,0.30063897,0.14836729,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.26940376,0.5388075,0.80821127,1.0815194,1.3509232,3.0063896,4.657952,6.3134184,7.968885,9.6243515,7.699481,5.774611,3.8497405,1.9248703,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,2.6237583,4.8687897,7.1177254,9.366661,11.611692,10.0265045,8.437413,6.8483214,5.263134,3.6740425,3.0063896,2.338737,1.6710842,1.0034313,0.3357786,0.26940376,0.20302892,0.13665408,0.06637484,0.0,0.7106012,1.4212024,2.1318035,2.8385005,3.5491016,2.8385005,2.1318035,1.4212024,0.7106012,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.07418364,0.07027924,0.06637484,0.06637484,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.40996224,0.62079996,0.8316377,1.038571,1.2494087,1.33921,1.4251068,1.5110037,1.6008049,1.6867018,1.5461433,1.4016805,1.261122,1.116659,0.97610056,0.93315214,0.8941081,0.8550641,0.8160201,0.77307165,0.6559396,0.5388075,0.42167544,0.30454338,0.18741131,0.1796025,0.1717937,0.1639849,0.15617609,0.14836729,0.24207294,0.3357786,0.42557985,0.5192855,0.61299115,0.57785153,0.5427119,0.5075723,0.47243267,0.43729305,0.77307165,1.1127546,1.4485333,1.7882162,2.1239948,2.1864653,2.2489357,2.3114061,2.3738766,2.436347,2.3699722,2.3035975,2.233318,2.1669433,2.1005683,1.8233559,1.5500476,1.2767396,0.999527,0.7262188,0.9917182,1.261122,1.5266213,1.796025,2.0615244,2.5964274,3.1274261,3.6584249,4.193328,4.7243266,4.716518,4.7087092,4.7009,4.6930914,4.689187,4.2089458,3.7287042,3.2484627,2.7682211,2.2879796,2.1122816,1.9365835,1.7608855,1.5890918,1.4133936,1.3509232,1.2923572,1.2337911,1.1713207,1.1127546,0.9956226,0.8823949,0.76916724,0.6520352,0.5388075,0.47243267,0.40605783,0.3435874,0.27721256,0.21083772,0.22645533,0.24207294,0.25769055,0.27330816,0.28892577,0.46071947,0.63251317,0.80430686,0.97610056,1.1517987,1.2572175,1.3665408,1.4719596,1.5812829,1.6867018,2.1864653,2.6862288,3.1859922,3.6857557,4.185519,4.7087092,5.2279944,5.74728,6.266566,6.785851,7.6643414,8.542832,9.421323,10.295909,11.174399,11.92014,12.665881,13.411622,14.153459,14.899199,15.992432,17.085665,18.178898,19.268225,20.361458,21.25947,22.157482,23.055496,23.953508,24.85152,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22645533,0.44900626,0.6754616,0.9019169,1.1244678,2.5183394,3.9161155,5.309987,6.703859,8.101635,8.734148,9.366661,9.999174,10.631687,11.2642,9.733675,8.207053,6.6804323,5.153811,3.6232853,3.4710135,3.3148375,3.1586614,3.0063896,2.8502135,3.1586614,3.4632049,3.7716527,4.0801005,4.388548,4.095718,3.802888,3.5100577,3.2172275,2.9243972,3.6818514,4.4393053,5.196759,5.9542136,6.7116675,7.988407,9.269051,10.545791,11.82253,13.09927,12.775204,12.4511385,12.123169,11.799104,11.475039,10.84643,10.221725,9.593117,8.964508,8.335898,7.703386,7.0708723,6.4383593,5.805846,5.173333,4.6735697,4.169902,3.6662338,3.1664703,2.6628022,3.513962,4.369026,5.2201858,6.0713453,6.9264097,7.7385254,8.554545,9.370565,10.186585,10.998701,10.213917,9.425227,8.636538,7.8517528,7.0630636,7.094299,7.1294384,7.1606736,7.191909,7.223144,6.735094,6.2431393,5.755089,5.263134,4.775084,4.572055,4.369026,4.165997,3.9668727,3.7638438,4.8883114,6.016684,7.1450562,8.273428,9.4018,10.741011,12.084125,13.427239,14.770353,16.113468,16.535143,16.95682,17.378494,17.804073,18.22575,20.462973,22.700195,24.937418,27.17464,29.411861,30.227882,31.043901,31.856018,32.67204,33.48806,32.039524,30.590992,29.146362,27.69783,26.249296,24.055023,21.860748,19.666473,17.468296,15.274021,15.894821,16.515621,17.136421,17.753317,18.374117,27.323008,36.275803,45.22469,54.17358,63.126377,62.150276,61.174175,60.201977,59.22588,58.24978,54.618683,50.991493,47.3604,43.729305,40.09821,38.743385,37.388557,36.03373,34.6789,33.324074,28.252254,23.180437,18.108618,13.036799,7.9610763,7.773665,7.5823493,7.3910336,7.2036223,7.012306,9.518932,12.021654,14.528281,17.031002,19.537628,16.64837,13.763018,10.87376,7.988407,5.099149,5.056201,5.0132523,4.9742084,4.93126,4.8883114,4.3455997,3.802888,3.260176,2.717464,2.174752,4.677474,7.180196,9.682918,12.185639,14.688361,12.915763,11.143164,9.370565,7.5979667,5.825368,5.579391,5.3334136,5.0913405,4.845363,4.5993857,4.40807,4.220659,4.029343,3.8380275,3.6506162,5.407597,7.164578,8.921559,10.67854,12.435521,10.373997,8.308568,6.2431393,4.1777105,2.1122816,4.4432096,6.7780423,9.108971,11.443803,13.774731,13.708356,13.645885,13.579511,13.513136,13.450665,15.723028,17.999294,20.27556,22.551826,24.82419,36.119625,47.415062,58.710495,70.005936,81.30137,70.903946,60.506523,50.1091,39.711674,29.314253,31.309402,33.308456,35.303604,37.302658,39.301712,35.409023,31.520239,27.631454,23.738766,19.849981,24.75391,29.653934,34.557865,39.461792,44.36182,41.332,38.298283,35.26456,32.23084,29.201025,32.129326,35.06153,37.989834,40.92204,43.85034,42.42914,41.004032,39.58283,38.16163,36.736523,31.4851,26.233679,20.978354,15.726933,10.475512,12.5058,14.53609,16.56638,18.596668,20.623053,21.43517,22.24338,23.055496,23.863707,24.675823,19.943687,15.211552,10.475512,5.743376,1.0112402,8.980125,16.94901,24.91399,32.882877,40.85176,42.675117,44.498474,46.325733,48.14909,49.97635,44.873295,39.774147,34.674995,29.575848,24.476698,19.611813,14.750832,9.885946,5.024966,0.1639849,3.1703746,6.1767645,9.187058,12.193448,15.199838,12.330102,9.460366,6.590631,3.7208953,0.8511597,0.7106012,0.5700427,0.42948425,0.28892577,0.14836729,0.3318742,0.5153811,0.698888,0.8784905,1.0619974,0.92924774,0.79649806,0.6637484,0.5309987,0.39824903,0.9019169,1.4016805,1.901444,2.4012074,2.900971,2.4871042,2.0732377,1.6632754,1.2494087,0.8355421,0.7066968,0.57785153,0.44900626,0.31625658,0.18741131,0.3631094,0.5427119,0.71841,0.8980125,1.0737107,0.9097257,0.74574083,0.58175594,0.41386664,0.24988174,0.6715572,1.0893283,1.5110037,1.9287747,2.35045,2.0263848,1.698415,1.3743496,1.0502841,0.7262188,0.6832704,0.64032197,0.59737355,0.5544251,0.5114767,0.62079996,0.7262188,0.8355421,0.94096094,1.0502841,0.9136301,0.78088045,0.6442264,0.5114767,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.359205,0.71841,1.0815194,1.4407244,1.7999294,2.4012074,3.0063896,3.6076677,4.2089458,4.814128,3.8497405,2.8892577,1.9248703,0.96438736,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,3.2055142,6.223617,9.24172,12.2559185,15.274021,13.09927,10.924518,8.749765,6.575013,4.4002614,3.611572,2.8189783,2.0302892,1.2415999,0.44900626,0.359205,0.26940376,0.1796025,0.08980125,0.0,0.92924774,1.8584955,2.7916477,3.7208953,4.650143,3.7208953,2.7916477,1.8584955,0.92924774,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.093705654,0.08589685,0.078088045,0.07027924,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.06637484,0.09761006,0.12884527,0.1639849,0.29283017,0.42167544,0.5544251,0.6832704,0.81211567,0.97610056,1.1361811,1.3001659,1.4641509,1.6242313,1.53443,1.4446288,1.3548276,1.2650263,1.175225,1.1439898,1.1088502,1.077615,1.0463798,1.0112402,0.8472553,0.6832704,0.5192855,0.3513962,0.18741131,0.19131571,0.19131571,0.19522011,0.19912452,0.19912452,0.26549935,0.3318742,0.39434463,0.46071947,0.5231899,0.5075723,0.48805028,0.47243267,0.45681506,0.43729305,0.8745861,1.3118792,1.7491722,2.1864653,2.6237583,2.6003318,2.5769055,2.5495746,2.5261483,2.4988174,2.4090161,2.3192148,2.2294137,2.1396124,2.0498111,1.7999294,1.5500476,1.3001659,1.0502841,0.80040246,1.1010414,1.4055848,1.7062237,2.0107672,2.3114061,2.87364,3.4319696,3.9942036,4.552533,5.1108627,5.1030536,5.0913405,5.083532,5.0718184,5.0640097,4.5837684,4.1074314,3.631094,3.1508527,2.6745155,2.475391,2.2762666,2.0732377,1.8741131,1.6749885,1.6320401,1.5890918,1.5461433,1.5031948,1.4641509,1.3040704,1.1478943,0.9917182,0.8316377,0.6754616,0.58175594,0.48414588,0.39044023,0.29673457,0.19912452,0.19522011,0.19131571,0.1835069,0.1796025,0.1756981,0.26940376,0.359205,0.45291066,0.5466163,0.63641757,0.7106012,0.78088045,0.8550641,0.92924774,0.999527,1.4251068,1.8506867,2.2762666,2.7018464,3.1235218,3.5100577,3.8965936,4.279225,4.6657605,5.0483923,6.196286,7.3402762,8.484266,9.628256,10.77615,11.596075,12.419904,13.243732,14.063657,14.8874855,15.890917,16.894348,17.893875,18.897306,19.900738,20.74409,21.583536,22.426888,23.270237,24.113588,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,1.8741131,3.2484627,4.6267166,6.001066,7.375416,8.300759,9.226103,10.151445,11.076789,11.998228,10.338858,8.675582,7.012306,5.349031,3.6857557,3.5881457,3.4866312,3.3890212,3.2875066,3.1859922,3.5608149,3.9356375,4.3143644,4.689187,5.0640097,4.73604,4.4119744,4.087909,3.7638438,3.435874,4.2362766,5.036679,5.8370814,6.6374836,7.437886,8.886419,10.338858,11.787391,13.235924,14.688361,14.301826,13.911386,13.524849,13.138313,12.751778,12.0606985,11.373524,10.686349,9.999174,9.311999,8.437413,7.562827,6.688241,5.813655,4.939069,4.4393053,3.9356375,3.435874,2.9361105,2.436347,3.2757936,4.1113358,4.950782,5.786324,6.6257706,7.6135845,8.601398,9.589212,10.573121,11.560935,10.838621,10.112402,9.386183,8.663869,7.9376497,7.461313,6.98888,6.5125427,6.036206,5.563773,4.900025,4.2362766,3.5764325,2.912684,2.2489357,2.135708,2.0263848,1.9131571,1.7999294,1.6867018,2.87364,4.0605783,5.251421,6.4383593,7.6252975,9.276859,10.924518,12.576079,14.223738,15.875299,16.874826,17.874353,18.87388,19.873407,20.876839,23.648964,26.424995,29.201025,31.97315,34.74918,35.2997,35.85022,36.40074,36.951263,37.501785,34.65157,31.801357,28.951143,26.10093,23.250715,20.73628,18.22575,15.711315,13.200784,10.686349,11.29934,11.912332,12.525322,13.138313,13.751305,25.71049,37.673576,49.636665,61.599754,73.56284,73.07479,72.58674,72.098694,71.61064,71.126495,66.90193,62.673466,58.448902,54.22434,49.999775,48.22327,46.450672,44.67417,42.901573,41.12507,33.97611,26.827148,19.674282,12.525322,5.376362,4.775084,4.173806,3.5764325,2.9751544,2.3738766,5.9620223,9.550168,13.138313,16.72646,20.310701,16.250122,12.189544,8.125061,4.0605783,0.0,0.1756981,0.3513962,0.5231899,0.698888,0.8745861,0.999527,1.1244678,1.2494087,1.3743496,1.4992905,4.2011366,6.899079,9.600925,12.298867,15.000713,12.013845,9.026978,6.036206,3.049338,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,1.2376955,2.2879796,3.338264,4.388548,5.4388323,4.5017757,3.5608149,2.6237583,1.6867018,0.74964523,3.7638438,6.774138,9.788337,12.798631,15.812829,14.450192,13.087557,11.72492,10.362284,8.999647,13.399908,17.800169,22.200432,26.600693,31.000954,44.11194,57.22292,70.33781,83.44879,96.563675,83.77676,70.989845,58.19902,45.4121,32.625187,35.924404,39.223625,42.52675,45.82597,49.12519,43.401337,37.673576,31.949724,26.22587,20.498112,26.56165,32.625187,38.68872,44.748356,50.81189,46.77474,42.737587,38.700436,34.663284,30.626131,34.948303,39.274384,43.60046,47.926537,52.24871,49.226704,46.20079,43.17488,40.148968,37.12306,31.114182,25.101402,19.088623,13.075843,7.0630636,9.776623,12.486279,15.199838,17.913397,20.623053,21.938837,23.250715,24.562595,25.874474,27.186354,21.95055,16.710842,11.475039,6.239235,0.999527,9.0386915,17.073952,25.113115,33.148376,41.18754,45.201263,49.211086,53.22481,57.238537,61.24836,55.001316,48.750366,42.49942,36.24847,30.001427,24.012074,18.026625,12.037272,6.0518236,0.062470436,3.814601,7.562827,11.311053,15.063184,18.81141,15.250595,11.685876,8.125061,4.564246,0.999527,0.81211567,0.62470436,0.43729305,0.24988174,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.37482262,0.3357786,0.30063897,0.26159495,0.22645533,0.18741131,0.8628729,1.5383345,2.2137961,2.8892577,3.5608149,2.9361105,2.3114061,1.6867018,1.0619974,0.43729305,0.38653582,0.3357786,0.28892577,0.23816854,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.14836729,0.1756981,0.19912452,0.22645533,0.24988174,0.77697605,1.3001659,1.8233559,2.35045,2.87364,2.35045,1.8233559,1.3001659,0.77307165,0.24988174,0.3240654,0.39824903,0.47633708,0.5505207,0.62470436,0.6481308,0.6754616,0.698888,0.7262188,0.74964523,0.60127795,0.44900626,0.30063897,0.14836729,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.44900626,0.9019169,1.3509232,1.7999294,2.2489357,1.7999294,1.3509232,0.9019169,0.44900626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.78727,7.57454,11.361811,15.14908,18.936352,16.175938,13.411622,10.651209,7.8868923,5.12648,4.21285,3.2992198,2.3855898,1.475864,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,1.1517987,2.2996929,3.4514916,4.5993857,5.7511845,4.5993857,3.4514916,2.2996929,1.1517987,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.1756981,0.22645533,0.27330816,0.3240654,0.37482262,0.61299115,0.8511597,1.0893283,1.3235924,1.5617609,1.5266213,1.4875772,1.4485333,1.4133936,1.3743496,1.3509232,1.3235924,1.3001659,1.2767396,1.2494087,1.038571,0.8238289,0.61299115,0.39824903,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,0.28892577,0.3240654,0.3631094,0.39824903,0.43729305,0.43729305,0.43729305,0.43729305,0.43729305,0.43729305,0.97610056,1.5110037,2.0498111,2.5886188,3.1235218,3.0141985,2.900971,2.787743,2.6745155,2.5612879,2.4480603,2.338737,2.2255092,2.1122816,1.999054,1.7765031,1.5500476,1.3235924,1.1010414,0.8745861,1.2142692,1.5500476,1.8858263,2.2255092,2.5612879,3.1508527,3.736513,4.3260775,4.911738,5.5013027,5.4856853,5.473972,5.462259,5.4505453,5.4388323,4.9624953,4.4861584,4.0137253,3.5373883,3.0610514,2.8385005,2.612045,2.3855898,2.1630387,1.9365835,1.9131571,1.8858263,1.8623998,1.8389735,1.8116426,1.6125181,1.4133936,1.2142692,1.0112402,0.81211567,0.6871748,0.5622339,0.43729305,0.31235218,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.1639849,0.19912452,0.23816854,0.27330816,0.31235218,0.6637484,1.0112402,1.3626363,1.7140326,2.0615244,2.3114061,2.5612879,2.8111696,3.0610514,3.310933,4.7243266,6.13772,7.551114,8.960603,10.373997,11.275913,12.173926,13.075843,13.973856,14.875772,15.789403,16.69913,17.612759,18.526388,19.436115,20.224804,21.013493,21.798277,22.586967,23.375656,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12884527,0.25378615,0.38263142,0.5114767,0.63641757,1.8897307,3.1430438,4.396357,5.645766,6.899079,7.8634663,8.831758,9.796145,10.760532,11.72492,10.604357,9.483793,8.36323,7.2465706,6.126007,5.903456,5.6809053,5.4583545,5.2358036,5.0132523,5.263134,5.5169206,5.7707067,6.0205884,6.2743745,5.7785153,5.2865605,4.7907014,4.2948427,3.7989833,4.8765984,5.9542136,7.0318284,8.109444,9.187058,10.2881,11.393045,12.494087,13.599033,14.700074,14.294017,13.891863,13.4858055,13.079747,12.67369,12.056794,11.4398985,10.823003,10.206107,9.589212,9.093353,8.597494,8.101635,7.605776,7.113821,6.126007,5.142098,4.1581883,3.174279,2.1864653,2.9868677,3.7833657,4.579864,5.376362,6.1767645,7.28171,8.39056,9.499411,10.604357,11.713207,11.252487,10.791768,10.331048,9.874233,9.413514,8.843472,8.273428,7.703386,7.1333427,6.5633,6.168956,5.7785153,5.3841705,4.9937305,4.5993857,4.8805027,5.165524,5.446641,5.7316628,6.012779,7.348085,8.683391,10.018696,11.354002,12.689307,13.638077,14.590752,15.543426,16.4961,17.448774,17.495626,17.538574,17.585428,17.628376,17.675228,20.06082,22.450314,24.835903,27.225397,29.610987,30.786211,31.957533,33.128853,34.304077,35.4754,34.42121,33.363117,32.30893,31.25474,30.200552,28.080462,25.960371,23.84028,21.72019,19.6001,18.623999,17.643993,16.667892,15.6917925,14.711788,23.805141,32.898495,41.991848,51.081295,60.17465,59.55775,58.940857,58.32396,57.707066,57.086266,54.134537,51.182808,48.231083,45.279354,42.32372,41.25001,40.1763,39.098682,38.024975,36.951263,30.419197,23.891037,17.358973,10.8308115,4.298747,4.029343,3.7599394,3.4905357,3.2211318,2.951728,5.677001,8.406178,11.131451,13.860628,16.585901,13.271063,9.952321,6.6335793,3.3187418,0.0,0.16008049,0.32016098,0.48024148,0.64032197,0.80040246,1.2962615,1.7882162,2.2840753,2.7799344,3.2757936,5.12648,6.9810715,8.831758,10.686349,12.537036,10.131924,7.726812,5.3217,2.9165885,0.5114767,0.44510186,0.37872702,0.30844778,0.24207294,0.1756981,0.1756981,0.1796025,0.1835069,0.1835069,0.18741131,2.979059,5.7707067,8.566258,11.357906,14.149553,11.849861,9.550168,7.250475,4.950782,2.6510892,4.650143,6.649197,8.648251,10.651209,12.650263,12.08803,11.525795,10.963562,10.401327,9.839094,14.30573,18.77627,23.24681,27.717352,32.187893,41.64045,51.093006,60.545567,69.99812,79.45068,69.13915,58.83153,48.520008,38.20848,27.900858,32.016098,36.135242,40.254387,44.36963,48.488773,42.2183,35.951736,29.685171,23.418604,17.148134,22.04035,26.928663,31.820879,36.70919,41.601406,39.30562,37.00983,34.71404,32.41825,30.126368,33.058575,35.994686,38.930794,41.866905,44.79911,42.167545,39.535976,36.90441,34.26894,31.637371,27.580698,23.527927,19.471254,15.418485,11.361811,13.466284,15.570756,17.679134,19.783606,21.888079,21.903696,21.919313,21.931028,21.946646,21.962263,17.964155,13.962143,9.964035,5.9620223,1.9639144,8.574067,15.188125,21.802181,28.412334,35.026394,38.5833,42.140213,45.697124,49.254036,52.810944,47.305737,41.804436,36.29923,30.79402,25.288813,21.884174,18.479536,15.070992,11.666354,8.261715,9.815667,11.373524,12.927476,14.481428,16.039284,13.513136,10.986988,8.460839,5.938596,3.4124475,2.7486992,2.0810463,1.4172981,0.75354964,0.08589685,0.12884527,0.1717937,0.21474212,0.25769055,0.30063897,0.26940376,0.23816854,0.21083772,0.1796025,0.14836729,0.6949836,1.2415999,1.7843118,2.330928,2.87364,2.463678,2.0537157,1.6437533,1.2337911,0.8238289,0.7027924,0.58175594,0.45681506,0.3357786,0.21083772,0.3318742,0.44900626,0.5661383,0.6832704,0.80040246,0.92534333,1.0502841,1.175225,1.3001659,1.4251068,1.8467822,2.2684577,2.6940374,3.1157131,3.5373883,2.893162,2.25284,1.6086137,0.96829176,0.3240654,0.5075723,0.6910792,0.8706817,1.0541886,1.2376955,1.1127546,0.9878138,0.8628729,0.737932,0.61299115,0.49195468,0.3709182,0.25378615,0.13274968,0.011713207,0.20693332,0.40215343,0.59737355,0.79259366,0.9878138,0.8433509,0.7027924,0.5583295,0.41777104,0.27330816,0.31625658,0.3553006,0.39434463,0.43338865,0.47633708,0.41777104,0.359205,0.30063897,0.24597734,0.18741131,0.5114767,0.8316377,1.1557031,1.475864,1.7999294,1.9834363,2.1630387,2.3465457,2.5300527,2.7135596,2.1708477,1.6281357,1.0854238,0.5427119,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,3.1508527,6.153338,9.155824,12.158309,15.160794,12.978233,10.791768,8.609207,6.422742,4.2362766,3.4788225,2.7213683,1.9639144,1.2064602,0.44900626,0.5075723,0.5661383,0.62079996,0.679366,0.737932,1.5734742,2.4090161,3.240654,4.0761957,4.911738,3.951255,2.9907722,2.0341935,1.0737107,0.113227665,0.16008049,0.20693332,0.25378615,0.30063897,0.3513962,0.28111696,0.21474212,0.14836729,0.078088045,0.011713207,0.042948425,0.07418364,0.10151446,0.13274968,0.1639849,0.14055848,0.12103647,0.10151446,0.08199245,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.1717937,0.21474212,0.26159495,0.30454338,0.3513962,0.5388075,0.7301232,0.92143893,1.1088502,1.3001659,1.2767396,1.2533131,1.2337911,1.2103647,1.1869383,1.175225,1.1635119,1.1517987,1.1361811,1.1244678,0.95657855,0.78868926,0.62079996,0.45681506,0.28892577,0.27330816,0.26159495,0.24988174,0.23816854,0.22645533,0.24988174,0.27330816,0.30063897,0.3240654,0.3513962,0.359205,0.3709182,0.37872702,0.39044023,0.39824903,0.8238289,1.2494087,1.6749885,2.1005683,2.5261483,2.4597735,2.3933985,2.330928,2.2645533,2.1981785,2.1239948,2.0459068,1.9678187,1.8897307,1.8116426,1.6086137,1.4055848,1.2064602,1.0034313,0.80040246,1.1244678,1.4485333,1.7765031,2.1005683,2.4246337,2.9361105,3.4514916,3.9629683,4.474445,4.985922,4.939069,4.892216,4.845363,4.7985106,4.7516575,4.322173,3.8965936,3.4671092,3.0415294,2.612045,2.4324427,2.25284,2.0732377,1.893635,1.7140326,1.698415,1.6867018,1.6749885,1.6632754,1.6515622,1.4953861,1.33921,1.1869383,1.0307622,0.8745861,0.77697605,0.679366,0.58175594,0.48414588,0.38653582,0.3553006,0.3240654,0.28892577,0.25769055,0.22645533,0.21474212,0.20693332,0.19522011,0.1835069,0.1756981,0.19522011,0.21474212,0.23426414,0.25378615,0.27330816,0.5544251,0.8355421,1.116659,1.3938715,1.6749885,1.8819219,2.084951,2.2918842,2.494913,2.7018464,3.8575494,5.0132523,6.17286,7.328563,8.488171,9.296382,10.100689,10.9089,11.717112,12.525322,13.528754,14.53609,15.539521,16.546856,17.550287,18.362404,19.174519,19.986635,20.79875,21.610867,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15617609,0.30844778,0.46462387,0.62079996,0.77307165,1.9053483,3.0337205,4.165997,5.2943697,6.426646,7.4300776,8.433509,9.440845,10.444276,11.4516115,10.87376,10.295909,9.718058,9.140205,8.562354,8.218767,7.871275,7.5276875,7.1841,6.8366084,6.969358,7.098203,7.2270484,7.355894,7.4886436,6.8209906,6.1572423,5.493494,4.825841,4.1620927,5.5169206,6.871748,8.226576,9.581403,10.936231,11.693685,12.447234,13.200784,13.958238,14.711788,14.2901125,13.868437,13.446761,13.021181,12.599506,12.05289,11.506273,10.955752,10.409137,9.86252,9.749292,9.63216,9.518932,9.4018,9.288573,7.816613,6.348558,4.8765984,3.408543,1.9365835,2.6940374,3.4514916,4.2089458,4.9663997,5.7238536,6.9537406,8.179723,9.405705,10.6355915,11.861574,11.666354,11.471134,11.275913,11.080693,10.889378,10.221725,9.557977,8.894228,8.226576,7.562827,7.4417906,7.3168497,7.195813,7.0708723,6.949836,7.629202,8.304664,8.98403,9.659492,10.338858,11.818625,13.302299,14.785972,16.26574,17.749413,18.003199,18.26089,18.514675,18.768461,19.026152,18.116426,17.206701,16.29307,15.383345,14.473619,16.476578,18.475632,20.474686,22.47374,24.476698,26.268818,28.064844,29.860868,31.656893,33.449013,34.19085,34.928783,35.67062,36.40855,37.150387,35.42074,33.694992,31.969246,30.239595,28.51385,25.944754,23.37956,20.810465,18.241367,15.676175,21.895887,28.119505,34.34312,40.56674,46.786453,46.04071,45.291065,44.545326,43.79568,43.04994,41.371048,39.688248,38.009357,36.330463,34.65157,34.27675,33.89802,33.523197,33.148376,32.773552,26.866192,20.954927,15.043662,9.136301,3.2250361,3.2836022,3.3460727,3.4046388,3.4632049,3.5256753,5.3919797,7.2582836,9.128492,10.994797,12.861101,10.2881,7.719003,5.1460023,2.5730011,0.0,0.14446288,0.28892577,0.43338865,0.58175594,0.7262188,1.5890918,2.455869,3.3187418,4.185519,5.0483923,6.055728,7.0591593,8.066495,9.069926,10.073358,8.253906,6.4305506,4.607195,2.7838387,0.96438736,0.80430686,0.6442264,0.48414588,0.3240654,0.1639849,0.1678893,0.1717937,0.1756981,0.1835069,0.18741131,4.7243266,9.257338,13.794253,18.327265,22.86418,19.20185,15.539521,11.873287,8.210958,4.548629,5.5364423,6.524256,7.5120697,8.499884,9.487698,9.725866,9.964035,10.198298,10.436467,10.674636,15.215456,19.756275,24.297094,28.834011,33.374832,39.168964,44.95919,50.753326,56.543552,62.337685,54.505455,46.673225,38.840992,31.008762,23.176533,28.111696,33.042957,37.982025,42.913284,47.84845,41.039173,34.229893,27.420616,20.61134,13.798158,17.519053,21.236044,24.953035,28.670025,32.387016,31.836496,31.28207,30.73155,30.177126,29.626604,31.168842,32.714985,34.26113,35.803368,37.34951,35.108383,32.871162,30.630035,28.388908,26.151686,24.051117,21.954454,19.85779,17.761126,15.664462,17.159847,18.659138,20.154524,21.653814,23.1492,21.868557,20.58401,19.303364,18.018816,16.738173,13.973856,11.213444,8.449126,5.688714,2.9243972,8.113348,13.298394,18.487345,23.676296,28.861341,31.965342,35.065437,38.169437,41.273438,44.37353,39.614067,34.8546,30.095133,25.335667,20.5762,19.75237,18.928543,18.108618,17.284788,16.46096,15.820638,15.18422,14.543899,13.903577,13.263254,11.775677,10.2881,8.800523,7.3129454,5.825368,4.6813784,3.541293,2.397303,1.2533131,0.113227665,0.13665408,0.15617609,0.1796025,0.20302892,0.22645533,0.20302892,0.1796025,0.15617609,0.13665408,0.113227665,0.5270943,0.94096094,1.358732,1.7725986,2.1864653,1.9912452,1.796025,1.6008049,1.4055848,1.2142692,1.0190489,0.8238289,0.62860876,0.43338865,0.23816854,0.48414588,0.7340276,0.98000497,1.2259823,1.475864,1.698415,1.9248703,2.1513257,2.3738766,2.6003318,2.920493,3.240654,3.5608149,3.8809757,4.2011366,3.4397783,2.67842,1.9209659,1.1596074,0.39824903,0.6910792,0.98000497,1.2689307,1.5617609,1.8506867,1.5734742,1.3001659,1.0268579,0.74964523,0.47633708,0.38653582,0.29673457,0.20693332,0.113227665,0.023426414,0.41386664,0.80430686,1.1947471,1.5851873,1.9756275,1.639849,1.3040704,0.96829176,0.63641757,0.30063897,0.42948425,0.5583295,0.6910792,0.8199245,0.94876975,0.8355421,0.71841,0.60518235,0.48805028,0.37482262,0.5700427,0.76526284,0.96048295,1.1557031,1.3509232,2.1669433,2.979059,3.795079,4.6110992,5.423215,4.3416953,3.2562714,2.1708477,1.0854238,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,2.5183394,4.73604,6.9537406,9.171441,11.389141,9.780528,8.171914,6.5633,4.958591,3.349977,2.7486992,2.1435168,1.542239,0.94096094,0.3357786,0.5661383,0.79259366,1.0190489,1.2494087,1.475864,1.9951496,2.514435,3.0337205,3.5569105,4.0761957,3.3031244,2.533957,1.7647898,0.9956226,0.22645533,0.32016098,0.41386664,0.5114767,0.60518235,0.698888,0.5661383,0.42948425,0.29673457,0.16008049,0.023426414,0.058566034,0.093705654,0.12884527,0.1639849,0.19912452,0.1717937,0.14446288,0.11713207,0.08980125,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.1639849,0.20693332,0.24597734,0.28502136,0.3240654,0.46852827,0.60908675,0.75354964,0.8941081,1.038571,1.0307622,1.0229534,1.0151446,1.0073358,0.999527,0.999527,0.999527,0.999527,0.999527,0.999527,0.8784905,0.75354964,0.63251317,0.5114767,0.38653582,0.3513962,0.31235218,0.27330816,0.23816854,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,0.26159495,0.28111696,0.30063897,0.3240654,0.3435874,0.3631094,0.6754616,0.9878138,1.3001659,1.6125181,1.9248703,1.9092526,1.8897307,1.8741131,1.8545911,1.8389735,1.796025,1.7530766,1.7101282,1.6671798,1.6242313,1.4446288,1.2650263,1.0854238,0.9058213,0.7262188,1.038571,1.3509232,1.6632754,1.9756275,2.2879796,2.7252727,3.1625657,3.5998588,4.037152,4.474445,4.3924527,4.31046,4.2284675,4.1464753,4.0605783,3.6818514,3.3031244,2.9243972,2.541766,2.1630387,2.0263848,1.893635,1.756981,1.6242313,1.4875772,1.4875772,1.4875772,1.4875772,1.4875772,1.4875772,1.3782539,1.2689307,1.1557031,1.0463798,0.93705654,0.8667773,0.79649806,0.7262188,0.6559396,0.58566034,0.5466163,0.5075723,0.46852827,0.42557985,0.38653582,0.3553006,0.3240654,0.28892577,0.25769055,0.22645533,0.22645533,0.23035973,0.23426414,0.23426414,0.23816854,0.44900626,0.6559396,0.8667773,1.077615,1.2884527,1.4485333,1.6086137,1.7686942,1.9287747,2.0888553,2.9907722,3.892689,4.794606,5.6965227,6.5984397,7.3168497,8.031356,8.745861,9.460366,10.174872,11.272009,12.369146,13.466284,14.56342,15.660558,16.500004,17.33945,18.174992,19.010534,19.849981,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1835069,0.3631094,0.5466163,0.7301232,0.9136301,1.9209659,2.9283018,3.9356375,4.942973,5.950309,6.996689,8.039165,9.085544,10.131924,11.174399,11.139259,11.10412,11.06898,11.033841,10.998701,10.534078,10.065549,9.597021,9.128492,8.663869,8.671678,8.679486,8.683391,8.691199,8.699008,7.8634663,7.0318284,6.196286,5.3607445,4.5252023,6.1572423,7.7892823,9.421323,11.053363,12.689307,13.095366,13.501423,13.911386,14.317443,14.723501,14.286208,13.845011,13.403813,12.96652,12.525322,12.0489855,11.568744,11.092407,10.61607,10.135828,10.401327,10.666827,10.932326,11.197825,11.4633255,9.507219,7.551114,5.5989127,3.6428072,1.6867018,2.4051118,3.1235218,3.8419318,4.5564375,5.2748475,6.621866,7.968885,9.315904,10.666827,12.013845,12.084125,12.154405,12.220779,12.291059,12.361338,11.603884,10.8425255,10.081166,9.323712,8.562354,8.710721,8.859089,9.0035515,9.151918,9.300286,10.373997,11.443803,12.517513,13.591225,14.661031,16.29307,17.921206,19.553246,21.181383,22.813423,22.36832,21.927124,21.485926,21.040823,20.599627,18.733322,16.870922,15.004618,13.138313,11.275913,12.888432,14.50095,16.113468,17.725986,19.338505,21.75533,24.172153,26.58898,29.005804,31.426535,33.96049,36.49445,39.028404,41.566265,44.100224,42.76492,41.42961,40.094307,38.759003,37.423695,33.269413,29.111223,24.953035,20.794846,16.636658,19.99054,23.340517,26.694399,30.048279,33.39826,32.52367,31.64518,30.76669,29.888199,29.013613,28.603651,28.197594,27.791534,27.381573,26.975515,27.29958,27.623646,27.951616,28.27568,28.599747,23.309282,18.018816,12.728352,7.4417906,2.1513257,2.541766,2.9283018,3.3187418,3.7091823,4.0996222,5.1069584,6.114294,7.1216297,8.128965,9.136301,7.309041,5.481781,3.6545205,1.8272603,0.0,0.12884527,0.26159495,0.39044023,0.5192855,0.6481308,1.8858263,3.1196175,4.3534083,5.591104,6.824895,6.9810715,7.141152,7.297328,7.453504,7.6135845,6.3719845,5.134289,3.892689,2.6510892,1.4133936,1.1596074,0.9058213,0.6559396,0.40215343,0.14836729,0.15617609,0.1639849,0.1717937,0.1796025,0.18741131,6.46569,12.743969,19.022247,25.296621,31.574902,26.549934,21.52497,16.500004,11.475039,6.4500723,6.426646,6.3993154,6.375889,6.348558,6.3251314,7.363703,8.398369,9.43694,10.475512,11.514082,16.121277,20.732376,25.343475,29.95067,34.561768,36.693573,38.825375,40.961082,43.092888,45.22469,39.86785,34.514915,29.158075,23.805141,18.448301,24.20339,29.954575,35.705757,41.460846,47.212032,39.860043,32.508053,25.156063,17.804073,10.44818,12.993851,15.539521,18.085192,20.630861,23.176533,24.36347,25.554314,26.745155,27.935999,29.12684,29.279112,29.43529,29.591465,29.743736,29.899912,28.053131,26.206348,24.355661,22.508879,20.662096,20.521538,20.38098,20.244326,20.103767,19.96321,20.853413,21.743616,22.63382,23.524023,24.414227,21.833418,19.252607,16.671797,14.090988,11.514082,9.987461,8.460839,6.9381227,5.4115014,3.8887846,7.648724,11.412568,15.176412,18.936352,22.700195,25.34738,27.994564,30.641748,33.288933,35.93612,31.922394,27.908667,23.891037,19.877312,15.863586,17.624472,19.381453,21.142338,22.903223,24.664108,21.82561,18.991013,16.156416,13.32182,10.487225,10.0382185,9.589212,9.136301,8.687295,8.238289,6.617962,4.997635,3.377308,1.756981,0.13665408,0.14055848,0.14055848,0.14446288,0.14836729,0.14836729,0.13665408,0.12103647,0.10541886,0.08980125,0.07418364,0.359205,0.6442264,0.92924774,1.2142692,1.4992905,1.5188124,1.5383345,1.5617609,1.5812829,1.6008049,1.3314011,1.0659018,0.79649806,0.5309987,0.26159495,0.64032197,1.0190489,1.3938715,1.7725986,2.1513257,2.475391,2.7994564,3.1235218,3.4514916,3.775557,3.9942036,4.2089458,4.4275923,4.646239,4.860981,3.9863946,3.1079042,2.2294137,1.3509232,0.47633708,0.8706817,1.2689307,1.6671798,2.0654287,2.463678,2.0380979,1.6125181,1.1869383,0.76135844,0.3357786,0.27721256,0.21864653,0.15617609,0.09761006,0.039044023,0.62079996,1.2064602,1.7921207,2.377781,2.9634414,2.436347,1.9092526,1.3782539,0.8511597,0.3240654,0.5466163,0.76526284,0.98390937,1.2064602,1.4251068,1.2533131,1.0815194,0.9058213,0.7340276,0.5622339,0.62860876,0.698888,0.76526284,0.8316377,0.9019169,2.3465457,3.795079,5.2436123,6.688241,8.136774,6.5086384,4.884407,3.2562714,1.6281357,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08980125,0.1796025,0.26940376,0.359205,0.44900626,1.8819219,3.3148375,4.747753,6.180669,7.6135845,6.5828223,5.55206,4.521298,3.4905357,2.463678,2.0146716,1.5656652,1.1205635,0.6715572,0.22645533,0.62079996,1.0190489,1.4172981,1.815547,2.2137961,2.416825,2.6237583,2.8267872,3.0337205,3.2367494,2.6588979,2.077142,1.4992905,0.91753453,0.3357786,0.48024148,0.62079996,0.76526284,0.9058213,1.0502841,0.8472553,0.6442264,0.44119745,0.23816854,0.039044023,0.078088045,0.11713207,0.15617609,0.19912452,0.23816854,0.20302892,0.1678893,0.13274968,0.09761006,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.16008049,0.19522011,0.23035973,0.26549935,0.30063897,0.39434463,0.48805028,0.58566034,0.679366,0.77307165,0.78088045,0.78868926,0.79649806,0.80430686,0.81211567,0.8238289,0.8394465,0.8511597,0.8628729,0.8745861,0.79649806,0.71841,0.6442264,0.5661383,0.48805028,0.42557985,0.3631094,0.30063897,0.23816854,0.1756981,0.1756981,0.1756981,0.1756981,0.1756981,0.1756981,0.20693332,0.23426414,0.26549935,0.29673457,0.3240654,0.5231899,0.7262188,0.92534333,1.1244678,1.3235924,1.3548276,1.3860629,1.4133936,1.4446288,1.475864,1.4680552,1.4602464,1.4524376,1.4446288,1.43682,1.2806439,1.1205635,0.96438736,0.80821127,0.6481308,0.94876975,1.2494087,1.5500476,1.8506867,2.1513257,2.514435,2.87364,3.2367494,3.5998588,3.9629683,3.8458362,3.7287042,3.611572,3.4905357,3.3734035,3.0415294,2.7096553,2.377781,2.0459068,1.7140326,1.6242313,1.53443,1.4407244,1.3509232,1.261122,1.2767396,1.2884527,1.3001659,1.3118792,1.3235924,1.261122,1.1947471,1.1283722,1.0659018,0.999527,0.95657855,0.9136301,0.8706817,0.8316377,0.78868926,0.7418364,0.6910792,0.6442264,0.59737355,0.5505207,0.4958591,0.44119745,0.38653582,0.3318742,0.27330816,0.26159495,0.24597734,0.23035973,0.21474212,0.19912452,0.339683,0.48024148,0.62079996,0.76135844,0.9019169,1.0151446,1.1283722,1.2455044,1.358732,1.475864,2.1239948,2.7682211,3.416352,4.0644827,4.7126136,5.3334136,5.958118,6.578918,7.2036223,7.824422,9.0152645,10.206107,11.393045,12.583888,13.774731,14.637604,15.500477,16.36335,17.226223,18.089096,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21083772,0.42167544,0.62860876,0.8394465,1.0502841,1.9365835,2.8189783,3.7052777,4.591577,5.473972,6.559396,7.6448197,8.730244,9.815667,10.901091,11.408664,11.916236,12.423808,12.93138,13.438952,12.849388,12.2559185,11.666354,11.076789,10.487225,10.373997,10.256865,10.143637,10.0265045,9.913278,8.905942,7.90251,6.899079,5.891743,4.8883114,6.7975645,8.706817,10.61607,12.529227,14.438479,14.4970455,14.555612,14.618082,14.676648,14.739119,14.278399,13.821584,13.364769,12.907954,12.4511385,12.041177,11.6351185,11.229061,10.819098,10.413041,11.057267,11.701493,12.34572,12.993851,13.638077,11.197825,8.757574,6.3173227,3.8770714,1.43682,2.1161861,2.7916477,3.4710135,4.1464753,4.825841,6.2938967,7.758047,9.226103,10.694158,12.162213,12.497992,12.83377,13.165645,13.501423,13.837202,12.982138,12.127073,11.272009,10.416945,9.561881,9.979652,10.397423,10.815194,11.232965,11.650736,13.118792,14.586847,16.050997,17.519053,18.987108,20.76361,22.544018,24.320522,26.097025,27.873528,26.733442,25.593357,24.453272,23.313187,22.1731,19.354122,16.535143,13.716166,10.893282,8.074304,9.300286,10.526268,11.748346,12.974329,14.200311,17.237936,20.279465,23.320995,26.35862,29.400148,33.73013,38.060112,42.390095,46.720078,51.05006,50.1091,49.164234,48.22327,47.278408,46.337444,40.590164,34.842884,29.095606,23.348326,17.601046,18.081287,18.565434,19.045673,19.52982,20.013966,19.00663,17.99539,16.988054,15.980719,14.973383,15.84016,16.703033,17.56981,18.436588,19.29946,20.326319,21.349272,22.37613,23.399082,24.425941,19.756275,15.086611,10.413041,5.743376,1.0737107,1.796025,2.514435,3.2367494,3.9551594,4.6735697,4.8219366,4.970304,5.1186714,5.263134,5.4115014,4.3299823,3.2484627,2.1630387,1.0815194,0.0,0.113227665,0.23035973,0.3435874,0.46071947,0.57394713,2.1786566,3.7833657,5.3919797,6.996689,8.601398,7.910319,7.2192397,6.5281606,5.840986,5.1499066,4.493967,3.8341231,3.1781836,2.5183394,1.8623998,1.5188124,1.1713207,0.8277333,0.48414588,0.13665408,0.14836729,0.15617609,0.1678893,0.1756981,0.18741131,8.207053,16.226696,24.246338,32.26598,40.289528,33.901924,27.514322,21.12672,14.739119,8.351517,7.3129454,6.2743745,5.2358036,4.2011366,3.1625657,5.001539,6.8366084,8.675582,10.510651,12.349625,17.031002,21.708477,26.389854,31.071234,35.748707,34.222084,32.695465,31.168842,29.638317,28.111696,25.234152,22.356607,19.479063,16.601519,13.723974,20.295082,26.866192,33.433395,40.004505,46.575615,38.680912,30.786211,22.89151,14.992905,7.098203,8.472553,9.8429985,11.217348,12.591698,13.962143,16.894348,19.826555,22.75876,25.690968,28.623173,27.389381,26.15559,24.921799,23.684105,22.450314,20.99397,19.541533,18.085192,16.628849,15.176412,16.991959,18.81141,20.626957,22.44641,24.261955,24.546976,24.828094,25.109211,25.394232,25.67535,21.798277,17.921206,14.044135,10.163159,6.2860875,6.001066,5.7121406,5.423215,5.138193,4.8492675,7.1880045,9.526741,11.861574,14.200311,16.539047,18.729418,20.92369,23.114061,25.308336,27.498705,24.23072,20.958832,17.690847,14.418958,11.150972,15.492668,19.834364,24.17606,28.521658,32.863354,27.83058,22.801708,17.772839,12.743969,7.7111945,8.300759,8.886419,9.475985,10.061645,10.651209,8.550641,6.453977,4.357313,2.260649,0.1639849,0.14446288,0.12884527,0.10932326,0.093705654,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.19131571,0.3474918,0.5036679,0.6559396,0.81211567,1.0463798,1.2806439,1.5188124,1.7530766,1.9873407,1.6476578,1.3079748,0.96829176,0.62860876,0.28892577,0.79649806,1.3040704,1.8116426,2.3192148,2.8267872,3.2484627,3.6740425,4.0996222,4.5252023,4.950782,5.0640097,5.181142,5.2943697,5.4115014,5.5247293,4.5291066,3.533484,2.541766,1.5461433,0.5505207,1.0541886,1.5617609,2.0654287,2.5690966,3.076669,2.4988174,1.9248703,1.3509232,0.77307165,0.19912452,0.1717937,0.14055848,0.10932326,0.078088045,0.05075723,0.8316377,1.6086137,2.3894942,3.1703746,3.951255,3.2289407,2.5105307,1.7882162,1.0698062,0.3513962,0.659844,0.96829176,1.2806439,1.5890918,1.901444,1.6710842,1.4407244,1.2103647,0.98000497,0.74964523,0.6910792,0.62860876,0.5700427,0.5114767,0.44900626,2.5300527,4.6110992,6.688241,8.769287,10.850334,8.679486,6.5086384,4.3416953,2.1708477,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12103647,0.23816854,0.359205,0.48024148,0.60127795,1.2494087,1.893635,2.541766,3.1898966,3.8380275,3.3851168,2.9322062,2.4792955,2.0263848,1.5734742,1.2806439,0.9917182,0.698888,0.40605783,0.113227665,0.679366,1.2494087,1.815547,2.3816853,2.951728,2.8385005,2.7291772,2.619854,2.5105307,2.4012074,2.0107672,1.620327,1.2298868,0.8394465,0.44900626,0.64032197,0.8316377,1.0190489,1.2103647,1.4016805,1.1283722,0.8589685,0.58956474,0.32016098,0.05075723,0.093705654,0.14055848,0.1835069,0.23035973,0.27330816,0.23426414,0.19131571,0.14836729,0.10541886,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.15617609,0.1835069,0.21474212,0.24597734,0.27330816,0.3240654,0.3709182,0.41777104,0.46462387,0.5114767,0.5349031,0.5583295,0.58175594,0.60127795,0.62470436,0.6481308,0.6754616,0.698888,0.7262188,0.74964523,0.71841,0.6832704,0.6520352,0.62079996,0.58566034,0.4997635,0.41386664,0.3240654,0.23816854,0.14836729,0.13665408,0.12494087,0.113227665,0.10151446,0.08589685,0.12884527,0.1678893,0.20693332,0.24597734,0.28892577,0.37482262,0.46071947,0.5505207,0.63641757,0.7262188,0.80430686,0.8784905,0.95657855,1.0346665,1.1127546,1.1400855,1.1674163,1.1947471,1.2220778,1.2494087,1.116659,0.98000497,0.8433509,0.7106012,0.57394713,0.8628729,1.1517987,1.43682,1.7257458,2.0107672,2.2996929,2.5886188,2.87364,3.1625657,3.4514916,3.2992198,3.1430438,2.9907722,2.8385005,2.6862288,2.4012074,2.1161861,1.8311646,1.5461433,1.261122,1.2181735,1.1713207,1.1283722,1.0815194,1.038571,1.0619974,1.0893283,1.1127546,1.1361811,1.1635119,1.1439898,1.1205635,1.1010414,1.0815194,1.0619974,1.0463798,1.0307622,1.0190489,1.0034313,0.9878138,0.93315214,0.8784905,0.8238289,0.76916724,0.7106012,0.63641757,0.5583295,0.48024148,0.40215343,0.3240654,0.29283017,0.26159495,0.22645533,0.19522011,0.1639849,0.23426414,0.30063897,0.3709182,0.44119745,0.5114767,0.58175594,0.6520352,0.7223144,0.79259366,0.8628729,1.2533131,1.6476578,2.0380979,2.4324427,2.8267872,3.3538816,3.8848803,4.415879,4.9468775,5.473972,6.75852,8.039165,9.323712,10.604357,11.888905,12.775204,13.661504,14.551707,15.438006,16.324306,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23816854,0.47633708,0.7106012,0.94876975,1.1869383,1.9482968,2.7135596,3.474918,4.2362766,5.001539,6.126007,7.250475,8.374943,9.499411,10.6238785,11.674163,12.724447,13.774731,14.825015,15.875299,15.160794,14.450192,13.735687,13.025085,12.31058,12.076316,11.838148,11.599979,11.361811,11.123642,9.948417,8.773191,7.601871,6.426646,5.251421,7.437886,9.6243515,11.810817,14.001186,16.187653,15.8987255,15.613705,15.324779,15.035853,14.750832,14.274494,13.798158,13.325725,12.849388,12.373051,12.037272,11.701493,11.361811,11.0260315,10.686349,11.713207,12.73616,13.763018,14.785972,15.812829,12.888432,9.964035,7.0357327,4.1113358,1.1869383,1.8233559,2.463678,3.1000953,3.736513,4.376835,5.9620223,7.551114,9.136301,10.725393,12.31058,12.911859,13.513136,14.114414,14.711788,15.313066,14.364296,13.411622,12.4628525,11.514082,10.561408,11.248583,11.935758,12.626837,13.314012,14.001186,15.863586,17.725986,19.588387,21.450787,23.313187,25.238056,27.162926,29.087797,31.012667,32.93754,31.098564,29.263494,27.424522,25.585548,23.750479,19.974922,16.199366,12.423808,8.648251,4.8765984,5.7121406,6.551587,7.387129,8.226576,9.062118,12.724447,16.386776,20.049105,23.711435,27.373764,33.49977,39.62578,45.751785,51.87389,57.999897,57.449375,56.898853,56.348335,55.801716,55.251198,47.91092,40.574547,33.23818,25.901804,18.56153,16.175938,13.786445,11.400854,9.01136,6.6257706,5.4856853,4.349504,3.213323,2.0732377,0.93705654,3.076669,5.212377,7.3519893,9.487698,11.623405,13.349152,15.074897,16.800642,18.526388,20.24823,16.199366,12.150499,8.101635,4.0488653,0.0,1.0502841,2.1005683,3.1508527,4.2011366,5.251421,4.5369153,3.8263142,3.1118085,2.4012074,1.6867018,1.3509232,1.0112402,0.6754616,0.3357786,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,2.475391,4.4510183,6.426646,8.398369,10.373997,8.835662,7.3012323,5.7628975,4.224563,2.6862288,2.612045,2.5378613,2.463678,2.3855898,2.3114061,1.8741131,1.43682,0.999527,0.5622339,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,9.948417,19.713327,29.474333,39.239243,49.000248,41.25001,33.49977,25.749533,17.999294,10.249056,8.1992445,6.1494336,4.0996222,2.0498111,0.0,2.639376,5.2748475,7.914223,10.549695,13.189071,17.936825,22.688482,27.436235,32.187893,36.935646,31.750599,26.56165,21.376602,16.187653,10.998701,10.600452,10.198298,9.80005,9.4018,8.999647,16.386776,23.773905,31.161034,38.548164,45.939198,37.501785,29.064371,20.623053,12.185639,3.7482262,3.951255,4.1503797,4.349504,4.548629,4.7516575,9.425227,14.098797,18.77627,23.44984,28.12341,25.499651,22.875893,20.24823,17.624472,15.000713,13.938716,12.8767185,11.810817,10.748819,9.686822,13.462379,17.237936,21.013493,24.78905,28.560703,28.236637,27.91257,27.588507,27.26444,26.936472,21.763138,16.585901,11.412568,6.239235,1.0619974,2.0107672,2.9634414,3.912211,4.860981,5.813655,6.7233806,7.6370106,8.550641,9.464272,10.373997,12.111456,13.848915,15.586374,17.323833,19.061293,16.539047,14.012899,11.486752,8.960603,6.4383593,13.364769,20.287273,27.213684,34.13619,41.0626,33.83555,26.612406,19.385357,12.162213,4.939069,6.5633,8.187531,9.811763,11.435994,13.06413,10.487225,7.914223,5.337318,2.7643168,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.57394713,1.0268579,1.475864,1.9248703,2.3738766,1.9639144,1.5500476,1.1361811,0.7262188,0.31235218,0.94876975,1.5890918,2.2255092,2.8619268,3.4983444,4.025439,4.548629,5.0757227,5.5989127,6.126007,6.13772,6.1494336,6.1611466,6.1767645,6.1884775,5.0757227,3.9629683,2.8502135,1.737459,0.62470436,1.2376955,1.8506867,2.463678,3.076669,3.6857557,2.9634414,2.2372224,1.5110037,0.78868926,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,1.038571,2.0107672,2.9868677,3.9629683,4.939069,4.025439,3.1118085,2.1981785,1.2884527,0.37482262,0.77697605,1.175225,1.5734742,1.9756275,2.3738766,2.0888553,1.7999294,1.5110037,1.2259823,0.93705654,0.74964523,0.5622339,0.37482262,0.18741131,0.0,2.7135596,5.423215,8.136774,10.850334,13.563893,10.850334,8.136774,5.423215,2.7135596,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14836729,0.30063897,0.44900626,0.60127795,0.74964523,0.61299115,0.47633708,0.3357786,0.19912452,0.062470436,0.18741131,0.31235218,0.43729305,0.5622339,0.6871748,0.5505207,0.41386664,0.27330816,0.13665408,0.0,0.737932,1.475864,2.2137961,2.951728,3.6857557,3.2640803,2.8385005,2.4129205,1.9873407,1.5617609,1.3626363,1.1635119,0.96438736,0.76135844,0.5622339,0.80040246,1.038571,1.2767396,1.5110037,1.7491722,1.4133936,1.0737107,0.737932,0.39824903,0.062470436,0.113227665,0.1639849,0.21083772,0.26159495,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.1756981,0.19912452,0.22645533,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.28892577,0.3240654,0.3631094,0.39824903,0.43729305,0.47633708,0.5114767,0.5505207,0.58566034,0.62470436,0.63641757,0.6481308,0.6637484,0.6754616,0.6871748,0.57394713,0.46071947,0.3513962,0.23816854,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.22645533,0.19912452,0.1756981,0.14836729,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,0.74964523,0.81211567,0.8745861,0.93705654,0.999527,1.0619974,0.94876975,0.8394465,0.7262188,0.61299115,0.4997635,0.77307165,1.0502841,1.3235924,1.6008049,1.8741131,2.0888553,2.2996929,2.514435,2.7252727,2.9361105,2.7486992,2.5612879,2.3738766,2.1864653,1.999054,1.7608855,1.5266213,1.2884527,1.0502841,0.81211567,0.81211567,0.81211567,0.81211567,0.81211567,0.81211567,0.8511597,0.8862993,0.92534333,0.96438736,0.999527,1.0268579,1.0502841,1.0737107,1.1010414,1.1244678,1.1361811,1.1517987,1.1635119,1.175225,1.1869383,1.1244678,1.0619974,0.999527,0.93705654,0.8745861,0.77307165,0.6754616,0.57394713,0.47633708,0.37482262,0.3240654,0.27330816,0.22645533,0.1756981,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.14836729,0.1756981,0.19912452,0.22645533,0.24988174,0.38653582,0.5231899,0.6637484,0.80040246,0.93705654,1.3743496,1.8116426,2.2489357,2.6862288,3.1235218,4.5017757,5.8761253,7.250475,8.624825,9.999174,10.912805,11.826434,12.73616,13.64979,14.56342,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19912452,0.39434463,0.59346914,0.78868926,0.9878138,1.815547,2.6432803,3.4710135,4.298747,5.12648,6.3173227,7.5081654,8.702912,9.893755,11.088503,12.455043,13.821584,15.188125,16.55857,17.92511,17.30431,16.679607,16.058807,15.434102,14.813302,14.469715,14.126127,13.786445,13.442857,13.09927,12.041177,10.983084,9.928895,8.870802,7.812709,9.499411,11.186112,12.8767185,14.56342,16.250122,15.74255,15.234978,14.727406,14.219833,13.712261,13.271063,12.825961,12.384764,11.943566,11.498465,11.935758,12.373051,12.814248,13.251541,13.688834,14.821111,15.957292,17.093473,18.22575,19.36193,16.226696,13.087557,9.948417,6.813182,3.6740425,5.805846,7.941554,10.073358,12.205161,14.336966,15.711315,17.08176,18.45611,19.826555,21.200905,21.891983,22.583063,23.278046,23.969126,24.664108,23.86761,23.071114,22.278519,21.482021,20.685524,20.634766,20.58401,20.529346,20.47859,20.423927,20.83389,21.243853,21.653814,22.063778,22.47374,23.820759,25.163872,26.510891,27.854006,29.201025,27.96333,26.725634,25.487938,24.250242,23.012547,19.959305,16.906061,13.856724,10.803481,7.7502384,7.984503,8.218767,8.456935,8.691199,8.925464,11.6351185,14.344774,17.054428,19.764084,22.47374,27.276154,32.074665,36.87708,41.67559,46.4741,46.688843,46.89968,47.11442,47.32526,47.5361,41.121166,34.70623,28.291298,21.876366,15.461433,14.399435,13.333533,12.267632,11.20173,10.135828,9.511124,8.886419,8.261715,7.6370106,7.012306,7.4886436,7.968885,8.445222,8.921559,9.4018,11.810817,14.223738,16.636658,19.049578,21.4625,17.17156,12.8767185,8.58578,4.290938,0.0,0.8862993,1.7686942,2.6549935,3.541293,4.423688,3.8809757,3.3343596,2.7916477,2.2450314,1.698415,1.3626363,1.0268579,0.6871748,0.3513962,0.011713207,0.23426414,0.45291066,0.6715572,0.8941081,1.1127546,2.6432803,4.173806,5.704332,7.230953,8.761478,7.9259367,7.094299,6.2587566,5.423215,4.5876727,4.21285,3.8380275,3.4632049,3.0883822,2.7135596,4.041056,5.3724575,6.703859,8.031356,9.362757,7.523783,5.688714,3.8497405,2.0107672,0.1756981,8.0040245,15.828446,23.656773,31.4851,39.313427,33.82774,28.342056,22.85637,17.370686,11.888905,9.511124,7.1333427,4.755562,2.377781,0.0,2.4402514,4.8805027,7.320754,9.761005,12.201257,15.668366,19.13938,22.610394,26.081408,29.548515,25.40204,21.251661,17.101282,12.950902,8.800523,8.480362,8.160201,7.8400397,7.519879,7.1997175,13.314012,19.4244,25.538694,31.649084,37.76338,31.371872,24.976461,18.584955,12.193448,5.7980375,5.5013027,5.2045684,4.9078336,4.6110992,4.3143644,7.9923115,11.674163,15.35211,19.03396,22.711908,21.122816,19.533724,17.94073,16.351637,14.762545,13.759113,12.755682,11.756155,10.752724,9.749292,13.845011,17.94073,22.036446,26.12826,30.223978,28.783253,27.346434,25.905708,24.464985,23.02426,18.95197,14.875772,10.799577,6.7233806,2.6510892,3.5569105,4.466636,5.3724575,6.278279,7.1880045,8.800523,10.413041,12.025558,13.638077,15.250595,17.72989,20.209187,22.688482,25.17168,27.650976,23.500597,19.350218,15.199838,11.0494585,6.899079,12.412095,17.92511,23.438128,28.951143,34.464157,29.283016,24.10578,18.928543,13.751305,8.574067,9.639969,10.705871,11.771772,12.83377,13.899672,11.197825,8.495979,5.794133,3.0883822,0.38653582,0.31235218,0.23816854,0.1639849,0.08589685,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.031235218,0.046852827,0.06637484,0.08199245,0.10151446,0.46462387,0.8316377,1.1947471,1.5617609,1.9248703,1.6047094,1.2845483,0.96438736,0.6442264,0.3240654,0.8316377,1.33921,1.8467822,2.3543546,2.8619268,3.8887846,4.911738,5.938596,6.9615493,7.988407,7.3832245,6.7780423,6.17286,5.5676775,4.9624953,4.1894236,3.416352,2.6432803,1.8741131,1.1010414,1.6749885,2.2489357,2.8267872,3.4007344,3.9746814,3.408543,2.8463092,2.280171,1.7140326,1.1517987,0.92924774,0.7106012,0.48805028,0.26940376,0.05075723,0.9917182,1.9287747,2.8697357,3.8106966,4.7516575,3.998108,3.2484627,2.4988174,1.7491722,0.999527,1.3040704,1.6047094,1.9092526,2.2098918,2.514435,2.3348327,2.1591344,1.979532,1.8038338,1.6242313,1.3274968,1.0307622,0.7340276,0.43338865,0.13665408,2.280171,4.423688,6.5633,8.706817,10.850334,8.679486,6.5086384,4.3416953,2.1708477,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.12103647,0.23816854,0.359205,0.48024148,0.60127795,0.5349031,0.46852827,0.40605783,0.339683,0.27330816,0.46071947,0.6442264,0.8316377,1.0151446,1.1986516,1.3782539,1.5539521,1.7335546,1.9092526,2.0888553,2.260649,2.4324427,2.6042364,2.77603,2.951728,2.6081407,2.2684577,1.9287747,1.5890918,1.2494087,1.1010414,0.95657855,0.80821127,0.659844,0.5114767,0.78088045,1.0463798,1.3157835,1.5812829,1.8506867,1.4992905,1.1439898,0.79259366,0.44119745,0.08589685,0.14446288,0.20302892,0.26159495,0.31625658,0.37482262,0.31625658,0.25378615,0.19522011,0.13665408,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.13274968,0.1639849,0.19912452,0.23035973,0.26159495,0.26940376,0.27721256,0.28502136,0.29283017,0.30063897,0.3553006,0.40996224,0.46462387,0.5192855,0.57394713,0.57785153,0.58175594,0.58175594,0.58566034,0.58566034,0.62079996,0.6559396,0.6910792,0.7262188,0.76135844,0.6442264,0.5270943,0.40996224,0.29283017,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.1835069,0.1717937,0.15617609,0.14055848,0.12494087,0.22255093,0.32016098,0.41777104,0.5153811,0.61299115,0.6676528,0.7223144,0.77697605,0.8316377,0.8862993,0.79649806,0.7066968,0.61689556,0.5270943,0.43729305,0.7262188,1.0112402,1.3001659,1.5890918,1.8741131,2.0068626,2.1396124,2.2723622,2.4051118,2.5378613,2.3816853,2.2216048,2.0654287,1.9092526,1.7491722,1.5539521,1.358732,1.1635119,0.96829176,0.77307165,0.8277333,0.8784905,0.93315214,0.98390937,1.038571,1.0073358,0.97610056,0.94876975,0.91753453,0.8862993,0.9097257,0.93315214,0.95657855,0.97610056,0.999527,1.038571,1.0815194,1.1205635,1.1596074,1.1986516,1.1283722,1.0580931,0.9917182,0.92143893,0.8511597,0.77697605,0.7066968,0.63251317,0.5583295,0.48805028,0.45681506,0.42557985,0.39824903,0.3670138,0.3357786,0.3240654,0.31235218,0.30063897,0.28892577,0.27330816,0.27721256,0.28111696,0.28111696,0.28502136,0.28892577,0.39824903,0.5075723,0.61689556,0.7262188,0.8394465,1.1908426,1.542239,1.893635,2.2489357,2.6003318,3.7208953,4.845363,5.9659266,7.0903945,8.210958,8.968412,9.725866,10.48332,11.240774,11.998228,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15617609,0.31625658,0.47243267,0.62860876,0.78868926,1.678893,2.5730011,3.4632049,4.357313,5.251421,6.5086384,7.7697606,9.030883,10.2881,11.549222,13.235924,14.918721,16.605423,18.28822,19.974922,19.443924,18.90902,18.378021,17.843119,17.31212,16.863113,16.41801,15.969006,15.523903,15.074897,14.133936,13.196879,12.2559185,11.314958,10.373997,11.560935,12.751778,13.938716,15.125654,16.312593,15.586374,14.856251,14.130032,13.403813,12.67369,12.263727,11.8537655,11.443803,11.033841,10.6238785,11.838148,13.048512,14.262781,15.473146,16.687416,17.93292,19.178425,20.423927,21.669432,22.911032,19.561056,16.211079,12.861101,9.511124,6.1611466,9.788337,13.415526,17.04662,20.67381,24.300999,25.456703,26.61631,27.772013,28.931622,30.087324,30.872108,31.656893,32.441677,33.226463,34.01125,33.370926,32.73451,32.094185,31.453865,30.813543,30.020948,29.228355,28.435762,27.643167,26.850574,25.8081,24.765623,23.723148,22.680674,21.638197,22.40346,23.168722,23.933987,24.69925,25.460608,24.82419,24.187773,23.551353,22.911032,22.274614,19.943687,17.616663,15.285735,12.954806,10.6238785,10.256865,9.889851,9.522837,9.155824,8.78881,10.545791,12.302772,14.059752,15.816733,17.573715,21.048632,24.52355,27.998468,31.473387,34.948303,35.924404,36.900505,37.876606,38.8488,39.8249,34.33141,28.84182,23.348326,17.854832,12.361338,12.619028,12.8767185,13.134409,13.392099,13.64979,13.536563,13.423335,13.314012,13.200784,13.087557,11.904523,10.721489,9.538455,8.359325,7.1762915,10.276386,13.376482,16.476578,19.576674,22.67677,18.139853,13.606842,9.069926,4.533011,0.0,0.71841,1.4407244,2.1591344,2.8814487,3.5998588,3.2211318,2.8463092,2.4675822,2.0888553,1.7140326,1.3743496,1.038571,0.698888,0.3631094,0.023426414,0.3631094,0.7066968,1.0463798,1.3860629,1.7257458,2.8111696,3.8965936,4.9781127,6.0635366,7.1489606,7.016211,6.883461,6.7507114,6.621866,6.4891167,5.813655,5.138193,4.462732,3.78727,3.1118085,6.211904,9.308095,12.404286,15.504381,18.600573,14.9109125,11.225157,7.535496,3.8497405,0.1639849,6.055728,11.947471,17.839214,23.730957,29.626604,26.405472,23.184341,19.96321,16.745981,13.524849,10.819098,8.113348,5.4115014,2.7057507,0.0,2.241127,4.4861584,6.727285,8.968412,11.213444,13.403813,15.594183,17.780647,19.971018,22.161386,19.049578,15.93777,12.825961,9.714153,6.5984397,6.3602715,6.1181984,5.8800297,5.6418614,5.3997884,10.237343,15.074897,19.91245,24.750006,29.58756,25.24196,20.892456,16.542952,12.197352,7.8517528,7.055255,6.2587566,5.466163,4.6696653,3.873167,6.559396,9.245625,11.931853,14.614178,17.300406,16.745981,16.191557,15.633226,15.078801,14.524376,13.583415,12.63855,11.697589,10.756628,9.811763,14.227642,18.64352,23.0594,27.471375,31.887253,29.333775,26.77639,24.222912,21.665527,19.11205,16.136894,13.16174,10.186585,7.211431,4.2362766,5.1030536,5.9659266,6.832704,7.6955767,8.562354,10.87376,13.189071,15.500477,17.811884,20.12329,23.348326,26.569458,29.794493,33.015625,36.23676,30.462147,24.687536,18.912924,13.138313,7.363703,11.4633255,15.562947,19.662569,23.762192,27.861814,24.730484,21.603058,18.471727,15.344301,12.212971,12.716639,13.224211,13.727879,14.231546,14.739119,11.908427,9.077735,6.2470436,3.416352,0.58566034,0.47633708,0.3631094,0.24988174,0.13665408,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.03513962,0.046852827,0.05466163,0.06637484,0.07418364,0.3553006,0.63641757,0.9136301,1.1947471,1.475864,1.2494087,1.0190489,0.79259366,0.5661383,0.3357786,0.7145056,1.0932326,1.4719596,1.8467822,2.2255092,3.7482262,5.2748475,6.801469,8.324185,9.850807,8.628729,7.406651,6.180669,4.958591,3.736513,3.3031244,2.87364,2.4402514,2.0068626,1.5734742,2.1122816,2.6510892,3.1859922,3.7247996,4.263607,3.8575494,3.4514916,3.049338,2.6432803,2.2372224,1.796025,1.358732,0.91753453,0.47633708,0.039044023,0.94096094,1.8467822,2.7526035,3.6584249,4.564246,3.9746814,3.3890212,2.7994564,2.2137961,1.6242313,1.8311646,2.0341935,2.241127,2.4441557,2.6510892,2.5808098,2.514435,2.4480603,2.3816853,2.3114061,1.9053483,1.4992905,1.0893283,0.6832704,0.27330816,1.8467822,3.4202564,4.9937305,6.5633,8.136774,6.5086384,4.884407,3.2562714,1.6281357,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.08980125,0.1796025,0.26940376,0.359205,0.44900626,0.45681506,0.46462387,0.47243267,0.48024148,0.48805028,0.7340276,0.97610056,1.2220778,1.4680552,1.7140326,2.2059872,2.697942,3.1898966,3.6818514,4.173806,3.7833657,3.3890212,2.998581,2.6042364,2.2137961,1.9561055,1.7023194,1.4485333,1.1908426,0.93705654,0.8433509,0.74574083,0.6520352,0.5583295,0.46071947,0.76135844,1.0580931,1.3548276,1.6515622,1.9482968,1.5812829,1.2142692,0.8472553,0.48024148,0.113227665,0.1756981,0.24207294,0.30844778,0.3709182,0.43729305,0.3670138,0.29673457,0.22645533,0.15617609,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.113227665,0.15617609,0.19522011,0.23426414,0.27330816,0.28892577,0.30454338,0.32016098,0.3357786,0.3513962,0.42167544,0.4958591,0.5661383,0.64032197,0.7106012,0.679366,0.6481308,0.61689556,0.58175594,0.5505207,0.60908675,0.6637484,0.7223144,0.78088045,0.8394465,0.7145056,0.59346914,0.46852827,0.3474918,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.14446288,0.14055848,0.13665408,0.12884527,0.12494087,0.19522011,0.26549935,0.3357786,0.40605783,0.47633708,0.5231899,0.5700427,0.61689556,0.6637484,0.7106012,0.6442264,0.57785153,0.5114767,0.44119745,0.37482262,0.6754616,0.97610056,1.2767396,1.5734742,1.8741131,1.9287747,1.979532,2.0341935,2.084951,2.135708,2.0107672,1.8819219,1.7530766,1.6281357,1.4992905,1.3470187,1.1947471,1.0424755,0.8902037,0.737932,0.8433509,0.94876975,1.0541886,1.1557031,1.261122,1.1635119,1.0659018,0.96829176,0.8706817,0.77307165,0.79649806,0.8160201,0.8355421,0.8550641,0.8745861,0.94096094,1.0112402,1.077615,1.1439898,1.2142692,1.1361811,1.0580931,0.98000497,0.9019169,0.8238289,0.78088045,0.7340276,0.6910792,0.6442264,0.60127795,0.58956474,0.58175594,0.5700427,0.5583295,0.5505207,0.5231899,0.4997635,0.47633708,0.44900626,0.42557985,0.40605783,0.38653582,0.3631094,0.3435874,0.3240654,0.40605783,0.49195468,0.57394713,0.6559396,0.737932,1.0034313,1.2728351,1.5383345,1.8077383,2.0732377,2.9439192,3.814601,4.6852827,5.5559645,6.426646,7.027924,7.629202,8.234385,8.835662,9.43694,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11713207,0.23426414,0.3513962,0.46852827,0.58566034,1.5461433,2.5027218,3.4593005,4.415879,5.376362,6.703859,8.031356,9.358852,10.686349,12.013845,14.016804,16.015858,18.018816,20.021774,22.024733,21.583536,21.138433,20.697237,20.256039,19.810938,19.260416,18.705992,18.15547,17.601046,17.050524,16.226696,15.406772,14.582942,13.759113,12.939189,13.626364,14.313539,15.000713,15.687888,16.375063,15.426293,14.481428,13.532659,12.583888,11.639023,11.260296,10.881569,10.506746,10.128019,9.749292,11.736633,13.723974,15.711315,17.698656,19.685997,21.040823,22.39565,23.754383,25.109211,26.464039,22.899319,19.338505,15.773785,12.212971,8.648251,13.770826,18.893402,24.015978,29.138554,34.26113,35.205994,36.146957,37.09182,38.032784,38.973743,39.852234,40.730724,41.609215,42.483803,43.362293,42.878147,42.394,41.90595,41.421803,40.937656,39.40713,37.872704,36.338272,34.807747,33.273315,30.778402,28.28349,25.788576,23.293663,20.79875,20.986162,21.169668,21.353176,21.540586,21.724094,21.688955,21.64991,21.610867,21.575727,21.536682,19.931974,18.32336,16.714746,15.1061325,13.501423,12.529227,11.560935,10.588739,9.620447,8.648251,9.456462,10.260769,11.065076,11.869383,12.67369,14.825015,16.976341,19.123762,21.275087,23.426414,25.163872,26.90133,28.63879,30.37625,32.11371,27.541653,22.973503,18.401447,13.833297,9.261242,10.8425255,12.423808,14.001186,15.582469,17.163752,17.562002,17.964155,18.362404,18.764557,19.162806,16.320402,13.477997,10.6355915,7.793187,4.950782,8.738052,12.525322,16.312593,20.099863,23.887133,19.11205,14.33306,9.554072,4.7789884,0.0,0.5544251,1.1088502,1.6632754,2.2216048,2.77603,2.5651922,2.3543546,2.1435168,1.9365835,1.7257458,1.3860629,1.0502841,0.7106012,0.37482262,0.039044023,0.4958591,0.95657855,1.4172981,1.8780174,2.338737,2.979059,3.619381,4.2557983,4.8961205,5.5364423,6.1064854,6.676528,7.2465706,7.816613,8.386656,7.4144597,6.4383593,5.462259,4.4861584,3.513962,8.378847,13.243732,18.108618,22.973503,27.838388,22.301945,16.761599,11.225157,5.688714,0.14836729,4.1074314,8.066495,12.021654,15.980719,19.935879,18.983204,18.026625,17.073952,16.117373,15.160794,12.130978,9.097258,6.0635366,3.0337205,0.0,2.0459068,4.0918136,6.133816,8.179723,10.22563,11.135355,12.045081,12.954806,13.864532,14.774258,12.70102,10.6238785,8.550641,6.473499,4.4002614,4.240181,4.0801005,3.9200199,3.7599394,3.5998588,7.1606736,10.725393,14.286208,17.850927,21.411741,19.108145,16.808453,14.504854,12.201257,9.901564,8.609207,7.3168497,6.0205884,4.728231,3.435874,5.12648,6.817086,8.507692,10.198298,11.888905,12.369146,12.845484,13.325725,13.805966,14.286208,13.403813,12.521418,11.639023,10.756628,9.874233,14.610273,19.346313,24.07845,28.81449,33.55053,29.88039,26.210253,22.540113,18.869976,15.199838,13.325725,11.4516115,9.573594,7.699481,5.825368,6.649197,7.4691215,8.292951,9.116779,9.936704,12.950902,15.961197,18.975395,21.989594,24.999887,28.96676,32.92973,36.896603,40.85957,44.826443,37.423695,30.024853,22.62601,15.223265,7.824422,10.514555,13.200784,15.8870125,18.573242,21.263374,20.177952,19.096432,18.014912,16.933393,15.851873,15.793307,15.738646,15.683984,15.629322,15.57466,12.619028,9.659492,6.703859,3.7443218,0.78868926,0.63641757,0.48805028,0.3357786,0.18741131,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.042948425,0.046852827,0.046852827,0.05075723,0.24597734,0.44119745,0.63641757,0.8316377,1.0268579,0.8902037,0.75354964,0.62079996,0.48414588,0.3513962,0.59737355,0.8433509,1.0932326,1.33921,1.5890918,3.611572,5.6379566,7.6643414,9.686822,11.713207,9.874233,8.031356,6.192382,4.3534083,2.5105307,2.4207294,2.3270237,2.233318,2.1435168,2.0498111,2.5495746,3.049338,3.5491016,4.0488653,4.548629,4.3065557,4.0605783,3.814601,3.5686235,3.3265507,2.6667068,2.0068626,1.3431144,0.6832704,0.023426414,0.8941081,1.7647898,2.6354716,3.506153,4.376835,3.951255,3.5256753,3.1000953,2.6745155,2.2489357,2.358259,2.463678,2.5730011,2.67842,2.787743,2.8306916,2.87364,2.9165885,2.9556324,2.998581,2.4831998,1.9639144,1.4485333,0.92924774,0.41386664,1.4133936,2.416825,3.4202564,4.423688,5.423215,4.3416953,3.2562714,2.1708477,1.0854238,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.37872702,0.46071947,0.5388075,0.62079996,0.698888,1.0034313,1.3118792,1.6164225,1.9209659,2.2255092,3.0337205,3.8419318,4.646239,5.45445,6.262661,5.3060827,4.349504,3.3890212,2.4324427,1.475864,1.3040704,1.1361811,0.96438736,0.79649806,0.62470436,0.58175594,0.5388075,0.4958591,0.45681506,0.41386664,0.7418364,1.0659018,1.3938715,1.7218413,2.0498111,1.6671798,1.2845483,0.9019169,0.5192855,0.13665408,0.21083772,0.28111696,0.3553006,0.42557985,0.4997635,0.42167544,0.339683,0.26159495,0.1796025,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.09761006,0.14446288,0.19131571,0.23816854,0.28892577,0.30844778,0.3318742,0.3553006,0.37872702,0.39824903,0.49195468,0.58175594,0.6715572,0.76135844,0.8511597,0.78088045,0.7145056,0.6481308,0.58175594,0.5114767,0.59346914,0.6715572,0.75354964,0.8316377,0.9136301,0.78478485,0.6559396,0.5309987,0.40215343,0.27330816,0.21864653,0.1639849,0.10932326,0.05466163,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.10541886,0.10932326,0.113227665,0.12103647,0.12494087,0.1678893,0.21083772,0.25378615,0.29673457,0.3357786,0.37872702,0.41777104,0.45681506,0.4958591,0.5388075,0.49195468,0.44900626,0.40215343,0.359205,0.31235218,0.62470436,0.93705654,1.2494087,1.5617609,1.8741131,1.8467822,1.8194515,1.7921207,1.7647898,1.737459,1.639849,1.542239,1.4446288,1.3470187,1.2494087,1.1400855,1.0307622,0.92143893,0.80821127,0.698888,0.8589685,1.0151446,1.1713207,1.3314011,1.4875772,1.3235924,1.1557031,0.9917182,0.8277333,0.6637484,0.679366,0.698888,0.7145056,0.7340276,0.74964523,0.8433509,0.94096094,1.0346665,1.1283722,1.2259823,1.1400855,1.0541886,0.96829176,0.8862993,0.80040246,0.78088045,0.76526284,0.74574083,0.7301232,0.7106012,0.7223144,0.7340276,0.7418364,0.75354964,0.76135844,0.7262188,0.6871748,0.6481308,0.61299115,0.57394713,0.5309987,0.48805028,0.44900626,0.40605783,0.3631094,0.41777104,0.47243267,0.5270943,0.58175594,0.63641757,0.8199245,1.0034313,1.1869383,1.3665408,1.5500476,2.1669433,2.7838387,3.4007344,4.0215344,4.6384296,5.083532,5.532538,5.9815445,6.426646,6.8756523,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.078088045,0.15617609,0.23426414,0.30844778,0.38653582,1.4094892,2.4324427,3.455396,4.478349,5.5013027,6.8951745,8.289046,9.686822,11.080693,12.4745655,14.79378,17.1169,19.436115,21.75533,24.074545,23.723148,23.371752,23.01645,22.665054,22.31366,21.653814,20.997875,20.341936,19.682093,19.026152,18.319456,17.616663,16.909966,16.20327,15.500477,15.687888,15.875299,16.062712,16.250122,16.437534,15.270117,14.102701,12.935285,11.767868,10.600452,10.256865,9.909373,9.565785,9.218294,8.874706,11.639023,14.399435,17.163752,19.924164,22.688482,24.152632,25.616783,27.080935,28.548988,30.01314,26.237583,22.462027,18.68647,14.9109125,11.139259,17.753317,24.371279,30.98924,37.6072,44.225163,44.95138,45.681507,46.407726,47.133945,47.864067,48.83236,49.804554,50.772846,51.74114,52.713333,52.381462,52.05349,51.721615,51.393646,51.06177,48.78941,46.517048,44.244686,41.972324,39.699963,35.752613,31.805262,27.85791,23.910559,19.96321,19.568865,19.170614,18.77627,18.381926,17.987581,18.549814,19.11205,19.674282,20.236517,20.79875,19.916355,19.030056,18.143757,17.261362,16.375063,14.801589,13.232019,11.6585455,10.085071,8.511597,8.36323,8.218767,8.070399,7.9220324,7.773665,8.601398,9.425227,10.249056,11.076789,11.900618,14.399435,16.898252,19.400974,21.899792,24.39861,20.751898,17.105186,13.458474,9.811763,6.1611466,9.066022,11.966993,14.871868,17.772839,20.67381,21.58744,22.50107,23.410795,24.324427,25.238056,20.73628,16.234505,11.728825,7.2270484,2.7252727,7.1997175,11.674163,16.148607,20.626957,25.101402,20.080341,15.059279,10.0382185,5.0210614,0.0,0.39044023,0.78088045,1.1713207,1.5617609,1.9482968,1.9092526,1.8663043,1.8233559,1.7804074,1.737459,1.4016805,1.0619974,0.7262188,0.38653582,0.05075723,0.62860876,1.2103647,1.7882162,2.3699722,2.951728,3.1469483,3.338264,3.533484,3.7287042,3.9239242,5.196759,6.4695945,7.7424297,9.0152645,10.2881,9.01136,7.7385254,6.461786,5.1889505,3.912211,10.545791,17.175465,23.809046,30.442625,37.076202,29.689075,22.301945,14.9109125,7.523783,0.13665408,2.1591344,4.181615,6.2040954,8.226576,10.249056,11.560935,12.86891,14.180789,15.488764,16.800642,13.438952,10.081166,6.719476,3.3616903,0.0,1.8467822,3.6935644,5.5442514,7.3910336,9.237816,8.866898,8.495979,8.128965,7.758047,7.387129,6.348558,5.3138914,4.2753205,3.2367494,2.1981785,2.1200905,2.0380979,1.9600099,1.8819219,1.7999294,4.087909,6.375889,8.663869,10.951848,13.235924,12.978233,12.720543,12.466757,12.209065,11.951375,10.159255,8.371038,6.578918,4.7907014,2.998581,3.6935644,4.388548,5.083532,5.7785153,6.473499,7.988407,9.503315,11.018223,12.533132,14.051944,13.228115,12.404286,11.584361,10.760532,9.936704,14.992905,20.049105,25.101402,30.157602,35.213802,30.427008,25.644114,20.857317,16.07052,11.287627,10.510651,9.737579,8.960603,8.187531,7.4144597,8.191436,8.972317,9.753197,10.534078,11.311053,15.024139,18.737226,22.450314,26.163399,29.876486,34.58129,39.29,43.99871,48.703514,53.412224,44.385246,35.36217,26.339098,17.31212,8.289046,9.561881,10.838621,12.111456,13.388195,14.661031,15.629322,16.59371,17.558098,18.522484,19.486872,18.87388,18.256985,17.643993,17.027098,16.414106,13.325725,10.241247,7.1567693,4.0722914,0.9878138,0.80040246,0.61299115,0.42557985,0.23816854,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.046852827,0.039044023,0.03513962,0.031235218,0.023426414,0.13665408,0.24597734,0.3553006,0.46462387,0.57394713,0.5309987,0.48805028,0.44900626,0.40605783,0.3631094,0.48024148,0.59737355,0.7145056,0.8316377,0.94876975,3.474918,6.001066,8.52331,11.0494585,13.575606,11.115833,8.659965,6.2040954,3.7443218,1.2884527,1.53443,1.7843118,2.0302892,2.2762666,2.5261483,2.9868677,3.4514916,3.912211,4.376835,4.8375545,4.7516575,4.6657605,4.5837684,4.4978714,4.4119744,3.533484,2.6510892,1.7725986,0.8941081,0.011713207,0.8472553,1.6827974,2.5183394,3.3538816,4.1894236,3.9239242,3.6623292,3.4007344,3.1391394,2.87364,2.8853533,2.893162,2.9048753,2.9165885,2.9243972,3.076669,3.2289407,3.3812122,3.533484,3.6857557,3.0610514,2.4324427,1.8038338,1.1791295,0.5505207,0.98390937,1.4133936,1.8467822,2.280171,2.7135596,2.1708477,1.6281357,1.0854238,0.5427119,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.30063897,0.45681506,0.60908675,0.76135844,0.9136301,1.2767396,1.6437533,2.0068626,2.3738766,2.736986,3.8614538,4.9820175,6.1064854,7.2270484,8.351517,6.8287997,5.3060827,3.7833657,2.260649,0.737932,0.6520352,0.5661383,0.48414588,0.39824903,0.31235218,0.3240654,0.3318742,0.3435874,0.3513962,0.3631094,0.71841,1.077615,1.43682,1.7921207,2.1513257,1.7530766,1.3548276,0.95657855,0.5583295,0.1639849,0.24207294,0.3240654,0.40215343,0.48414588,0.5622339,0.47243267,0.38263142,0.29283017,0.20302892,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.078088045,0.13665408,0.19131571,0.24597734,0.30063897,0.3318742,0.359205,0.39044023,0.42167544,0.44900626,0.5583295,0.6637484,0.77307165,0.8784905,0.9878138,0.8862993,0.78088045,0.679366,0.57785153,0.47633708,0.57785153,0.679366,0.78088045,0.8862993,0.9878138,0.8550641,0.7223144,0.58956474,0.45681506,0.3240654,0.26159495,0.19522011,0.12884527,0.06637484,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.06637484,0.078088045,0.093705654,0.10932326,0.12494087,0.14055848,0.15617609,0.1717937,0.1835069,0.19912452,0.23426414,0.26549935,0.29673457,0.3318742,0.3631094,0.339683,0.31625658,0.29673457,0.27330816,0.24988174,0.57394713,0.9019169,1.2259823,1.5500476,1.8741131,1.7686942,1.6593709,1.5539521,1.4446288,1.33921,1.2689307,1.2025559,1.1361811,1.0659018,0.999527,0.93315214,0.8667773,0.79649806,0.7301232,0.6637484,0.8706817,1.0815194,1.2923572,1.5031948,1.7140326,1.4797685,1.2494087,1.0151446,0.78088045,0.5505207,0.5661383,0.58175594,0.59346914,0.60908675,0.62470436,0.74574083,0.8706817,0.9917182,1.116659,1.2376955,1.1439898,1.0541886,0.96048295,0.8667773,0.77307165,0.78478485,0.79649806,0.80430686,0.8160201,0.8238289,0.8550641,0.8862993,0.9136301,0.94486535,0.97610056,0.92534333,0.8745861,0.8238289,0.77307165,0.7262188,0.659844,0.59346914,0.5309987,0.46462387,0.39824903,0.42557985,0.45681506,0.48414588,0.5114767,0.5388075,0.63641757,0.7340276,0.8316377,0.92924774,1.0268579,1.3899672,1.756981,2.1200905,2.4831998,2.8502135,3.1430438,3.435874,3.7287042,4.0215344,4.3143644,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,1.2767396,2.3621633,3.4514916,4.5369153,5.6262436,7.08649,8.550641,10.010887,11.475039,12.939189,15.57466,18.214037,20.849508,23.488884,26.124355,25.86276,25.601166,25.335667,25.074072,24.812477,24.051117,23.285854,22.524496,21.763138,21.00178,20.412214,19.826555,19.23699,18.651329,18.061766,17.749413,17.437061,17.124708,16.812357,16.500004,15.113941,13.723974,12.337912,10.951848,9.561881,9.249529,8.937177,8.624825,8.312472,8.00012,11.537509,15.074897,18.612286,22.149673,25.687063,27.260536,28.837915,30.411388,31.988768,33.56224,29.575848,25.589453,21.599154,17.612759,13.626364,21.735807,29.849155,37.9625,46.07585,54.189198,54.700676,55.21215,55.72363,56.23901,56.75049,57.812485,58.87448,59.936478,60.998478,62.064377,61.88868,61.712982,61.537285,61.361588,61.185886,58.175594,55.161396,52.1511,49.1369,46.12661,40.726818,35.32703,29.92334,24.52355,19.123762,18.151566,17.175465,16.199366,15.223265,14.251068,15.410676,16.574188,17.7377,18.90121,20.06082,19.900738,19.736753,19.576674,19.412687,19.248703,17.073952,14.899199,12.724447,10.549695,8.374943,7.2739015,6.1767645,5.0757227,3.9746814,2.87364,2.3738766,1.8741131,1.3743496,0.8745861,0.37482262,3.638903,6.899079,10.163159,13.423335,16.687416,13.962143,11.23687,8.511597,5.786324,3.0610514,7.2856145,11.514082,15.738646,19.96321,24.187773,25.612879,27.037985,28.463093,29.888199,31.313307,25.148254,18.987108,12.825961,6.66091,0.4997635,5.661383,10.823003,15.988527,21.150146,26.311768,21.048632,15.789403,10.526268,5.263134,0.0,0.22645533,0.44900626,0.6754616,0.9019169,1.1244678,1.2494087,1.3743496,1.4992905,1.6242313,1.7491722,1.4133936,1.0737107,0.737932,0.39824903,0.062470436,0.76135844,1.4641509,2.1630387,2.8619268,3.5608149,3.310933,3.0610514,2.8111696,2.5612879,2.3114061,4.2870336,6.262661,8.238289,10.213917,12.185639,10.612165,9.0386915,7.461313,5.8878384,4.3143644,12.712734,21.111103,29.513376,37.911747,46.31402,37.076202,27.838388,18.600573,9.362757,0.12494087,0.21083772,0.30063897,0.38653582,0.47633708,0.5622339,4.138666,7.7111945,11.287627,14.864059,18.436588,14.750832,11.061172,7.375416,3.6857557,0.0,1.6515622,3.2992198,4.950782,6.5984397,8.250002,6.5984397,4.950782,3.2992198,1.6515622,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0112402,2.0263848,3.0376248,4.0488653,5.0640097,6.8483214,8.636538,10.424754,12.212971,14.001186,11.713207,9.425227,7.137247,4.8492675,2.5612879,2.260649,1.9639144,1.6632754,1.3626363,1.0619974,3.611572,6.1611466,8.710721,11.2642,13.813775,13.048512,12.287154,11.525795,10.764437,9.999174,15.375536,20.747993,26.124355,31.500717,36.873177,30.973623,25.074072,19.174519,13.274967,7.375416,7.699481,8.023546,8.351517,8.675582,8.999647,9.737579,10.475512,11.213444,11.951375,12.689307,17.101282,21.513256,25.925232,30.337206,34.74918,40.199726,45.650272,51.100815,56.55136,62.001907,51.3507,40.69949,30.048279,19.400974,8.749765,8.6131115,8.476458,8.335898,8.1992445,8.062591,11.076789,14.087084,17.101282,20.111576,23.125774,21.95055,20.775324,19.6001,18.424873,17.24965,14.036326,10.826907,7.6135845,4.4002614,1.1869383,0.96438736,0.737932,0.5114767,0.28892577,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.1756981,0.22645533,0.27330816,0.3240654,0.37482262,0.3631094,0.3513962,0.3357786,0.3240654,0.31235218,3.338264,6.364176,9.386183,12.412095,15.438006,12.361338,9.288573,6.211904,3.1391394,0.062470436,0.6481308,1.2376955,1.8233559,2.4129205,2.998581,3.4241607,3.8497405,4.2753205,4.7009,5.12648,5.2006636,5.2748475,5.349031,5.423215,5.5013027,4.4002614,3.2992198,2.1981785,1.1010414,0.0,0.80040246,1.6008049,2.4012074,3.2016098,3.998108,3.900498,3.7989833,3.7013733,3.5998588,3.4983444,3.4124475,3.3265507,3.2367494,3.1508527,3.0610514,3.3265507,3.5881457,3.8497405,4.1113358,4.376835,3.638903,2.900971,2.1630387,1.4251068,0.6871748,0.5505207,0.41386664,0.27330816,0.13665408,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22645533,0.44900626,0.6754616,0.9019169,1.1244678,1.5500476,1.9756275,2.4012074,2.8267872,3.2484627,4.689187,6.126007,7.562827,8.999647,10.436467,8.351517,6.262661,4.173806,2.0888553,0.0,0.0,0.0,0.0,0.0,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.698888,1.0893283,1.475864,1.8623998,2.2489357,1.8389735,1.4251068,1.0112402,0.60127795,0.18741131,0.27330816,0.3631094,0.44900626,0.5388075,0.62470436,0.5231899,0.42557985,0.3240654,0.22645533,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.3513962,0.38653582,0.42557985,0.46071947,0.4997635,0.62470436,0.74964523,0.8745861,0.999527,1.1244678,0.9878138,0.8511597,0.7106012,0.57394713,0.43729305,0.5622339,0.6871748,0.81211567,0.93705654,1.0619974,0.92534333,0.78868926,0.6481308,0.5114767,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.5231899,0.8628729,1.1986516,1.5383345,1.8741131,1.6867018,1.4992905,1.3118792,1.1244678,0.93705654,0.9019169,0.8628729,0.8238289,0.78868926,0.74964523,0.7262188,0.698888,0.6754616,0.6481308,0.62470436,0.8862993,1.1517987,1.4133936,1.6749885,1.9365835,1.6359446,1.33921,1.038571,0.737932,0.43729305,0.44900626,0.46071947,0.47633708,0.48805028,0.4997635,0.6481308,0.80040246,0.94876975,1.1010414,1.2494087,1.1517987,1.0502841,0.94876975,0.8511597,0.74964523,0.78868926,0.8238289,0.8628729,0.9019169,0.93705654,0.9878138,1.038571,1.0893283,1.1361811,1.1869383,1.1244678,1.0619974,0.999527,0.93705654,0.8745861,0.78868926,0.698888,0.61299115,0.5231899,0.43729305,0.43729305,0.43729305,0.43729305,0.43729305,0.43729305,0.44900626,0.46071947,0.47633708,0.48805028,0.4997635,0.61299115,0.7262188,0.8394465,0.94876975,1.0619974,1.1986516,1.33921,1.475864,1.6125181,1.7491722,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,1.1400855,2.0810463,3.018103,3.959064,4.900025,6.481308,8.058686,9.639969,11.221252,12.798631,14.840633,16.88654,18.928543,20.970545,23.012547,22.911032,22.813423,22.711908,22.614298,22.512783,22.391747,22.266806,22.14577,22.020828,21.899792,21.39222,20.884647,20.377075,19.869503,19.36193,18.694279,18.026625,17.358973,16.69132,16.023666,14.700074,13.376482,12.0489855,10.725393,9.4018,9.8312845,10.260769,10.690253,11.119738,11.549222,15.063184,18.58105,22.095013,25.608974,29.12684,30.954102,32.78136,34.60862,36.435883,38.26314,35.213802,32.16056,29.111223,26.061886,23.012547,29.341583,35.67062,42.00356,48.332596,54.661633,55.645542,56.625546,57.609455,58.593365,59.573368,60.27226,60.971146,61.66613,62.365017,63.063904,61.68565,60.311302,58.93695,57.562603,56.18825,54.15406,52.115963,50.081768,48.047573,46.013382,40.996223,35.98297,30.965815,25.952562,20.93931,19.924164,18.90902,17.893875,16.87873,15.863586,16.847496,17.831406,18.81922,19.803127,20.787037,19.721136,18.651329,17.585428,16.515621,15.449719,16.39068,17.335546,18.276506,19.221373,20.162333,17.027098,13.891863,10.756628,7.621393,4.4861584,3.7013733,2.9165885,2.1318035,1.3470187,0.5622339,3.2289407,5.891743,8.55845,11.221252,13.887959,11.607788,9.327617,7.0474463,4.7672753,2.4871042,5.8683167,9.253433,12.634645,16.015858,19.400974,20.529346,21.661623,22.789995,23.918367,25.050644,20.119385,15.192029,10.260769,5.3295093,0.39824903,4.533011,8.663869,12.798631,16.92949,21.06425,16.8514,12.63855,8.4257,4.21285,0.0,0.18741131,0.37482262,0.5622339,0.74964523,0.93705654,1.0659018,1.1908426,1.319688,1.4485333,1.5734742,1.358732,1.1439898,0.92924774,0.7145056,0.4997635,1.1361811,1.7765031,2.4129205,3.049338,3.6857557,3.5451972,3.4007344,3.260176,3.1157131,2.9751544,4.4314966,5.891743,7.348085,8.804427,10.260769,8.960603,7.656533,6.356367,5.0522966,3.7482262,10.436467,17.124708,23.81295,30.50119,37.18943,29.774971,22.364416,14.949956,7.535496,0.12494087,0.21083772,0.30063897,0.38653582,0.47633708,0.5622339,3.4593005,6.3524623,9.249529,12.142691,15.035853,12.357433,9.679013,6.996689,4.318269,1.6359446,2.7486992,3.8614538,4.9742084,6.086963,7.1997175,5.840986,4.4861584,3.1274261,1.7686942,0.41386664,0.3474918,0.28111696,0.21864653,0.15227169,0.08589685,0.46071947,0.8316377,1.2064602,1.5773785,1.9482968,2.3855898,2.8189783,3.2562714,3.68966,4.126953,6.250948,8.378847,10.506746,12.634645,14.762545,12.704925,10.647305,8.589685,6.532065,4.474445,4.154284,3.8341231,3.513962,3.193801,2.87364,5.3334136,7.793187,10.256865,12.716639,15.176412,14.614178,14.048039,13.4858055,12.923572,12.361338,17.761126,23.15701,28.556799,33.952682,39.348564,33.058575,26.768581,20.47859,14.188598,7.898606,8.55845,9.218294,9.878138,10.541886,11.20173,11.927949,12.654168,13.384291,14.11051,14.836729,17.698656,20.560583,23.426414,26.28834,29.150267,34.140095,39.12992,44.119747,49.109573,54.099396,45.509712,36.92003,28.330343,19.740658,11.150972,10.346666,9.546264,8.741957,7.941554,7.137247,11.240774,15.344301,19.443924,23.54745,27.650976,25.382519,23.114061,20.845604,18.58105,16.312593,13.239828,10.167064,7.094299,4.0215344,0.94876975,0.76916724,0.58956474,0.40996224,0.23035973,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.1835069,0.23426414,0.28111696,0.3279698,0.37482262,0.5466163,0.7145056,0.8862993,1.0541886,1.2259823,3.4593005,5.688714,7.9220324,10.155351,12.388668,9.956225,7.5276875,5.099149,2.6667068,0.23816854,0.8316377,1.4290112,2.0224805,2.6159496,3.213323,3.4710135,3.7287042,3.9863946,4.2440853,4.5017757,4.478349,4.4588275,4.4393053,4.4197836,4.4002614,3.521771,2.639376,1.7608855,0.8784905,0.0,0.64032197,1.2806439,1.9209659,2.5612879,3.2016098,3.1469483,3.096191,3.0415294,2.9907722,2.9361105,3.0024853,3.06886,3.1313305,3.1977055,3.2640803,3.5530062,3.8419318,4.1308575,4.423688,4.7126136,3.8809757,3.049338,2.2137961,1.3821584,0.5505207,0.44119745,0.3318742,0.21864653,0.10932326,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1796025,0.359205,0.5388075,0.71841,0.9019169,1.2415999,1.5812829,1.9209659,2.260649,2.6003318,3.7482262,4.900025,6.0518236,7.1997175,8.351517,6.703859,5.056201,3.408543,1.7608855,0.113227665,0.20693332,0.30063897,0.39824903,0.49195468,0.58566034,0.5192855,0.45291066,0.38653582,0.31625658,0.24988174,0.5583295,0.8706817,1.1791295,1.4914817,1.7999294,1.475864,1.1517987,0.8238289,0.4997635,0.1756981,0.24597734,0.31625658,0.38653582,0.45681506,0.5231899,0.44119745,0.359205,0.27721256,0.19522011,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05466163,0.10932326,0.1639849,0.21864653,0.27330816,0.30454338,0.3357786,0.3631094,0.39434463,0.42557985,0.5270943,0.62860876,0.7340276,0.8355421,0.93705654,0.8316377,0.7262188,0.62079996,0.5192855,0.41386664,0.5388075,0.6676528,0.79649806,0.92143893,1.0502841,0.93315214,0.8160201,0.698888,0.58175594,0.46071947,0.37872702,0.29283017,0.20693332,0.12103647,0.039044023,0.046852827,0.058566034,0.06637484,0.078088045,0.08589685,0.10932326,0.12884527,0.14836729,0.1678893,0.18741131,0.16008049,0.13274968,0.10541886,0.078088045,0.05075723,0.07418364,0.093705654,0.11713207,0.14055848,0.1639849,0.1796025,0.19912452,0.21474212,0.23426414,0.24988174,0.60127795,0.95657855,1.3079748,1.6593709,2.0107672,1.8077383,1.6008049,1.397776,1.1908426,0.9878138,0.92143893,0.8589685,0.79259366,0.7262188,0.6637484,0.6871748,0.7106012,0.737932,0.76135844,0.78868926,1.1400855,1.4914817,1.8467822,2.1981785,2.5495746,2.3621633,2.174752,1.9873407,1.7999294,1.6125181,1.4212024,1.2259823,1.0346665,0.8433509,0.6481308,0.75354964,0.8589685,0.96438736,1.0698062,1.175225,1.0893283,0.999527,0.9136301,0.8238289,0.737932,0.76916724,0.79649806,0.8277333,0.8589685,0.8862993,0.92143893,0.95657855,0.9917182,1.0268579,1.0619974,1.0190489,0.97610056,0.93315214,0.8941081,0.8511597,0.78868926,0.7301232,0.6715572,0.60908675,0.5505207,0.5661383,0.58566034,0.60127795,0.62079996,0.63641757,0.64032197,0.6442264,0.6442264,0.6481308,0.6481308,0.79649806,0.94486535,1.0932326,1.2415999,1.3860629,1.5110037,1.6359446,1.7608855,1.8858263,2.0107672,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.042948425,0.08589685,0.12884527,0.1717937,0.21083772,1.0034313,1.796025,2.5886188,3.3812122,4.173806,5.872221,7.570636,9.269051,10.963562,12.661977,14.11051,15.559043,17.003672,18.452206,19.900738,19.96321,20.025679,20.08815,20.15062,20.21309,20.728472,21.247757,21.763138,22.282423,22.801708,22.372225,21.946646,21.51716,21.091581,20.662096,19.639143,18.61619,17.593237,16.574188,15.551234,14.286208,13.025085,11.763964,10.498938,9.237816,10.409137,11.584361,12.755682,13.927003,15.098324,18.592764,22.0833,25.57774,29.068275,32.562714,34.64376,36.7209,38.80195,40.882996,42.964043,40.85176,38.73948,36.623295,34.511013,32.39873,36.947357,41.495987,46.044617,50.58934,55.13797,56.590405,58.042843,59.49528,60.94772,62.400158,62.732033,63.063904,63.39578,63.73156,64.06343,61.486526,58.913525,56.33662,53.76362,51.186714,50.12862,49.074432,48.01634,46.958244,45.900154,41.26953,36.638912,32.00829,27.381573,22.750952,21.696764,20.63867,19.584482,18.530293,17.476105,18.284315,19.088623,19.896833,20.705046,21.513256,19.541533,17.565907,15.594183,13.622459,11.650736,15.711315,19.767988,23.828568,27.889145,31.949724,26.780294,21.610867,16.441439,11.268105,6.098676,5.02887,3.959064,2.8892577,1.8194515,0.74964523,2.8189783,4.884407,6.9537406,9.019169,11.088503,9.253433,7.4183645,5.5832953,3.7482262,1.9131571,4.4510183,6.9927845,9.530646,12.072412,14.614178,15.445815,16.281357,17.1169,17.952442,18.787983,15.090515,11.393045,7.6955767,3.998108,0.30063897,3.4007344,6.504734,9.608734,12.708829,15.812829,12.650263,9.487698,6.3251314,3.1625657,0.0,0.14836729,0.30063897,0.44900626,0.60127795,0.74964523,0.8784905,1.0112402,1.1400855,1.2689307,1.4016805,1.3079748,1.2142692,1.1205635,1.0307622,0.93705654,1.5110037,2.0888553,2.6628022,3.2367494,3.8106966,3.775557,3.7443218,3.7091823,3.6740425,3.638903,4.575959,5.5169206,6.4578815,7.3988423,8.335898,7.309041,6.278279,5.2475166,4.2167544,3.1859922,8.164105,13.138313,18.112522,23.086731,28.06094,22.47374,16.88654,11.29934,5.7121406,0.12494087,0.21083772,0.30063897,0.38653582,0.47633708,0.5622339,2.77603,4.9937305,7.2075267,9.421323,11.639023,9.964035,8.292951,6.621866,4.9468775,3.2757936,3.8497405,4.423688,5.001539,5.575486,6.1494336,5.083532,4.0215344,2.9556324,1.8897307,0.8238289,0.6949836,0.5661383,0.43338865,0.30454338,0.1756981,0.92143893,1.6632754,2.4090161,3.154757,3.900498,3.7560349,3.6154766,3.4710135,3.330455,3.1859922,5.6535745,8.121157,10.588739,13.056321,15.523903,13.696643,11.869383,10.042123,8.214863,6.387602,6.0479193,5.708236,5.368553,5.02887,4.689187,7.0591593,9.4291315,11.799104,14.169076,16.539047,16.175938,15.812829,15.449719,15.086611,14.723501,20.146715,25.566027,30.985336,36.404648,41.823956,35.143524,28.466997,21.786564,15.1061325,8.4257,9.421323,10.413041,11.408664,12.404286,13.399908,14.118319,14.836729,15.551234,16.269644,16.988054,18.299932,19.611813,20.92369,22.23557,23.551353,28.080462,32.609566,37.138676,41.671684,46.20079,39.668728,33.140568,26.608501,20.080341,13.548276,12.084125,10.61607,9.148014,7.6799593,6.211904,11.404759,16.597614,21.790468,26.983324,32.176178,28.81449,25.456703,22.095013,18.733322,15.375536,12.44333,9.511124,6.578918,3.6467118,0.7106012,0.57785153,0.44119745,0.30844778,0.1717937,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.19522011,0.23816854,0.28502136,0.3318742,0.37482262,0.7262188,1.0815194,1.4329157,1.7843118,2.135708,3.5764325,5.017157,6.4578815,7.898606,9.339331,7.551114,5.7668023,3.9824903,2.1981785,0.41386664,1.0151446,1.6164225,2.2216048,2.822883,3.4241607,3.513962,3.6037633,3.6935644,3.7833657,3.873167,3.7599394,3.6467118,3.5295796,3.416352,3.2992198,2.639376,1.979532,1.319688,0.659844,0.0,0.48024148,0.96048295,1.4407244,1.9209659,2.4012074,2.3933985,2.3894942,2.3855898,2.3816853,2.3738766,2.592523,2.8111696,3.0259118,3.2445583,3.4632049,3.7794614,4.095718,4.415879,4.732136,5.0483923,4.123049,3.193801,2.2684577,1.33921,0.41386664,0.3318742,0.24597734,0.1639849,0.08199245,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13665408,0.26940376,0.40605783,0.5388075,0.6754616,0.92924774,1.1869383,1.4407244,1.6945106,1.9482968,2.8111696,3.6740425,4.5369153,5.3997884,6.262661,5.056201,3.8458362,2.639376,1.4329157,0.22645533,0.41386664,0.60518235,0.79649806,0.98390937,1.175225,0.97610056,0.78088045,0.58175594,0.38653582,0.18741131,0.42167544,0.6520352,0.8862993,1.116659,1.3509232,1.1127546,0.8745861,0.63641757,0.39824903,0.1639849,0.21474212,0.26940376,0.32016098,0.3709182,0.42557985,0.359205,0.29673457,0.23035973,0.1639849,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.093705654,0.14055848,0.19131571,0.23816854,0.26159495,0.28111696,0.30454338,0.3279698,0.3513962,0.42948425,0.5114767,0.58956474,0.6715572,0.74964523,0.679366,0.60518235,0.5309987,0.46071947,0.38653582,0.5192855,0.6481308,0.77697605,0.9058213,1.038571,0.94096094,0.8433509,0.74574083,0.6481308,0.5505207,0.45681506,0.359205,0.26549935,0.1717937,0.07418364,0.093705654,0.113227665,0.13665408,0.15617609,0.1756981,0.19131571,0.20693332,0.21864653,0.23426414,0.24988174,0.20693332,0.1639849,0.12103647,0.078088045,0.039044023,0.058566034,0.078088045,0.09761006,0.11713207,0.13665408,0.1717937,0.20693332,0.24207294,0.27721256,0.31235218,0.679366,1.0463798,1.4133936,1.7843118,2.1513257,1.9287747,1.7062237,1.4836729,1.261122,1.038571,0.94486535,0.8511597,0.76135844,0.6676528,0.57394713,0.6481308,0.7262188,0.80040246,0.8745861,0.94876975,1.3938715,1.8350691,2.2762666,2.7213683,3.1625657,3.0883822,3.0141985,2.9361105,2.8619268,2.787743,2.3894942,1.9912452,1.5969005,1.1986516,0.80040246,0.8589685,0.92143893,0.98000497,1.038571,1.1010414,1.0268579,0.94876975,0.8745861,0.80040246,0.7262188,0.74574083,0.76916724,0.79259366,0.8160201,0.8394465,0.8589685,0.8784905,0.8980125,0.91753453,0.93705654,0.9136301,0.8941081,0.8706817,0.8472553,0.8238289,0.79259366,0.76135844,0.7262188,0.6949836,0.6637484,0.698888,0.7340276,0.76916724,0.80430686,0.8394465,0.8316377,0.8238289,0.8160201,0.80821127,0.80040246,0.98390937,1.1635119,1.3470187,1.5305257,1.7140326,1.8233559,1.9365835,2.0498111,2.1630387,2.2762666,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.08980125,0.13665408,0.1796025,0.22645533,0.8706817,1.5149081,2.1591344,2.803361,3.4514916,5.263134,7.0786815,8.894228,10.709775,12.525322,13.376482,14.231546,15.0827055,15.933866,16.788929,17.01148,17.237936,17.460487,17.686943,17.913397,19.069101,20.228708,21.38441,22.544018,23.699722,23.35223,23.004738,22.657246,22.309755,21.962263,20.58401,19.205755,17.831406,16.453152,15.074897,13.8762455,12.67369,11.475039,10.276386,9.073831,10.990892,12.90405,14.821111,16.734268,18.651329,22.118439,25.589453,29.060467,32.53148,35.99859,38.33342,40.66435,42.999184,45.33011,47.661037,46.485813,45.31449,44.139267,42.964043,41.78882,44.553135,47.31745,50.081768,52.846085,55.614307,57.53527,59.456238,61.381107,63.302074,65.226944,65.1918,65.16057,65.12933,65.09419,65.06296,61.287403,57.511845,53.73629,49.96073,46.18908,46.107086,46.029,45.947006,45.86892,45.786926,41.54284,37.298756,33.050766,28.80668,24.562595,23.469362,22.372225,21.278992,20.181856,19.088623,19.717232,20.34584,20.978354,21.606962,22.239475,19.36193,16.484386,13.602938,10.729298,7.8517528,15.028045,22.204336,29.384531,36.56082,43.737114,36.533493,29.32987,22.122343,14.918721,7.7111945,6.356367,5.001539,3.6467118,2.2918842,0.93705654,2.4090161,3.8770714,5.349031,6.817086,8.289046,6.899079,5.5091114,4.1191444,2.7291772,1.33921,3.0337205,4.732136,6.4305506,8.128965,9.823476,10.366188,10.904996,11.443803,11.986515,12.525322,10.061645,7.5940623,5.1303844,2.6667068,0.19912452,2.2723622,4.3455997,6.4188375,8.488171,10.561408,8.449126,6.336845,4.224563,2.1122816,0.0,0.113227665,0.22645533,0.3357786,0.44900626,0.5622339,0.6949836,0.8277333,0.96048295,1.0932326,1.2259823,1.2533131,1.2845483,1.3157835,1.3431144,1.3743496,1.8858263,2.4012074,2.912684,3.4241607,3.9356375,4.009821,4.084005,4.154284,4.2284675,4.298747,4.7243266,5.1460023,5.5676775,5.989353,6.4110284,5.6535745,4.8961205,4.138666,3.3812122,2.6237583,5.8878384,9.148014,12.412095,15.676175,18.936352,15.176412,11.412568,7.648724,3.8887846,0.12494087,0.21083772,0.30063897,0.38653582,0.47633708,0.5622339,2.096664,3.631094,5.169429,6.703859,8.238289,7.570636,6.9068875,6.2431393,5.579391,4.911738,4.950782,4.985922,5.024966,5.0640097,5.099149,4.3260775,3.5569105,2.7838387,2.0107672,1.2376955,1.0424755,0.8472553,0.6520352,0.45681506,0.26159495,1.3782539,2.4988174,3.6154766,4.732136,5.8487945,5.1303844,4.4119744,3.68966,2.97125,2.2489357,5.056201,7.8634663,10.670732,13.481901,16.289165,14.688361,13.091461,11.49456,9.897659,8.300759,7.941554,7.578445,7.2192397,6.860035,6.5008297,8.781001,11.061172,13.341343,15.621513,17.901684,17.7377,17.573715,17.413633,17.24965,17.085665,22.5284,27.971138,33.413876,38.856613,44.299347,37.228474,30.161507,23.090635,16.019762,8.94889,10.280292,11.611692,12.939189,14.27059,15.601992,16.30869,17.015385,17.722082,18.42878,19.13938,18.90121,18.663042,18.424873,18.186707,17.948538,22.020828,26.089216,30.161507,34.229893,38.298283,33.82774,29.361105,24.890564,20.420023,15.949483,13.817679,11.685876,9.554072,7.4183645,5.2865605,11.568744,17.850927,24.137014,30.419197,36.70138,32.24646,27.795439,23.340517,18.889498,14.438479,11.642927,8.85128,6.0596323,3.2679846,0.47633708,0.38653582,0.29673457,0.20693332,0.113227665,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.031235218,0.06637484,0.09761006,0.12884527,0.1639849,0.20693332,0.24597734,0.28892577,0.3318742,0.37482262,0.9097257,1.4446288,1.979532,2.514435,3.049338,3.697469,4.3455997,4.9937305,5.6418614,6.2860875,5.1460023,4.0059166,2.8658314,1.7257458,0.58566034,1.1986516,1.8077383,2.416825,3.0259118,3.638903,3.5608149,3.4827268,3.4046388,3.3265507,3.2484627,3.0415294,2.8306916,2.619854,2.4090161,2.1981785,1.7608855,1.319688,0.8784905,0.44119745,0.0,0.32016098,0.64032197,0.96048295,1.2806439,1.6008049,1.6437533,1.6867018,1.7257458,1.7686942,1.8116426,2.182561,2.5534792,2.9243972,3.2914112,3.6623292,4.0059166,4.3534083,4.6969957,5.040583,5.388075,4.365122,3.3421683,2.3192148,1.2962615,0.27330816,0.21864653,0.1639849,0.10932326,0.05466163,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08980125,0.1796025,0.26940376,0.359205,0.44900626,0.62079996,0.78868926,0.96048295,1.1283722,1.3001659,1.8741131,2.4480603,3.0259118,3.5998588,4.173806,3.408543,2.639376,1.8741131,1.1049459,0.3357786,0.62079996,0.9058213,1.1908426,1.475864,1.7608855,1.43682,1.1088502,0.78088045,0.45291066,0.12494087,0.28111696,0.43338865,0.58956474,0.74574083,0.9019169,0.74964523,0.60127795,0.44900626,0.30063897,0.14836729,0.1835069,0.21864653,0.25378615,0.28892577,0.3240654,0.27721256,0.23035973,0.1835069,0.13665408,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.21474212,0.23035973,0.24597734,0.26159495,0.27330816,0.3318742,0.39044023,0.44900626,0.5036679,0.5622339,0.5231899,0.48414588,0.44119745,0.40215343,0.3631094,0.4958591,0.62860876,0.76135844,0.8941081,1.0268579,0.94876975,0.8706817,0.79259366,0.7145056,0.63641757,0.5309987,0.42557985,0.3240654,0.21864653,0.113227665,0.14055848,0.1717937,0.20302892,0.23426414,0.26159495,0.27330816,0.28111696,0.29283017,0.30063897,0.31235218,0.25378615,0.19912452,0.14055848,0.08199245,0.023426414,0.042948425,0.058566034,0.078088045,0.093705654,0.113227665,0.1639849,0.21864653,0.26940376,0.3240654,0.37482262,0.75745404,1.1400855,1.5227169,1.9053483,2.2879796,2.0459068,1.8077383,1.5656652,1.3274968,1.0893283,0.96829176,0.8472553,0.7262188,0.60908675,0.48805028,0.61299115,0.737932,0.8628729,0.9878138,1.1127546,1.6437533,2.1786566,2.7096553,3.240654,3.775557,3.8106966,3.8497405,3.8887846,3.9239242,3.9629683,3.3616903,2.7565079,2.15523,1.5539521,0.94876975,0.96438736,0.98000497,0.9956226,1.0112402,1.0268579,0.96438736,0.9019169,0.8394465,0.77307165,0.7106012,0.7262188,0.7418364,0.75745404,0.77307165,0.78868926,0.79259366,0.79649806,0.80430686,0.80821127,0.81211567,0.80821127,0.80821127,0.80430686,0.80430686,0.80040246,0.79649806,0.78868926,0.78478485,0.78088045,0.77307165,0.8277333,0.8784905,0.93315214,0.98390937,1.038571,1.0190489,1.0034313,0.98390937,0.96829176,0.94876975,1.1674163,1.3860629,1.6008049,1.8194515,2.0380979,2.135708,2.2372224,2.338737,2.436347,2.5378613,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.093705654,0.14055848,0.19131571,0.23816854,0.7340276,1.2337911,1.7296503,2.2294137,2.7252727,4.657952,6.590631,8.52331,10.455989,12.388668,12.6463585,12.90405,13.16174,13.415526,13.673217,14.063657,14.450192,14.836729,15.223265,15.613705,17.409729,19.205755,21.005684,22.801708,24.601639,24.332235,24.066736,23.79733,23.531832,23.262428,21.528873,19.799223,18.06567,16.332115,14.59856,13.462379,12.326198,11.186112,10.049932,8.913751,11.568744,14.227642,16.88654,19.541533,22.200432,25.648018,29.095606,32.543194,35.99078,39.438366,42.023083,44.607796,47.19251,49.777225,52.36194,52.12377,51.889507,51.651337,51.41317,51.175,52.15891,53.138916,54.122826,55.106735,56.08674,58.480137,60.873535,63.266933,65.656425,68.04983,67.65158,67.25333,66.858986,66.46073,66.062485,61.088276,56.11407,51.135956,46.161747,41.18754,42.085552,42.983566,43.881577,44.775684,45.6737,41.816147,37.954693,34.09324,30.235691,26.374237,25.24196,24.10578,22.969599,21.833418,20.701141,21.15405,21.603058,22.05597,22.508879,22.96179,19.178425,15.398962,11.615597,7.832231,4.0488653,14.344774,24.640682,34.936592,45.228596,55.524506,46.28669,37.044968,27.80325,18.565434,9.323712,7.6838636,6.044015,4.4041657,2.7643168,1.1244678,1.999054,2.8697357,3.7443218,4.6150036,5.4856853,4.5408196,3.5959544,2.6510892,1.7062237,0.76135844,1.6164225,2.4714866,3.3265507,4.181615,5.036679,5.282656,5.5286336,5.7707067,6.016684,6.262661,5.02887,3.7989833,2.5651922,1.3314011,0.10151446,1.1439898,2.1864653,3.2289407,4.271416,5.3138914,4.251894,3.1859922,2.1239948,1.0619974,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.5114767,0.6442264,0.78088045,0.9136301,1.0502841,1.2025559,1.3548276,1.5070993,1.6593709,1.8116426,2.260649,2.7135596,3.1625657,3.611572,4.0605783,4.2440853,4.423688,4.60329,4.7828927,4.9624953,4.8687897,4.7711797,4.677474,4.5837684,4.4861584,4.0020123,3.5178664,3.0337205,2.5456703,2.0615244,3.611572,5.1616197,6.7116675,8.261715,9.811763,7.8751793,5.938596,3.998108,2.0615244,0.12494087,0.21083772,0.30063897,0.38653582,0.47633708,0.5622339,1.4172981,2.2723622,3.1274261,3.9824903,4.8375545,5.181142,5.520825,5.8644123,6.2079997,6.551587,6.0518236,5.548156,5.0483923,4.548629,4.0488653,3.5686235,3.0883822,2.6081407,2.1318035,1.6515622,1.3899672,1.1283722,0.8706817,0.60908675,0.3513962,1.8389735,3.330455,4.8219366,6.309514,7.800996,6.5008297,5.2045684,3.9083066,2.6081407,1.3118792,4.4588275,7.605776,10.756628,13.903577,17.050524,15.683984,14.313539,12.946998,11.580457,10.213917,9.8312845,9.452558,9.073831,8.691199,8.312472,10.502842,12.693212,14.883581,17.073952,19.26432,19.29946,19.338505,19.373644,19.412687,19.451733,24.91399,30.380154,35.846317,41.308575,46.77474,39.313427,31.856018,24.394705,16.933393,9.475985,11.139259,12.806439,14.469715,16.136894,17.800169,18.499058,19.194042,19.89293,20.591818,21.2868,19.498585,17.714273,15.926057,14.13784,12.349625,15.961197,19.568865,23.180437,26.788103,30.399675,27.99066,25.581644,23.168722,20.759706,18.35069,15.551234,12.755682,9.956225,7.1606736,4.3612175,11.736633,19.108145,26.479656,33.851166,41.22658,35.67843,30.134176,24.589926,19.045673,13.501423,10.84643,8.19534,5.5442514,2.8892577,0.23816854,0.19131571,0.14836729,0.10151446,0.058566034,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.21474212,0.25378615,0.29673457,0.3357786,0.37482262,1.0932326,1.8116426,2.5261483,3.2445583,3.9629683,3.8185053,3.6740425,3.5256753,3.3812122,3.2367494,2.7408905,2.2489357,1.7530766,1.2572175,0.76135844,1.3782539,1.999054,2.6159496,3.232845,3.8497405,3.6037633,3.3616903,3.1157131,2.8697357,2.6237583,2.3192148,2.0146716,1.7101282,1.4055848,1.1010414,0.8784905,0.659844,0.44119745,0.21864653,0.0,0.16008049,0.32016098,0.48024148,0.64032197,0.80040246,0.8902037,0.98000497,1.0698062,1.1596074,1.2494087,1.7725986,2.2957885,2.8189783,3.338264,3.8614538,4.2362766,4.607195,4.9781127,5.3529353,5.7238536,4.607195,3.4905357,2.3738766,1.2533131,0.13665408,0.10932326,0.08199245,0.05466163,0.027330816,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.08980125,0.13665408,0.1796025,0.22645533,0.30844778,0.39434463,0.48024148,0.5661383,0.6481308,0.93705654,1.2259823,1.5110037,1.7999294,2.0888553,1.7608855,1.4329157,1.1049459,0.77697605,0.44900626,0.8316377,1.2103647,1.5890918,1.9717231,2.35045,1.893635,1.43682,0.97610056,0.5192855,0.062470436,0.14055848,0.21864653,0.29673457,0.3709182,0.44900626,0.38653582,0.3240654,0.26159495,0.19912452,0.13665408,0.15617609,0.1717937,0.19131571,0.20693332,0.22645533,0.19522011,0.1639849,0.13665408,0.10541886,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.06637484,0.09761006,0.12884527,0.1639849,0.1717937,0.1756981,0.1835069,0.19131571,0.19912452,0.23426414,0.26940376,0.30454338,0.339683,0.37482262,0.3670138,0.359205,0.3513962,0.3435874,0.3357786,0.47243267,0.60908675,0.7418364,0.8784905,1.0112402,0.95657855,0.8980125,0.8394465,0.78088045,0.7262188,0.60908675,0.4958591,0.37872702,0.26549935,0.14836729,0.19131571,0.23035973,0.26940376,0.30844778,0.3513962,0.3553006,0.359205,0.3631094,0.3709182,0.37482262,0.30063897,0.23035973,0.15617609,0.08589685,0.011713207,0.027330816,0.042948425,0.058566034,0.07418364,0.08589685,0.15617609,0.22645533,0.29673457,0.3670138,0.43729305,0.8355421,1.2337911,1.6281357,2.0263848,2.4246337,2.1669433,1.9092526,1.6515622,1.3938715,1.1361811,0.9917182,0.8433509,0.6949836,0.5466163,0.39824903,0.57394713,0.74964523,0.92534333,1.1010414,1.2767396,1.8975395,2.5183394,3.1430438,3.7638438,4.388548,4.5369153,4.689187,4.8375545,4.985922,5.138193,4.3299823,3.521771,2.7135596,1.9092526,1.1010414,1.0698062,1.038571,1.0112402,0.98000497,0.94876975,0.9019169,0.8511597,0.80040246,0.74964523,0.698888,0.7066968,0.7145056,0.7223144,0.7301232,0.737932,0.7262188,0.71841,0.7066968,0.698888,0.6871748,0.7066968,0.7223144,0.7418364,0.75745404,0.77307165,0.79649806,0.8199245,0.8433509,0.8667773,0.8862993,0.95657855,1.0268579,1.097137,1.1674163,1.2376955,1.2103647,1.183034,1.1557031,1.1283722,1.1010414,1.3509232,1.6047094,1.8584955,2.1083772,2.3621633,2.4480603,2.5378613,2.6237583,2.7135596,2.7994564,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.60127795,0.94876975,1.3001659,1.6515622,1.999054,4.0488653,6.098676,8.148487,10.198298,12.24811,11.912332,11.576552,11.23687,10.901091,10.561408,11.111929,11.66245,12.212971,12.763491,13.314012,15.750359,18.186707,20.626957,23.063305,25.499651,25.31224,25.124828,24.937418,24.750006,24.562595,22.47374,20.388788,18.299932,16.211079,14.126127,13.048512,11.974802,10.901091,9.823476,8.749765,12.150499,15.551234,18.95197,22.348799,25.749533,29.173695,32.601757,36.02592,39.45008,42.87424,45.71274,48.551243,51.385838,54.22434,57.06284,57.761726,58.460613,59.163406,59.862297,60.561184,59.76078,58.964283,58.16388,57.36348,56.563076,59.425003,62.28693,65.14886,68.01078,70.87662,70.11135,69.34999,68.58863,67.82337,67.06201,60.889153,54.712387,48.535625,42.362766,36.186,38.06402,39.93813,41.812244,43.686356,45.564373,42.089455,38.61454,35.135715,31.660797,28.18588,27.010654,25.839334,24.664108,23.488884,22.31366,22.586967,22.86418,23.137487,23.410795,23.68801,18.998821,14.313539,9.6243515,4.939069,0.24988174,13.661504,27.073126,40.48865,53.900272,67.3119,56.03598,44.763973,33.48806,22.212145,10.936231,9.01136,7.08649,5.1616197,3.2367494,1.3118792,1.5890918,1.8623998,2.135708,2.4129205,2.6862288,2.1864653,1.6867018,1.1869383,0.6871748,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.3240654,0.46071947,0.60127795,0.737932,0.8745861,1.1517987,1.4251068,1.698415,1.9756275,2.2489357,2.639376,3.0259118,3.4124475,3.7989833,4.1894236,4.474445,4.7633705,5.0483923,5.337318,5.6262436,5.0132523,4.4002614,3.78727,3.174279,2.5612879,2.35045,2.135708,1.9248703,1.7140326,1.4992905,1.33921,1.175225,1.0112402,0.8511597,0.6871748,0.57394713,0.46071947,0.3513962,0.23816854,0.12494087,0.21083772,0.30063897,0.38653582,0.47633708,0.5622339,0.737932,0.9136301,1.0893283,1.261122,1.43682,2.787743,4.138666,5.4856853,6.8366084,8.187531,7.1489606,6.114294,5.0757227,4.037152,2.998581,2.8111696,2.6237583,2.436347,2.2489357,2.0615244,1.737459,1.4133936,1.0893283,0.76135844,0.43729305,2.2996929,4.1620927,6.0244927,7.8868923,9.749292,7.8751793,6.001066,4.123049,2.2489357,0.37482262,3.8614538,7.348085,10.838621,14.325252,17.811884,16.675701,15.535617,14.399435,13.263254,12.123169,11.72492,11.326671,10.924518,10.526268,10.124115,12.224684,14.325252,16.42582,18.526388,20.623053,20.861221,21.09939,21.337559,21.575727,21.813896,27.29958,32.78917,38.274857,43.764446,49.25013,41.398376,33.55053,25.698776,17.850927,9.999174,11.998228,14.001186,16.00024,17.999294,19.998348,20.689428,21.376602,22.063778,22.750952,23.438128,20.099863,16.761599,13.423335,10.088976,6.7507114,9.901564,13.048512,16.199366,19.350218,22.50107,22.149673,21.798277,21.450787,21.09939,20.751898,17.288692,13.825488,10.362284,6.899079,3.435874,11.900618,20.361458,28.826202,37.28704,45.751785,39.110397,32.476818,25.83543,19.20185,12.564366,10.049932,7.5394006,5.024966,2.5105307,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.22645533,0.26159495,0.30063897,0.3357786,0.37482262,1.2767396,2.174752,3.076669,3.9746814,4.8765984,3.9356375,2.998581,2.0615244,1.1244678,0.18741131,0.3357786,0.48805028,0.63641757,0.78868926,0.93705654,1.5617609,2.1864653,2.8111696,3.435874,4.0605783,3.6506162,3.2367494,2.8267872,2.4129205,1.999054,1.6008049,1.1986516,0.80040246,0.39824903,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13665408,0.27330816,0.41386664,0.5505207,0.6871748,1.3626363,2.0380979,2.7135596,3.3890212,4.0605783,4.462732,4.860981,5.263134,5.661383,6.0635366,4.8492675,3.638903,2.4246337,1.2142692,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.113227665,0.22645533,0.3357786,0.44900626,0.5622339,1.038571,1.5110037,1.9873407,2.463678,2.9361105,2.35045,1.7608855,1.175225,0.58566034,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.21083772,0.23816854,0.26159495,0.28892577,0.31235218,0.44900626,0.58566034,0.7262188,0.8628729,0.999527,0.96438736,0.92534333,0.8862993,0.8511597,0.81211567,0.6871748,0.5622339,0.43729305,0.31235218,0.18741131,0.23816854,0.28892577,0.3357786,0.38653582,0.43729305,0.43729305,0.43729305,0.43729305,0.43729305,0.43729305,0.3513962,0.26159495,0.1756981,0.08589685,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.14836729,0.23816854,0.3240654,0.41386664,0.4997635,0.9136301,1.3235924,1.737459,2.1513257,2.5612879,2.2879796,2.0107672,1.737459,1.4641509,1.1869383,1.0112402,0.8394465,0.6637484,0.48805028,0.31235218,0.5388075,0.76135844,0.9878138,1.2142692,1.43682,2.1513257,2.8619268,3.5764325,4.2870336,5.001539,5.263134,5.5247293,5.786324,6.0518236,6.3134184,5.298274,4.2870336,3.2757936,2.260649,1.2494087,1.175225,1.1010414,1.0268579,0.94876975,0.8745861,0.8394465,0.80040246,0.76135844,0.7262188,0.6871748,0.6871748,0.6871748,0.6871748,0.6871748,0.6871748,0.6637484,0.63641757,0.61299115,0.58566034,0.5622339,0.60127795,0.63641757,0.6754616,0.7106012,0.74964523,0.80040246,0.8511597,0.9019169,0.94876975,0.999527,1.0893283,1.175225,1.261122,1.3509232,1.43682,1.4016805,1.3626363,1.3235924,1.2884527,1.2494087,1.5383345,1.8233559,2.1122816,2.4012074,2.6862288,2.7643168,2.8385005,2.912684,2.9868677,3.0610514,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.14836729,0.25769055,0.3670138,0.47633708,0.58566034,0.97610056,1.3626363,1.7491722,2.135708,2.5261483,4.1972322,5.8683167,7.5433054,9.21439,10.889378,10.741011,10.592644,10.444276,10.295909,10.151445,10.530173,10.9089,11.291532,11.6702585,12.0489855,14.161267,16.273548,18.38583,20.502016,22.614298,22.508879,22.40346,22.29804,22.192623,22.087204,20.486399,18.88169,17.280884,15.676175,14.07537,13.189071,12.306676,11.420377,10.534078,9.651682,12.4745655,15.3013525,18.124235,20.951023,23.773905,26.955994,30.134176,33.316265,36.49445,39.676537,41.710728,43.744923,45.779118,47.81331,49.85141,50.27699,50.70647,51.132053,51.561535,51.987118,50.6401,49.29308,47.94606,46.59904,45.25202,48.039764,50.831413,53.619156,56.410805,59.198547,59.49528,59.792015,60.084846,60.38158,60.67441,55.49327,50.316032,45.13489,39.953747,34.776512,35.904884,37.033257,38.16553,39.293903,40.42618,40.738533,41.050884,41.36324,41.67559,41.98794,37.228474,32.47291,27.713448,22.957886,18.19842,18.420969,18.639616,18.858263,19.080814,19.29946,15.601992,11.900618,8.1992445,4.5017757,0.80040246,11.408664,22.020828,32.62909,43.241257,53.849518,44.838154,35.826794,26.811531,17.800169,8.78881,7.523783,6.2587566,4.9937305,3.7287042,2.463678,2.4012074,2.338737,2.2762666,2.2137961,2.1513257,2.0068626,1.8584955,1.7140326,1.5695697,1.4251068,1.5617609,1.698415,1.8389735,1.9756275,2.1122816,2.4090161,2.7018464,2.998581,3.2914112,3.5881457,2.9439192,2.3035975,1.6593709,1.0190489,0.37482262,0.30844778,0.24597734,0.1796025,0.113227665,0.05075723,0.042948425,0.03513962,0.027330816,0.019522011,0.011713207,0.05075723,0.08589685,0.12494087,0.1639849,0.19912452,0.30844778,0.41386664,0.5231899,0.62860876,0.737932,1.43682,2.1318035,2.8306916,3.5256753,4.224563,4.056674,3.8887846,3.7208953,3.5569105,3.3890212,3.677947,3.9668727,4.2557983,4.548629,4.8375545,4.298747,3.7638438,3.2250361,2.6862288,2.1513257,1.9639144,1.7804074,1.5969005,1.4094892,1.2259823,1.0932326,0.96438736,0.8355421,0.7066968,0.57394713,0.48024148,0.38653582,0.28892577,0.19522011,0.10151446,0.21083772,0.32016098,0.42948425,0.5388075,0.6481308,1.0346665,1.4212024,1.8038338,2.1903696,2.5769055,3.3929255,4.2089458,5.02887,5.84489,6.66091,5.8097506,4.958591,4.1035266,3.252367,2.4012074,2.436347,2.4714866,2.5066261,2.541766,2.5769055,2.1396124,1.7062237,1.2689307,0.8355421,0.39824903,2.096664,3.7911747,5.4856853,7.180196,8.874706,7.9220324,6.969358,6.016684,5.0640097,4.1113358,6.348558,8.581876,10.819098,13.052417,15.285735,14.176885,13.06413,11.951375,10.838621,9.725866,9.6673,9.608734,9.554072,9.495506,9.43694,10.9089,12.380859,13.856724,15.328683,16.800642,16.95682,17.10909,17.265266,17.421442,17.573715,22.579159,27.580698,32.582237,37.583775,42.58922,36.228947,29.868677,23.508406,17.148134,10.787864,12.2793455,13.766922,15.258404,16.745981,18.237463,18.8036,19.373644,19.939783,20.50592,21.075964,18.303837,15.535617,12.763491,9.99527,7.223144,10.826907,14.426766,18.026625,21.626484,25.226343,26.179018,27.131691,28.084366,29.033134,29.98581,25.222439,20.459068,15.6917925,10.928422,6.1611466,12.603411,19.041769,25.484034,31.922394,38.360752,33.050766,27.744682,22.430792,17.120804,11.810817,9.753197,7.6916723,5.6340523,3.5725281,1.5110037,1.2103647,0.9058213,0.60518235,0.30063897,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.042948425,0.08589685,0.12884527,0.1717937,0.21083772,0.23426414,0.25378615,0.27330816,0.29283017,0.31235218,1.077615,1.8428779,2.6081407,3.3734035,4.138666,3.6428072,3.1469483,2.6510892,2.1591344,1.6632754,1.4797685,1.2962615,1.116659,0.93315214,0.74964523,1.3860629,2.0263848,2.6628022,3.2992198,3.9356375,3.611572,3.2836022,2.9556324,2.6276627,2.2996929,2.0341935,1.7686942,1.5031948,1.2415999,0.97610056,0.78088045,0.58566034,0.39044023,0.19522011,0.0,0.0,0.0,0.0,0.0,0.0,0.1639849,0.3240654,0.48805028,0.6481308,0.81211567,1.3509232,1.893635,2.4324427,2.97125,3.513962,3.8458362,4.1777105,4.5095844,4.841459,5.173333,4.138666,3.1039999,2.069333,1.0346665,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.44510186,0.8902037,1.3353056,1.7804074,2.2255092,1.7804074,1.3353056,0.8902037,0.44510186,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.093705654,0.19131571,0.28502136,0.37872702,0.47633708,0.8511597,1.2298868,1.6086137,1.9834363,2.3621633,1.8897307,1.4172981,0.94486535,0.47243267,0.0,0.0,0.0,0.0,0.0,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.12884527,0.12103647,0.113227665,0.10932326,0.10151446,0.093705654,0.08980125,0.08589685,0.078088045,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.10151446,0.10541886,0.10932326,0.10932326,0.113227665,0.12103647,0.12884527,0.13665408,0.14055848,0.14836729,0.1756981,0.19912452,0.22645533,0.24988174,0.27330816,0.38653582,0.4997635,0.61299115,0.7262188,0.8394465,0.8433509,0.8511597,0.8589685,0.8667773,0.8745861,0.77697605,0.679366,0.58175594,0.48414588,0.38653582,0.44119745,0.4958591,0.5544251,0.60908675,0.6637484,0.6637484,0.6637484,0.6637484,0.6637484,0.6637484,0.5661383,0.46852827,0.3709182,0.27330816,0.1756981,0.15617609,0.13665408,0.113227665,0.093705654,0.07418364,0.14836729,0.21864653,0.29283017,0.3631094,0.43729305,0.8667773,1.2962615,1.7257458,2.1591344,2.5886188,2.2840753,1.9756275,1.6710842,1.3665408,1.0619974,0.9097257,0.75745404,0.60518235,0.45291066,0.30063897,0.5231899,0.74574083,0.96829176,1.1908426,1.4133936,2.0927596,2.7721257,3.4514916,4.1308575,4.814128,4.9663997,5.1186714,5.270943,5.423215,5.575486,4.8492675,4.123049,3.4007344,2.6745155,1.9482968,1.9209659,1.893635,1.8663043,1.8389735,1.8116426,1.6359446,1.4641509,1.2884527,1.1127546,0.93705654,0.8902037,0.8433509,0.79649806,0.74574083,0.698888,0.6715572,0.6442264,0.61689556,0.58956474,0.5622339,0.58566034,0.60908675,0.62860876,0.6520352,0.6754616,0.7145056,0.75354964,0.79649806,0.8355421,0.8745861,0.94876975,1.0190489,1.0932326,1.1635119,1.2376955,1.2337911,1.2337911,1.2298868,1.2259823,1.2259823,1.475864,1.7257458,1.9756275,2.2255092,2.475391,2.7213683,2.97125,3.2172275,3.4632049,3.7130866,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.24597734,0.41386664,0.58566034,0.75354964,0.92534333,1.3509232,1.7765031,2.1981785,2.6237583,3.049338,4.3455997,5.6418614,6.9342184,8.23048,9.526741,9.565785,9.608734,9.651682,9.694631,9.737579,9.948417,10.159255,10.366188,10.577025,10.787864,12.576079,14.364296,16.148607,17.936825,5052.0,19.701614,19.678188,19.658665,19.635239,19.611813,18.495153,17.378494,16.261835,15.141272,14.024612,13.329629,12.634645,11.939662,11.2446785,10.549695,12.798631,15.051471,17.300406,19.549341,21.798277,24.734388,27.670498,30.60661,33.538815,36.474926,37.708717,38.938602,40.172394,41.406185,42.636074,42.792248,42.948425,43.100697,43.256874,43.413048,41.519413,39.621876,37.728237,35.8307,33.937065,36.65453,39.371994,42.089455,44.80692,47.524384,48.87921,50.230137,51.58106,52.935886,54.286808,50.101288,45.91577,41.734158,37.548637,33.363117,33.74575,34.132286,34.51882,34.90145,35.287987,39.38761,43.487232,47.586853,51.686478,55.7861,47.446297,39.10649,30.76669,22.426888,14.087084,14.251068,14.418958,14.582942,14.746927,14.9109125,12.201257,9.487698,6.774138,4.0605783,1.3509232,9.155824,16.964628,24.773432,32.57833,40.38714,33.636425,26.885714,20.138906,13.388195,6.6374836,6.0323014,5.4271193,4.8219366,4.2167544,3.611572,3.213323,2.8111696,2.4129205,2.0107672,1.6125181,1.8233559,2.0341935,2.241127,2.4519646,2.6628022,2.9243972,3.1859922,3.4514916,3.7130866,3.9746814,4.6150036,5.2553253,5.8956475,6.5359693,7.1762915,5.891743,4.60329,3.3187418,2.0341935,0.74964523,0.60908675,0.46462387,0.3240654,0.1796025,0.039044023,0.03513962,0.031235218,0.031235218,0.027330816,0.023426414,0.062470436,0.10151446,0.13665408,0.1756981,0.21083772,0.28892577,0.3670138,0.44510186,0.5231899,0.60127795,1.7218413,2.8385005,3.959064,5.0796275,6.2001905,5.477876,4.755562,4.0332475,3.310933,2.5886188,2.8814487,3.174279,3.4632049,3.7560349,4.0488653,3.5881457,3.1235218,2.6628022,2.1981785,1.737459,1.5812829,1.4212024,1.2650263,1.1088502,0.94876975,0.8511597,0.75354964,0.6559396,0.5583295,0.46071947,0.38653582,0.30844778,0.23035973,0.15227169,0.07418364,0.20693332,0.339683,0.47243267,0.60518235,0.737932,1.3314011,1.9287747,2.522244,3.1157131,3.7130866,3.998108,4.283129,4.5681505,4.853172,5.138193,4.4705405,3.802888,3.135235,2.4675822,1.7999294,2.05762,2.3153105,2.5730011,2.8306916,3.0883822,2.541766,1.999054,1.4524376,0.9058213,0.3631094,1.8897307,3.416352,4.9468775,6.473499,8.00012,7.968885,7.941554,7.910319,7.8790836,7.8517528,8.831758,9.815667,10.795672,11.779582,12.763491,11.674163,10.588739,9.499411,8.413987,7.3246584,7.60968,7.8947015,8.179723,8.464745,8.749765,9.593117,10.4403715,11.283723,12.130978,12.974329,13.048512,13.118792,13.192975,13.263254,13.337439,17.854832,22.372225,26.889618,31.407011,35.924404,31.055616,26.186827,21.314133,16.445343,11.576552,12.556558,13.536563,14.516567,15.4965725,16.476578,16.921679,17.370686,17.815788,18.264793,18.7138,16.511717,14.30573,12.103647,9.901564,7.699481,11.748346,15.801116,19.849981,23.898846,27.951616,30.204456,32.4612,34.71404,36.970783,39.223625,33.156185,27.088743,21.021301,14.95386,8.886419,13.306203,17.722082,22.141865,26.557745,30.973623,26.991133,23.008642,19.026152,15.043662,11.061172,9.456462,7.8478484,6.239235,4.630621,3.0259118,2.4207294,1.815547,1.2103647,0.60518235,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.093705654,0.14055848,0.19131571,0.23816854,0.23816854,0.24207294,0.24597734,0.24597734,0.24988174,0.8784905,1.5110037,2.1396124,2.7682211,3.4007344,3.3460727,3.2953155,3.240654,3.1898966,3.1391394,2.6237583,2.1083772,1.5929961,1.077615,0.5622339,1.2142692,1.8623998,2.514435,3.1625657,3.8106966,3.5686235,3.3265507,3.084478,2.8424048,2.6003318,2.4714866,2.338737,2.2098918,2.0810463,1.9482968,1.5617609,1.1713207,0.78088045,0.39044023,0.0,0.0,0.0,0.0,0.0,0.0,0.18741131,0.37482262,0.5622339,0.74964523,0.93705654,1.3431144,1.7491722,2.1513257,2.5573835,2.9634414,3.2289407,3.4905357,3.7560349,4.0215344,4.2870336,3.4280653,2.5730011,1.7140326,0.8589685,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.8902037,1.7804074,2.6706111,3.5608149,4.4510183,3.5608149,2.6706111,1.7804074,0.8902037,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.078088045,0.15617609,0.23426414,0.30844778,0.38653582,0.6676528,0.94876975,1.2259823,1.5070993,1.7882162,1.4290112,1.0737107,0.7145056,0.359205,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.13665408,0.12103647,0.10541886,0.08980125,0.07418364,0.078088045,0.078088045,0.08199245,0.08589685,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.078088045,0.08589685,0.08980125,0.093705654,0.10151446,0.10151446,0.10541886,0.10932326,0.10932326,0.113227665,0.13665408,0.1639849,0.18741131,0.21083772,0.23816854,0.3240654,0.41386664,0.4997635,0.58566034,0.6754616,0.7262188,0.78088045,0.8316377,0.8862993,0.93705654,0.8667773,0.79649806,0.7262188,0.6559396,0.58566034,0.6481308,0.7066968,0.76916724,0.8277333,0.8862993,0.8862993,0.8862993,0.8862993,0.8862993,0.8862993,0.78088045,0.6715572,0.5661383,0.45681506,0.3513962,0.29673457,0.24597734,0.19131571,0.14055848,0.08589685,0.14446288,0.20302892,0.26159495,0.31625658,0.37482262,0.8238289,1.2689307,1.717937,2.1630387,2.612045,2.2762666,1.9443923,1.6086137,1.2728351,0.93705654,0.80821127,0.679366,0.5466163,0.41777104,0.28892577,0.5075723,0.7262188,0.94876975,1.1674163,1.3860629,2.0341935,2.6823244,3.330455,3.978586,4.6267166,4.6657605,4.7087092,4.7516575,4.794606,4.8375545,4.4002614,3.9629683,3.5256753,3.0883822,2.6510892,2.6706111,2.690133,2.7096553,2.7291772,2.7486992,2.436347,2.1239948,1.8116426,1.4992905,1.1869383,1.0932326,0.9956226,0.9019169,0.80821127,0.7106012,0.6832704,0.6520352,0.62079996,0.59346914,0.5622339,0.5700427,0.57785153,0.58566034,0.59346914,0.60127795,0.62860876,0.659844,0.6910792,0.71841,0.74964523,0.80821127,0.8667773,0.92143893,0.98000497,1.038571,1.0698062,1.1010414,1.1361811,1.1674163,1.1986516,1.4133936,1.6242313,1.8389735,2.0498111,2.260649,2.6823244,3.1039999,3.521771,3.9434462,4.3612175,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.3435874,0.57394713,0.80430686,1.0307622,1.261122,1.7257458,2.1864653,2.6510892,3.1118085,3.5764325,4.493967,5.4115014,6.329036,7.2465706,8.164105,8.3944645,8.628729,8.859089,9.093353,9.323712,9.366661,9.405705,9.444749,9.483793,9.526741,10.986988,12.4511385,13.911386,15.375536,16.835783,16.898252,16.95682,17.019289,17.077856,17.136421,16.503908,15.871395,15.238882,14.606369,13.973856,13.470188,12.96652,12.458947,11.955279,11.4516115,13.1266,14.801589,16.476578,18.151566,19.826555,22.516687,25.202917,27.89305,30.583183,33.273315,33.706703,34.13619,34.565674,34.99516,35.42464,35.30751,35.190376,35.073246,34.956112,34.83898,32.394825,29.95067,27.510418,25.066263,22.62601,25.26929,27.916475,30.559757,33.203037,35.85022,38.25924,40.668255,43.081173,45.490192,47.899208,44.70931,41.519413,38.329517,35.13962,31.949724,31.590519,31.231314,30.868204,30.508999,30.149794,38.036686,45.92358,53.814377,61.701267,69.58816,57.664116,45.743977,33.81993,21.895887,9.975748,10.085071,10.194394,10.303718,10.413041,10.526268,8.800523,7.0747766,5.349031,3.6232853,1.901444,6.902983,11.908427,16.91387,21.919313,26.924759,22.4386,17.948538,13.462379,8.976221,4.4861584,4.5408196,4.5993857,4.6540475,4.7087092,4.7633705,4.025439,3.2875066,2.5495746,1.8116426,1.0737107,1.639849,2.2059872,2.7682211,3.3343596,3.900498,4.2870336,4.6735697,5.0640097,5.4505453,5.8370814,6.8209906,7.8088045,8.792714,9.776623,10.764437,8.835662,6.9068875,4.9781127,3.0532427,1.1244678,0.9058213,0.6832704,0.46462387,0.24597734,0.023426414,0.027330816,0.031235218,0.031235218,0.03513962,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.22645533,0.27330816,0.32016098,0.3670138,0.41386664,0.46071947,2.0068626,3.5491016,5.0913405,6.6335793,8.175818,6.899079,5.618435,4.3416953,3.0649557,1.7882162,2.0810463,2.377781,2.6706111,2.9673457,3.2640803,2.87364,2.4871042,2.1005683,1.7140326,1.3235924,1.1947471,1.0659018,0.93315214,0.80430686,0.6754616,0.60908675,0.5466163,0.48024148,0.41386664,0.3513962,0.28892577,0.23035973,0.1717937,0.10932326,0.05075723,0.20693332,0.359205,0.5153811,0.6715572,0.8238289,1.6281357,2.436347,3.240654,4.044961,4.8492675,4.60329,4.3534083,4.1074314,3.8614538,3.611572,3.1313305,2.6471848,2.1630387,1.6827974,1.1986516,1.678893,2.1591344,2.639376,3.1196175,3.5998588,2.9439192,2.2918842,1.6359446,0.98000497,0.3240654,1.6867018,3.0454338,4.4041657,5.7668023,7.125534,8.015738,8.909846,9.803954,10.694158,11.588266,11.318862,11.0494585,10.77615,10.506746,10.237343,9.175345,8.113348,7.0513506,5.989353,4.9234514,5.55206,6.180669,6.8092775,7.433982,8.062591,8.281238,8.495979,8.714626,8.933272,9.148014,9.140205,9.128492,9.120684,9.108971,9.101162,13.130505,17.163752,21.197,25.230247,29.263494,25.882282,22.50107,19.123762,15.74255,12.361338,12.83377,13.302299,13.770826,14.243259,14.711788,15.039758,15.367727,15.695697,16.023666,16.351637,14.7156925,13.079747,11.443803,9.811763,8.175818,12.67369,17.175465,21.673336,26.175114,30.67689,34.2338,37.79071,41.34762,44.90453,48.46144,41.093834,33.72232,26.350811,18.983204,11.611692,14.008995,16.402393,18.795792,21.193096,23.586494,20.931501,18.276506,15.621513,12.96652,10.311526,9.155824,8.0040245,6.8483214,5.6926184,4.5369153,3.631094,2.7213683,1.815547,0.9058213,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10541886,0.15617609,0.21083772,0.26159495,0.24597734,0.23426414,0.21864653,0.20302892,0.18741131,0.6832704,1.1791295,1.6710842,2.1669433,2.6628022,3.0532427,3.4436827,3.8341231,4.220659,4.6110992,3.7638438,2.9165885,2.069333,1.2220778,0.37482262,1.038571,1.698415,2.3621633,3.0259118,3.6857557,3.5295796,3.3734035,3.213323,3.057147,2.900971,2.9048753,2.9087796,2.9165885,2.920493,2.9243972,2.338737,1.756981,1.1713207,0.58566034,0.0,0.0,0.0,0.0,0.0,0.0,0.21083772,0.42557985,0.63641757,0.8511597,1.0619974,1.3314011,1.6008049,1.8741131,2.1435168,2.4129205,2.6081407,2.8072653,3.0063896,3.2016098,3.4007344,2.7213683,2.0380979,1.358732,0.679366,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,1.3353056,2.6706111,4.0059166,5.3412223,6.676528,5.3412223,4.0059166,2.6706111,1.3353056,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.48414588,0.6637484,0.8472553,1.0307622,1.2142692,0.96829176,0.7262188,0.48414588,0.24207294,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.06637484,0.09761006,0.12884527,0.1639849,0.14055848,0.11713207,0.093705654,0.07418364,0.05075723,0.058566034,0.07027924,0.078088045,0.08980125,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.058566034,0.06637484,0.07418364,0.078088045,0.08589685,0.08589685,0.08199245,0.078088045,0.078088045,0.07418364,0.10151446,0.12494087,0.14836729,0.1756981,0.19912452,0.26159495,0.3240654,0.38653582,0.44900626,0.5114767,0.60908675,0.7066968,0.80430686,0.9019169,0.999527,0.95657855,0.9136301,0.8706817,0.8316377,0.78868926,0.8511597,0.91753453,0.98390937,1.0463798,1.1127546,1.1127546,1.1127546,1.1127546,1.1127546,1.1127546,0.9956226,0.8784905,0.76135844,0.6442264,0.5231899,0.44119745,0.3553006,0.26940376,0.1835069,0.10151446,0.14055848,0.1835069,0.22645533,0.26940376,0.31235218,0.77697605,1.2415999,1.7062237,2.1708477,2.639376,2.2723622,1.9092526,1.542239,1.1791295,0.81211567,0.7066968,0.59737355,0.48805028,0.38263142,0.27330816,0.49195468,0.7106012,0.92924774,1.1439898,1.3626363,1.9756275,2.592523,3.2094188,3.8224099,4.4393053,4.369026,4.3026514,4.2362766,4.165997,4.0996222,3.951255,3.7989833,3.6506162,3.4983444,3.349977,3.416352,3.4866312,3.5530062,3.619381,3.6857557,3.2367494,2.787743,2.338737,1.8858263,1.43682,1.2962615,1.1517987,1.0112402,0.8667773,0.7262188,0.6910792,0.659844,0.62860876,0.59346914,0.5622339,0.5544251,0.5466163,0.5388075,0.5309987,0.5231899,0.5466163,0.5661383,0.58566034,0.60518235,0.62470436,0.6676528,0.7106012,0.75354964,0.79649806,0.8355421,0.9058213,0.97219616,1.038571,1.1088502,1.175225,1.3509232,1.5266213,1.698415,1.8741131,2.0498111,2.6432803,3.2367494,3.8263142,4.4197836,5.0132523,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.44119745,0.7301232,1.0190489,1.3118792,1.6008049,2.1005683,2.6003318,3.1000953,3.5998588,4.0996222,4.6384296,5.181142,5.7199492,6.2587566,6.801469,7.223144,7.6448197,8.066495,8.488171,8.913751,8.781001,8.652155,8.52331,8.39056,8.261715,9.4018,10.537982,11.674163,12.814248,13.950429,14.090988,14.235451,14.376009,14.520472,14.661031,14.516567,14.3682,14.219833,14.0714655,13.923099,13.610746,13.29449,12.978233,12.665881,12.349625,13.450665,14.551707,15.648844,16.749886,17.850927,20.295082,22.739239,25.183395,27.631454,30.075611,29.700788,29.32987,28.958952,28.58413,28.213211,27.822771,27.432331,27.04189,26.65145,26.26101,23.274141,20.28337,17.292597,14.301826,11.311053,13.884054,16.457056,19.030056,21.603058,24.17606,27.643167,31.110277,34.577385,38.044495,41.511604,39.31733,37.12306,34.928783,32.730602,30.53633,29.431385,28.326439,27.221493,26.116547,25.0116,36.685764,48.36383,60.037994,71.71216,83.38632,67.881935,52.377556,36.873177,21.368793,5.860508,5.919074,5.9737353,6.028397,6.083059,6.13772,5.3997884,4.661856,3.9239242,3.1859922,2.4480603,4.6540475,6.8561306,9.058213,11.260296,13.462379,11.23687,9.01136,6.785851,4.564246,2.338737,3.0532427,3.767748,4.482254,5.196759,5.911265,4.8375545,3.7638438,2.6862288,1.6125181,0.5388075,1.456342,2.377781,3.2992198,4.2167544,5.138193,5.64967,6.1611466,6.676528,7.1880045,7.699481,9.030883,10.358379,11.68978,13.021181,14.348679,11.779582,9.2104845,6.6413884,4.068387,1.4992905,1.2025559,0.9058213,0.60908675,0.30844778,0.011713207,0.019522011,0.027330816,0.03513962,0.042948425,0.05075723,0.08589685,0.12494087,0.1639849,0.19912452,0.23816854,0.25378615,0.27330816,0.28892577,0.30844778,0.3240654,2.2918842,4.2557983,6.2197127,8.183627,10.151445,8.316377,6.4852123,4.6540475,2.8189783,0.9878138,1.2845483,1.5812829,1.8819219,2.1786566,2.475391,2.1630387,1.8506867,1.5383345,1.2259823,0.9136301,0.80821127,0.7066968,0.60518235,0.5036679,0.39824903,0.3670138,0.3357786,0.30063897,0.26940376,0.23816854,0.19522011,0.15227169,0.10932326,0.06637484,0.023426414,0.20302892,0.37872702,0.5583295,0.7340276,0.9136301,1.9287747,2.9439192,3.959064,4.9742084,5.989353,5.2084727,4.4275923,3.6467118,2.8658314,2.0888553,1.7882162,1.4914817,1.1947471,0.8980125,0.60127795,1.3040704,2.0068626,2.7057507,3.408543,4.1113358,3.3460727,2.5808098,1.815547,1.0541886,0.28892577,1.4797685,2.6706111,3.8653584,5.056201,6.250948,8.066495,9.878138,11.693685,13.509232,15.324779,13.802062,12.2793455,10.756628,9.2339115,7.7111945,6.676528,5.6379566,4.5993857,3.5608149,2.5261483,3.49444,4.466636,5.434928,6.4032197,7.375416,6.9654536,6.5554914,6.1455293,5.735567,5.3256044,5.2318993,5.138193,5.0483923,4.9546866,4.860981,8.410083,11.959184,15.504381,19.053482,22.59868,20.70895,18.81922,16.92949,15.039758,13.150026,13.110983,13.0719385,13.028991,12.989946,12.950902,13.157836,13.364769,13.571702,13.778636,13.985569,12.919667,11.8537655,10.783959,9.718058,8.648251,13.599033,18.549814,23.500597,28.45138,33.39826,38.25924,43.12022,47.9812,52.838276,57.699257,49.02758,40.355904,31.684225,23.008642,14.336966,14.711788,15.0827055,15.453624,15.828446,16.199366,14.871868,13.544372,12.216875,10.889378,9.561881,8.859089,8.156297,7.453504,6.7507114,6.0518236,4.841459,3.631094,2.4207294,1.2103647,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.113227665,0.1717937,0.23035973,0.28892577,0.25378615,0.22255093,0.19131571,0.15617609,0.12494087,0.48414588,0.8433509,1.2064602,1.5656652,1.9248703,2.7565079,3.5881457,4.423688,5.2553253,6.086963,4.9078336,3.7287042,2.5456703,1.3665408,0.18741131,0.8628729,1.5383345,2.2137961,2.8892577,3.5608149,3.4905357,3.416352,3.3460727,3.2718892,3.2016098,3.338264,3.4788225,3.619381,3.7599394,3.900498,3.1196175,2.338737,1.5617609,0.78088045,0.0,0.0,0.0,0.0,0.0,0.0,0.23816854,0.47633708,0.7106012,0.94876975,1.1869383,1.3235924,1.456342,1.5929961,1.7257458,1.8623998,1.9912452,2.1239948,2.25284,2.3816853,2.514435,2.0107672,1.5070993,1.0034313,0.5036679,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,1.7804074,3.5608149,5.3412223,7.1216297,8.898132,7.1216297,5.3412223,3.5608149,1.7804074,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.042948425,0.08589685,0.12884527,0.1717937,0.21083772,0.29673457,0.38263142,0.46852827,0.5544251,0.63641757,0.5114767,0.38263142,0.25378615,0.12884527,0.0,0.0,0.0,0.0,0.0,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.14446288,0.113227665,0.08589685,0.05466163,0.023426414,0.042948425,0.058566034,0.078088045,0.093705654,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.03513962,0.046852827,0.05466163,0.06637484,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.19912452,0.23816854,0.27330816,0.31235218,0.3513962,0.49195468,0.63641757,0.77697605,0.92143893,1.0619974,1.0463798,1.0307622,1.0190489,1.0034313,0.9878138,1.0580931,1.1283722,1.1986516,1.2689307,1.33921,1.33921,1.33921,1.33921,1.33921,1.33921,1.2103647,1.0815194,0.95657855,0.8277333,0.698888,0.58175594,0.46462387,0.3474918,0.23035973,0.113227665,0.14055848,0.1678893,0.19522011,0.22255093,0.24988174,0.7340276,1.2142692,1.698415,2.1786566,2.6628022,2.2684577,1.8741131,1.475864,1.0815194,0.6871748,0.60127795,0.5192855,0.43338865,0.3474918,0.26159495,0.47633708,0.6910792,0.9058213,1.1205635,1.33921,1.9209659,2.5027218,3.084478,3.6662338,4.251894,4.0722914,3.8965936,3.716991,3.541293,3.3616903,3.4983444,3.638903,3.775557,3.912211,4.0488653,4.165997,4.279225,4.396357,4.5095844,4.6267166,4.037152,3.4514916,2.8619268,2.2762666,1.6867018,1.4992905,1.3079748,1.116659,0.92924774,0.737932,0.7027924,0.6676528,0.63251317,0.59737355,0.5622339,0.5388075,0.5192855,0.4958591,0.47243267,0.44900626,0.46071947,0.46852827,0.48024148,0.48805028,0.4997635,0.5270943,0.5544251,0.58175594,0.60908675,0.63641757,0.7418364,0.8433509,0.94486535,1.0463798,1.1517987,1.2884527,1.4251068,1.5617609,1.698415,1.8389735,2.6042364,3.3694992,4.1308575,4.8961205,5.661383,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.5388075,0.8862993,1.2376955,1.5890918,1.9365835,2.475391,3.0141985,3.5491016,4.087909,4.6267166,4.786797,4.950782,5.1108627,5.2748475,5.4388323,6.0518236,6.66091,7.2739015,7.8868923,8.499884,8.1992445,7.898606,7.601871,7.3012323,7.000593,7.812709,8.624825,9.43694,10.249056,11.061172,11.287627,11.514082,11.736633,11.963089,12.185639,12.525322,12.861101,13.200784,13.536563,13.8762455,13.751305,13.626364,13.501423,13.376482,13.251541,13.774731,14.301826,14.825015,15.348206,15.875299,18.073479,20.27556,22.47374,24.675823,26.874,25.698776,24.52355,23.348326,22.1731,21.00178,20.338032,19.674282,19.010534,18.35069,17.686943,14.149553,10.612165,7.0747766,3.5373883,0.0,2.4988174,5.001539,7.5003567,9.999174,12.501896,17.023193,21.548395,26.073599,30.5988,35.124004,33.92535,32.7267,31.524143,30.325493,29.12684,27.276154,25.425468,23.574781,21.724094,19.873407,35.338745,50.80018,66.26161,81.72695,97.18838,78.09976,59.011135,39.922512,20.837795,1.7491722,1.7491722,1.7491722,1.7491722,1.7491722,1.7491722,1.999054,2.2489357,2.4988174,2.7486992,2.998581,2.4012074,1.7999294,1.1986516,0.60127795,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,1.5617609,2.9361105,4.3143644,5.688714,7.0630636,5.64967,4.2362766,2.8267872,1.4133936,0.0,1.2767396,2.5495746,3.8263142,5.099149,6.375889,7.012306,7.648724,8.289046,8.925464,9.561881,11.23687,12.911859,14.586847,16.261835,17.936825,14.723501,11.514082,8.300759,5.087436,1.8741131,1.4992905,1.1244678,0.74964523,0.37482262,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.10151446,0.13665408,0.1756981,0.21083772,0.24988174,0.23816854,0.22645533,0.21083772,0.19912452,0.18741131,2.5769055,4.9624953,7.3519893,9.737579,12.123169,9.737579,7.3519893,4.9624953,2.5769055,0.18741131,0.48805028,0.78868926,1.0893283,1.3860629,1.6867018,1.4485333,1.2142692,0.97610056,0.737932,0.4997635,0.42557985,0.3513962,0.27330816,0.19912452,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.19912452,0.39824903,0.60127795,0.80040246,0.999527,2.2255092,3.4514916,4.6735697,5.899552,7.125534,5.813655,4.5017757,3.1859922,1.8741131,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.92534333,1.8506867,2.77603,3.7013733,4.6267166,3.7482262,2.87364,1.999054,1.1244678,0.24988174,1.2767396,2.2996929,3.3265507,4.349504,5.376362,8.113348,10.850334,13.58732,16.324306,19.061293,16.289165,13.513136,10.737106,7.9610763,5.1889505,4.173806,3.1625657,2.1513257,1.1361811,0.12494087,1.43682,2.7486992,4.0644827,5.376362,6.688241,5.64967,4.6110992,3.5764325,2.5378613,1.4992905,1.3235924,1.1517987,0.97610056,0.80040246,0.62470436,3.6857557,6.7507114,9.811763,12.8767185,15.93777,15.535617,15.137367,14.739119,14.336966,13.938716,13.388195,12.837675,12.287154,11.736633,11.186112,11.275913,11.361811,11.4516115,11.537509,11.623405,11.123642,10.6238785,10.124115,9.6243515,9.124588,14.524376,19.924164,25.323954,30.723742,36.12353,42.28858,48.449726,54.610874,60.775925,66.93707,56.961323,46.989483,37.013733,27.037985,17.062239,15.410676,13.763018,12.111456,10.4637985,8.812236,8.812236,8.812236,8.812236,8.812236,8.812236,8.562354,8.312472,8.062591,7.812709,7.562827,6.0518236,4.5369153,3.0259118,1.5110037,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.28892577,0.5114767,0.737932,0.96438736,1.1869383,2.463678,3.736513,5.0132523,6.2860875,7.562827,6.0518236,4.5369153,3.0259118,1.5110037,0.0,0.6871748,1.3743496,2.0615244,2.7486992,3.435874,3.4514916,3.4632049,3.474918,3.4866312,3.4983444,3.775557,4.0488653,4.3260775,4.5993857,4.8765984,3.900498,2.9243972,1.9482968,0.97610056,0.0,0.0,0.0,0.0,0.0,0.0,0.26159495,0.5231899,0.78868926,1.0502841,1.3118792,1.3118792,1.3118792,1.3118792,1.3118792,1.3118792,1.3743496,1.43682,1.4992905,1.5617609,1.6242313,1.3001659,0.97610056,0.6481308,0.3240654,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,2.2255092,4.4510183,6.676528,8.898132,11.123642,8.898132,6.676528,4.4510183,2.2255092,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.37482262,0.5622339,0.74964523,0.93705654,1.1244678,1.1361811,1.1517987,1.1635119,1.175225,1.1869383,1.261122,1.33921,1.4133936,1.4875772,1.5617609,1.5617609,1.5617609,1.5617609,1.5617609,1.5617609,1.4251068,1.2884527,1.1517987,1.0112402,0.8745861,0.7262188,0.57394713,0.42557985,0.27330816,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.6871748,1.1869383,1.6867018,2.1864653,2.6862288,2.260649,1.8389735,1.4133936,0.9878138,0.5622339,0.4997635,0.43729305,0.37482262,0.31235218,0.24988174,0.46071947,0.6754616,0.8862993,1.1010414,1.3118792,1.8623998,2.4129205,2.9634414,3.513962,4.0605783,3.775557,3.4866312,3.2016098,2.912684,2.6237583,3.049338,3.474918,3.900498,4.3260775,4.7516575,4.911738,5.0757227,5.2358036,5.3997884,5.563773,4.8375545,4.1113358,3.3890212,2.6628022,1.9365835,1.698415,1.4641509,1.2259823,0.9878138,0.74964523,0.7106012,0.6754616,0.63641757,0.60127795,0.5622339,0.5231899,0.48805028,0.44900626,0.41386664,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.38653582,0.39824903,0.41386664,0.42557985,0.43729305,0.57394713,0.7106012,0.8511597,0.9878138,1.1244678,1.2259823,1.3235924,1.4251068,1.5266213,1.6242313,2.5612879,3.4983444,4.4393053,5.376362,6.3134184,0.19912452,0.1796025,0.16008049,0.14055848,0.12103647,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.47243267,0.75745404,1.0424755,1.3274968,1.6125181,2.0927596,2.5730011,3.0532427,3.533484,4.0137253,4.3065557,4.60329,4.8961205,5.192855,5.4856853,5.833177,6.1767645,6.524256,6.8678436,7.211431,7.172387,7.1333427,7.094299,7.0513506,7.012306,7.7658563,8.52331,9.276859,10.034314,10.787864,11.20173,11.615597,12.033368,12.447234,12.861101,13.192975,13.520945,13.852819,14.180789,14.512663,14.415053,14.317443,14.219833,14.122223,14.024612,14.871868,15.7152195,16.55857,17.405825,18.249176,20.228708,22.20824,24.191677,26.171207,28.15074,26.729538,25.308336,23.891037,22.469835,21.048632,19.971018,18.889498,17.811884,16.730364,15.648844,14.590752,13.536563,12.47847,11.420377,10.362284,11.256392,12.146595,13.040704,13.930907,14.825015,18.440493,22.059874,25.679255,29.29473,32.914112,31.079042,29.243973,27.408903,25.573835,23.738766,22.305851,20.876839,19.447828,18.018816,16.585901,29.017517,41.449135,53.876846,66.308464,78.736176,63.84869,48.961205,34.07372,19.186234,4.298747,3.7482262,3.2016098,2.6510892,2.1005683,1.5500476,1.8819219,2.2137961,2.5456703,2.8814487,3.213323,2.5730011,1.9326792,1.2923572,0.6520352,0.011713207,0.039044023,0.06637484,0.093705654,0.12103647,0.14836729,1.2650263,2.3816853,3.49444,4.6110992,5.7238536,4.743849,3.7638438,2.7838387,1.8038338,0.8238289,1.7062237,2.5886188,3.4710135,4.3534083,5.2358036,5.735567,6.239235,6.7389984,7.238762,7.7385254,9.136301,10.534078,11.931853,13.325725,14.723501,12.216875,9.710248,7.2036223,4.6930914,2.1864653,1.7882162,1.3938715,0.9956226,0.59737355,0.19912452,0.1756981,0.15617609,0.13274968,0.10932326,0.08589685,0.12103647,0.15617609,0.19131571,0.22645533,0.26159495,0.26940376,0.27721256,0.28502136,0.29283017,0.30063897,2.1903696,4.0801005,5.969831,7.859562,9.749292,8.289046,6.824895,5.3607445,3.900498,2.436347,2.2294137,2.018576,1.8077383,1.5969005,1.3860629,1.5890918,1.7882162,1.9873407,2.1864653,2.3855898,2.1318035,1.8780174,1.6242313,1.3665408,1.1127546,1.1986516,1.2806439,1.3665408,1.4524376,1.5383345,1.5227169,1.5070993,1.4914817,1.475864,1.4641509,1.7335546,2.0068626,2.280171,2.5534792,2.8267872,3.6467118,4.4705405,5.2943697,6.114294,6.9381227,5.6418614,4.3416953,3.0454338,1.7491722,0.44900626,0.5036679,0.5544251,0.60908675,0.659844,0.7106012,1.3118792,1.9092526,2.5066261,3.1039999,3.7013733,3.3343596,2.97125,2.6042364,2.241127,1.8741131,2.5769055,3.279698,3.9824903,4.6852827,5.388075,8.246098,11.10412,13.958238,16.816261,19.674282,16.570284,13.466284,10.358379,7.2543793,4.1503797,4.0020123,3.853645,3.7091823,3.5608149,3.4124475,3.9317331,4.4510183,4.9742084,5.493494,6.012779,5.2436123,4.474445,3.7013733,2.9322062,2.1630387,2.241127,2.3192148,2.3933985,2.4714866,2.5495746,4.9468775,7.3402762,9.733675,12.130978,14.524376,14.243259,13.966047,13.68493,13.403813,13.1266,12.486279,11.849861,11.213444,10.573121,9.936704,10.22563,10.518459,10.807385,11.096312,11.389141,10.936231,10.48332,10.03041,9.577498,9.124588,13.661504,18.194515,22.73143,27.26444,31.801357,39.906895,48.00853,56.11407,64.219604,72.32515,60.963337,49.60543,38.24362,26.885714,15.523903,14.711788,13.899672,13.087557,12.27544,11.4633255,12.173926,12.880623,13.591225,14.301826,15.012426,13.466284,11.916236,10.370092,8.823949,7.2739015,5.8214636,4.365122,2.9087796,1.456342,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.59346914,0.8902037,1.1869383,1.4797685,1.7765031,1.8858263,1.9951496,2.1044729,2.2137961,2.3231194,3.06886,3.814601,4.560342,5.3060827,6.0518236,5.8761253,5.704332,5.532538,5.3607445,5.1889505,4.93126,4.677474,4.423688,4.165997,3.912211,3.7052777,3.4983444,3.2914112,3.0805733,2.87364,3.6349986,4.396357,5.153811,5.9151692,6.676528,5.4895897,4.3065557,3.1196175,1.9365835,0.74964523,0.60127795,0.44900626,0.30063897,0.14836729,0.0,0.21083772,0.42167544,0.62860876,0.8394465,1.0502841,1.0541886,1.0580931,1.0659018,1.0698062,1.0737107,1.1439898,1.2142692,1.2845483,1.3548276,1.4251068,1.2103647,0.9956226,0.78088045,0.5661383,0.3513962,0.30844778,0.26940376,0.23035973,0.19131571,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,1.7804074,3.5608149,5.3412223,7.1216297,8.898132,7.3051367,5.708236,4.11524,2.5183394,0.92534333,0.8823949,0.8394465,0.79649806,0.75354964,0.7106012,0.5700427,0.42557985,0.28502136,0.14055848,0.0,0.0,0.0,0.0,0.0,0.0,0.48024148,0.96048295,1.4407244,1.9209659,2.4012074,2.2957885,2.194274,2.0927596,1.9912452,1.8858263,1.8858263,1.8819219,1.8819219,1.8780174,1.8741131,1.6515622,1.4290112,1.2064602,0.98390937,0.76135844,0.679366,0.59346914,0.5075723,0.42167544,0.3357786,0.26940376,0.20302892,0.13665408,0.06637484,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.10932326,0.12103647,0.12884527,0.14055848,0.14836729,0.3240654,0.4997635,0.6754616,0.8511597,1.0268579,1.0307622,1.0346665,1.038571,1.0463798,1.0502841,1.097137,1.1439898,1.1908426,1.2415999,1.2884527,1.2962615,1.3040704,1.3118792,1.3157835,1.3235924,1.2689307,1.2103647,1.1517987,1.0932326,1.038571,0.8667773,0.698888,0.5270943,0.359205,0.18741131,0.19131571,0.19131571,0.19522011,0.19912452,0.19912452,0.6676528,1.1361811,1.6008049,2.069333,2.5378613,2.135708,1.737459,1.33921,0.93705654,0.5388075,0.48414588,0.43338865,0.37872702,0.3279698,0.27330816,0.45681506,0.64032197,0.8238289,1.0034313,1.1869383,1.6749885,2.1630387,2.6510892,3.1391394,3.6232853,3.3655949,3.1039999,2.8463092,2.5847144,2.3231194,2.6510892,2.979059,3.3070288,3.6349986,3.9629683,4.087909,4.21285,4.337791,4.462732,4.5876727,4.029343,3.4671092,2.9087796,2.3465457,1.7882162,1.6008049,1.4133936,1.2259823,1.038571,0.8511597,0.8160201,0.78088045,0.74574083,0.7106012,0.6754616,0.6481308,0.62470436,0.60127795,0.57394713,0.5505207,0.58175594,0.61689556,0.6481308,0.679366,0.7106012,0.7262188,0.7418364,0.75745404,0.77307165,0.78868926,0.8511597,0.91753453,0.98390937,1.0463798,1.1127546,1.1947471,1.2767396,1.358732,1.4407244,1.5266213,2.338737,3.154757,3.970777,4.786797,5.5989127,0.14836729,0.16008049,0.1717937,0.1796025,0.19131571,0.19912452,0.1796025,0.16008049,0.14055848,0.12103647,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.40605783,0.62860876,0.8472553,1.0659018,1.2884527,1.7101282,2.1318035,2.5534792,2.979059,3.4007344,3.8263142,4.2557983,4.6813784,5.1108627,5.5364423,5.6145306,5.6926184,5.7707067,5.8487945,5.9268827,6.1455293,6.364176,6.5867267,6.805373,7.0240197,7.7229075,8.421796,9.116779,9.815667,10.510651,11.115833,11.721016,12.326198,12.93138,13.536563,13.860628,14.180789,14.504854,14.828919,15.14908,15.078801,15.008522,14.938243,14.871868,14.801589,15.965101,17.128613,18.296028,19.459541,20.626957,22.383938,24.144823,25.905708,27.666594,29.423576,27.7603,26.09312,24.429846,22.76657,21.09939,19.604004,18.104713,16.609327,15.110037,13.610746,15.035853,16.457056,17.878258,19.303364,20.724567,20.010061,19.295555,18.58105,17.866545,17.148134,19.861694,22.57135,25.281004,27.99066,30.700315,28.228828,25.761246,23.289759,20.818274,18.35069,17.33945,16.32821,15.320874,14.309634,13.298394,22.696291,32.094185,41.492085,50.88998,60.287876,49.601524,38.911274,28.224924,17.538574,6.8483214,5.7511845,4.650143,3.5491016,2.4480603,1.3509232,1.7647898,2.1786566,2.5964274,3.0102942,3.4241607,2.7447948,2.0654287,1.3860629,0.7066968,0.023426414,0.042948425,0.058566034,0.078088045,0.093705654,0.113227665,0.96829176,1.8233559,2.67842,3.533484,4.388548,3.8419318,3.2914112,2.7447948,2.1981785,1.6515622,2.1396124,2.631567,3.1196175,3.611572,4.0996222,4.462732,4.825841,5.1889505,5.548156,5.911265,7.0318284,8.152391,9.272955,10.393518,11.514082,9.710248,7.9064145,6.1064854,4.3026514,2.4988174,2.0810463,1.6593709,1.2415999,0.8199245,0.39824903,0.3435874,0.28502136,0.22645533,0.1717937,0.113227665,0.14446288,0.1756981,0.21083772,0.24207294,0.27330816,0.30063897,0.3318742,0.359205,0.38653582,0.41386664,1.8038338,3.1977055,4.591577,5.9815445,7.375416,6.8366084,6.3017054,5.7628975,5.22409,4.689187,3.9668727,3.2484627,2.5261483,1.8077383,1.0893283,1.7257458,2.3621633,2.998581,3.638903,4.2753205,3.8419318,3.4046388,2.97125,2.533957,2.1005683,2.2684577,2.4402514,2.6081407,2.7799344,2.951728,2.9439192,2.9400148,2.9361105,2.9283018,2.9243972,3.2718892,3.6154766,3.959064,4.3065557,4.650143,5.0718184,5.4895897,5.911265,6.329036,6.7507114,5.466163,4.185519,2.900971,1.620327,0.3357786,0.5544251,0.77307165,0.9917182,1.2064602,1.4251068,1.6945106,1.9639144,2.233318,2.5066261,2.77603,2.920493,3.0649557,3.2094188,3.3538816,3.4983444,3.8809757,4.2597027,4.6384296,5.0210614,5.3997884,8.378847,11.354002,14.33306,17.308216,20.287273,16.8514,13.419431,9.983557,6.547683,3.1118085,3.8302186,4.548629,5.263134,5.9815445,6.699954,6.426646,6.153338,5.883934,5.610626,5.337318,4.83365,4.3338866,3.8302186,3.3265507,2.8267872,3.154757,3.4866312,3.814601,4.1464753,4.474445,6.2040954,7.929841,9.659492,11.385237,13.110983,12.950902,12.790822,12.630741,12.470661,12.31058,11.588266,10.862047,10.135828,9.413514,8.687295,9.17925,9.671205,10.163159,10.6590185,11.150972,10.744915,10.338858,9.936704,9.530646,9.124588,12.794726,16.464865,20.135002,23.805141,27.475279,37.521305,47.571236,57.617264,67.66329,77.71323,64.96535,52.22138,39.47741,26.733442,13.985569,14.012899,14.036326,14.063657,14.087084,14.114414,15.531713,16.952915,18.374117,19.791414,21.212618,18.366308,15.523903,12.677594,9.8312845,6.98888,5.591104,4.193328,2.795552,1.397776,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.113227665,0.1717937,0.23035973,0.28892577,0.92924774,1.5656652,2.2059872,2.8463092,3.4866312,3.4827268,3.4788225,3.4710135,3.4671092,3.4632049,3.677947,3.892689,4.1074314,4.322173,4.5369153,5.704332,6.871748,8.039165,9.20658,10.373997,9.17925,7.9805984,6.7819467,5.5832953,4.388548,3.959064,3.533484,3.1039999,2.67842,2.2489357,3.49444,4.7399445,5.985449,7.230953,8.476458,7.0786815,5.6848097,4.290938,2.893162,1.4992905,1.1986516,0.9019169,0.60127795,0.30063897,0.0,0.15617609,0.31625658,0.47243267,0.62860876,0.78868926,0.79649806,0.80821127,0.8160201,0.8277333,0.8394465,0.9136301,0.9917182,1.0698062,1.1478943,1.2259823,1.1205635,1.0151446,0.9097257,0.80430686,0.698888,0.59346914,0.49195468,0.38653582,0.28111696,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,1.3353056,2.6706111,4.0059166,5.3412223,6.676528,5.708236,4.743849,3.7794614,2.815074,1.8506867,1.7413634,1.6281357,1.5188124,1.4094892,1.3001659,1.038571,0.78088045,0.5192855,0.26159495,0.0,0.0,0.0,0.0,0.0,0.0,0.93315214,1.8702087,2.803361,3.7404175,4.6735697,4.493967,4.3143644,4.134762,3.9551594,3.775557,3.7443218,3.7130866,3.6857557,3.6545205,3.6232853,3.193801,2.7604125,2.3270237,1.893635,1.4641509,1.3040704,1.1478943,0.9917182,0.8316377,0.6754616,0.5388075,0.40605783,0.26940376,0.13665408,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.08199245,0.08980125,0.09761006,0.10541886,0.113227665,0.27330816,0.43729305,0.60127795,0.76135844,0.92534333,0.92143893,0.92143893,0.91753453,0.9136301,0.9136301,0.93315214,0.95267415,0.97219616,0.9917182,1.0112402,1.0268579,1.0424755,1.0580931,1.0737107,1.0893283,1.1088502,1.1322767,1.1557031,1.1791295,1.1986516,1.0112402,0.8199245,0.62860876,0.44119745,0.24988174,0.24207294,0.23426414,0.22645533,0.21864653,0.21083772,0.6481308,1.0815194,1.5188124,1.9522011,2.3855898,2.0107672,1.6359446,1.261122,0.8862993,0.5114767,0.46852827,0.42557985,0.38653582,0.3435874,0.30063897,0.45291066,0.60518235,0.75745404,0.9097257,1.0619974,1.4875772,1.9131571,2.338737,2.7643168,3.1859922,2.9556324,2.7213683,2.4910088,2.2567444,2.0263848,2.2567444,2.4831998,2.7135596,2.9439192,3.174279,3.2640803,3.349977,3.435874,3.5256753,3.611572,3.2172275,2.822883,2.4285383,2.0341935,1.6359446,1.4992905,1.3626363,1.2259823,1.0893283,0.94876975,0.91753453,0.8862993,0.8511597,0.8199245,0.78868926,0.77307165,0.76135844,0.74964523,0.737932,0.7262188,0.78868926,0.8550641,0.92143893,0.98390937,1.0502841,1.0659018,1.0854238,1.1010414,1.1205635,1.1361811,1.1283722,1.1205635,1.116659,1.1088502,1.1010414,1.1635119,1.2298868,1.2962615,1.358732,1.4251068,2.1161861,2.8111696,3.5022488,4.193328,4.8883114,0.10151446,0.14055848,0.1796025,0.21864653,0.26159495,0.30063897,0.26940376,0.23816854,0.21083772,0.1796025,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.3435874,0.4958591,0.6520352,0.80821127,0.96438736,1.3274968,1.6906061,2.05762,2.4207294,2.787743,3.3460727,3.9083066,4.466636,5.02887,5.5871997,5.395884,5.2084727,5.017157,4.825841,4.6384296,5.1186714,5.5989127,6.0791545,6.559396,7.0357327,7.676055,8.316377,8.956698,9.597021,10.237343,11.033841,11.826434,12.622932,13.419431,14.212025,14.528281,14.840633,15.15689,15.473146,15.789403,15.746454,15.7035055,15.660558,15.617609,15.57466,17.058334,18.54591,20.029583,21.513256,23.000834,24.539167,26.081408,27.619741,29.16198,30.700315,28.791061,26.88181,24.968653,23.0594,21.150146,19.233086,17.31993,15.406772,13.48971,11.576552,15.477051,19.381453,23.28195,27.186354,31.086851,28.763731,26.444517,24.121397,21.798277,19.475159,21.278992,23.078922,24.882755,26.68659,28.486519,25.382519,22.278519,19.170614,16.066616,12.962616,12.373051,11.783486,11.193921,10.600452,10.010887,16.378967,22.743143,29.107319,35.471493,41.83567,35.350456,28.861341,22.37613,15.8870125,9.4018,7.7502384,6.098676,4.4510183,2.7994564,1.1517987,1.6476578,2.1435168,2.6432803,3.1391394,3.638903,2.9165885,2.1981785,1.475864,0.75745404,0.039044023,0.046852827,0.05075723,0.058566034,0.06637484,0.07418364,0.6715572,1.2650263,1.8584955,2.455869,3.049338,2.9361105,2.8189783,2.7057507,2.5886188,2.475391,2.5730011,2.6706111,2.7682211,2.8658314,2.9634414,3.1859922,3.4124475,3.638903,3.8614538,4.087909,4.93126,5.7707067,6.6140575,7.4574084,8.300759,7.2036223,6.1064854,5.009348,3.9083066,2.8111696,2.3699722,1.9287747,1.4836729,1.0424755,0.60127795,0.5075723,0.41386664,0.3240654,0.23035973,0.13665408,0.1678893,0.19912452,0.22645533,0.25769055,0.28892577,0.3357786,0.38263142,0.42948425,0.47633708,0.5231899,1.4212024,2.3153105,3.2094188,4.1035266,5.001539,5.388075,5.774611,6.1611466,6.551587,6.9381227,5.708236,4.478349,3.2484627,2.018576,0.78868926,1.8623998,2.9361105,4.0137253,5.087436,6.1611466,5.548156,4.93126,4.318269,3.7013733,3.0883822,3.3421683,3.5959544,3.853645,4.1074314,4.3612175,4.369026,4.3729305,4.376835,4.380739,4.388548,4.806319,5.22409,5.6418614,6.055728,6.473499,6.493021,6.5086384,6.5281606,6.5437784,6.5633,5.2943697,4.029343,2.7604125,1.4914817,0.22645533,0.60908675,0.9917182,1.3743496,1.7530766,2.135708,2.0810463,2.0224805,1.9639144,1.9092526,1.8506867,2.5066261,3.1586614,3.814601,4.4705405,5.12648,5.181142,5.239708,5.298274,5.35684,5.4115014,8.511597,11.607788,14.703979,17.804073,20.900265,17.136421,13.368673,9.60483,5.840986,2.0732377,3.6584249,5.239708,6.8209906,8.406178,9.987461,8.921559,7.8556576,6.79366,5.727758,4.661856,4.4275923,4.193328,3.959064,3.7208953,3.4866312,4.068387,4.6540475,5.2358036,5.8175592,6.3993154,7.461313,8.519405,9.581403,10.639496,11.701493,11.6585455,11.619501,11.580457,11.541413,11.498465,10.686349,9.874233,9.062118,8.250002,7.437886,8.13287,8.827853,9.522837,10.217821,10.912805,10.553599,10.198298,9.839094,9.483793,9.124588,11.931853,14.735214,17.538574,20.34584,23.1492,35.13962,47.13004,59.12046,71.11088,83.101295,68.96736,54.841232,40.7112,26.581171,12.4511385,13.314012,14.176885,15.035853,15.8987255,16.761599,18.893402,21.021301,23.153105,25.281004,27.412807,23.270237,19.127666,14.985096,10.8425255,6.699954,5.3607445,4.0215344,2.67842,1.33921,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05466163,0.10932326,0.1639849,0.21864653,0.27330816,1.261122,2.2450314,3.2289407,4.2167544,5.2006636,5.0796275,4.958591,4.841459,4.7204223,4.5993857,4.283129,3.970777,3.6545205,3.338264,3.0259118,5.532538,8.039165,10.545791,13.056321,15.562947,13.423335,11.283723,9.14411,7.000593,4.860981,4.2167544,3.5686235,2.920493,2.2723622,1.6242313,3.3538816,5.083532,6.813182,8.546737,10.276386,8.671678,7.066968,5.4583545,3.853645,2.2489357,1.7999294,1.3509232,0.9019169,0.44900626,0.0,0.10541886,0.21083772,0.31625658,0.42167544,0.5231899,0.5388075,0.5544251,0.5700427,0.58566034,0.60127795,0.6832704,0.76916724,0.8550641,0.94096094,1.0268579,1.0307622,1.0346665,1.038571,1.0463798,1.0502841,0.8784905,0.7106012,0.5388075,0.3709182,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.8902037,1.7804074,2.6706111,3.5608149,4.4510183,4.11524,3.7794614,3.4436827,3.1118085,2.77603,2.5964274,2.4207294,2.241127,2.0654287,1.8858263,1.5110037,1.1322767,0.75354964,0.37872702,0.0,0.0,0.0,0.0,0.0,0.0,1.3899672,2.7799344,4.169902,5.559869,6.949836,6.6921453,6.434455,6.1767645,5.919074,5.661383,5.606722,5.548156,5.4895897,5.4310236,5.376362,4.732136,4.0918136,3.4475873,2.803361,2.1630387,1.9326792,1.7023194,1.4719596,1.2415999,1.0112402,0.80821127,0.60908675,0.40605783,0.20302892,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05466163,0.058566034,0.06637484,0.07027924,0.07418364,0.22645533,0.37482262,0.5231899,0.6754616,0.8238289,0.8160201,0.80430686,0.79649806,0.78478485,0.77307165,0.76916724,0.76135844,0.75354964,0.74574083,0.737932,0.76135844,0.78088045,0.80430686,0.8277333,0.8511597,0.95267415,1.0541886,1.1557031,1.261122,1.3626363,1.1517987,0.94096094,0.7340276,0.5231899,0.31235218,0.29673457,0.27721256,0.26159495,0.24207294,0.22645533,0.62860876,1.0307622,1.4329157,1.8350691,2.2372224,1.8858263,1.5383345,1.1869383,0.8394465,0.48805028,0.45681506,0.42167544,0.39044023,0.359205,0.3240654,0.44900626,0.5700427,0.6910792,0.8160201,0.93705654,1.3001659,1.6632754,2.0263848,2.3855898,2.7486992,2.5456703,2.338737,2.135708,1.9287747,1.7257458,1.8584955,1.9912452,2.1239948,2.2567444,2.3855898,2.436347,2.4871042,2.5378613,2.5886188,2.639376,2.4090161,2.1786566,1.9482968,1.717937,1.4875772,1.4016805,1.3118792,1.2259823,1.1361811,1.0502841,1.0190489,0.9917182,0.96048295,0.92924774,0.9019169,0.9019169,0.9019169,0.9019169,0.9019169,0.9019169,0.9956226,1.0932326,1.1908426,1.2884527,1.3860629,1.4055848,1.4290112,1.4485333,1.4680552,1.4875772,1.4055848,1.3274968,1.2494087,1.1674163,1.0893283,1.1361811,1.183034,1.2298868,1.2767396,1.3235924,1.893635,2.463678,3.0337205,3.6037633,4.173806,0.05075723,0.12103647,0.19131571,0.26159495,0.3318742,0.39824903,0.359205,0.32016098,0.28111696,0.23816854,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.27721256,0.3670138,0.45681506,0.5466163,0.63641757,0.94486535,1.2533131,1.5617609,1.8663043,2.174752,2.8658314,3.5608149,4.251894,4.9468775,5.6379566,5.181142,4.7243266,4.263607,3.8067923,3.349977,4.0918136,4.829746,5.571582,6.309514,7.0513506,7.633106,8.214863,8.796618,9.378374,9.964035,10.947944,11.931853,12.915763,13.903577,14.8874855,15.195933,15.504381,15.808925,16.117373,16.42582,16.410202,16.394585,16.378967,16.36335,16.351637,18.15547,19.959305,21.763138,23.570877,25.37471,26.694399,28.014086,29.333775,30.653461,31.97315,29.821825,27.666594,25.511364,23.356134,21.200905,18.866072,16.535143,14.204215,11.869383,9.538455,15.918248,22.301945,28.685644,35.06934,41.449135,37.521305,33.589573,29.661743,25.730011,21.798277,22.696291,23.590399,24.484507,25.378614,26.276627,22.53621,18.795792,15.055375,11.314958,7.57454,7.406651,7.2348576,7.0630636,6.8951745,6.7233806,10.05774,13.388195,16.722555,20.053009,23.38737,21.09939,18.81141,16.52343,14.239355,11.951375,9.749292,7.551114,5.349031,3.1508527,0.94876975,1.5305257,2.1083772,2.690133,3.2718892,3.8497405,3.0883822,2.330928,1.5695697,0.80821127,0.05075723,0.046852827,0.046852827,0.042948425,0.039044023,0.039044023,0.3709182,0.7066968,1.0424755,1.3782539,1.7140326,2.0302892,2.3465457,2.6667068,2.9829633,3.2992198,3.0063896,2.7096553,2.416825,2.1200905,1.8233559,1.9131571,1.999054,2.0888553,2.174752,2.260649,2.8267872,3.3929255,3.959064,4.521298,5.087436,4.6930914,4.3026514,3.9083066,3.5178664,3.1235218,2.6588979,2.194274,1.7296503,1.2650263,0.80040246,0.6715572,0.5466163,0.41777104,0.28892577,0.1639849,0.19131571,0.21864653,0.24597734,0.27330816,0.30063897,0.3670138,0.43338865,0.5036679,0.5700427,0.63641757,1.0346665,1.4329157,1.8311646,2.2294137,2.6237583,3.9356375,5.251421,6.5633,7.8751793,9.187058,7.445695,5.708236,3.9668727,2.2294137,0.48805028,1.999054,3.513962,5.024966,6.5359693,8.050878,7.2543793,6.461786,5.6652875,4.8687897,4.0761957,4.415879,4.755562,5.095245,5.434928,5.774611,5.7902284,5.805846,5.8214636,5.833177,5.8487945,6.3407493,6.8287997,7.320754,7.8088045,8.300759,7.914223,7.531592,7.1450562,6.75852,6.375889,5.1225758,3.8692627,2.6159496,1.3665408,0.113227665,0.659844,1.2064602,1.7530766,2.3035975,2.8502135,2.463678,2.0810463,1.6945106,1.3118792,0.92534333,2.0888553,3.2562714,4.4197836,5.5832953,6.7507114,6.4852123,6.2197127,5.9542136,5.688714,5.423215,8.644346,11.861574,15.078801,18.296028,21.513256,17.417538,13.32182,9.226103,5.134289,1.038571,3.4866312,5.930787,8.378847,10.826907,13.274967,11.416472,9.561881,7.703386,5.84489,3.9863946,4.0215344,4.0527697,4.084005,4.1191444,4.1503797,4.985922,5.8214636,6.6531014,7.4886436,8.324185,8.718531,9.108971,9.503315,9.893755,10.2881,10.366188,10.44818,10.526268,10.608261,10.686349,9.788337,8.886419,7.988407,7.08649,6.1884775,7.08649,7.9805984,8.878611,9.776623,10.674636,10.366188,10.053836,9.745388,9.43694,9.124588,11.065076,13.005564,14.946052,16.88654,18.823124,32.757935,46.688843,60.623653,74.55456,88.48937,72.97328,57.457184,41.94109,26.4289,10.912805,12.611219,14.313539,16.011953,17.714273,19.412687,22.251188,25.093594,27.932095,30.774498,33.613,28.174168,22.73143,17.292597,11.8537655,6.4110284,5.1303844,3.8458362,2.5651922,1.2806439,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10541886,0.15617609,0.21083772,0.26159495,1.5929961,2.9243972,4.251894,5.5832953,6.910792,6.676528,6.4422636,6.2079997,5.9737353,5.735567,4.892216,4.0488653,3.2016098,2.358259,1.5110037,5.3607445,9.20658,13.056321,16.902157,20.751898,17.66742,14.586847,11.502369,8.421796,5.337318,4.4705405,3.6037633,2.7330816,1.8663043,0.999527,3.213323,5.4310236,7.6448197,9.858616,12.076316,10.260769,8.445222,6.629675,4.814128,2.998581,2.4012074,1.7999294,1.1986516,0.60127795,0.0,0.05075723,0.10541886,0.15617609,0.21083772,0.26159495,0.28111696,0.30063897,0.3240654,0.3435874,0.3631094,0.45681506,0.5466163,0.64032197,0.7340276,0.8238289,0.94096094,1.0541886,1.1713207,1.2845483,1.4016805,1.1635119,0.92924774,0.6949836,0.46071947,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.44510186,0.8902037,1.3353056,1.7804074,2.2255092,2.5183394,2.815074,3.1118085,3.4046388,3.7013733,3.455396,3.2094188,2.9634414,2.7213683,2.475391,1.979532,1.4836729,0.9917182,0.4958591,0.0,0.0,0.0,0.0,0.0,0.0,1.8467822,3.68966,5.5364423,7.37932,9.226103,8.890324,8.554545,8.218767,7.8868923,7.551114,7.465217,7.37932,7.2934237,7.211431,7.125534,6.2743745,5.4193106,4.5681505,3.7130866,2.8619268,2.5612879,2.2567444,1.9561055,1.6515622,1.3509232,1.0815194,0.80821127,0.5388075,0.26940376,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.027330816,0.031235218,0.031235218,0.03513962,0.039044023,0.1756981,0.31235218,0.44900626,0.58566034,0.7262188,0.7066968,0.6910792,0.6715572,0.6559396,0.63641757,0.60127795,0.5661383,0.5309987,0.4958591,0.46071947,0.49195468,0.5231899,0.5544251,0.58175594,0.61299115,0.79649806,0.97610056,1.1596074,1.3431144,1.5266213,1.2962615,1.0659018,0.8355421,0.60518235,0.37482262,0.3474918,0.32016098,0.29283017,0.26549935,0.23816854,0.60908675,0.97610056,1.3470187,1.717937,2.0888553,1.7608855,1.43682,1.1127546,0.78868926,0.46071947,0.44119745,0.41777104,0.39434463,0.3709182,0.3513962,0.44119745,0.5349031,0.62860876,0.71841,0.81211567,1.1127546,1.4133936,1.7140326,2.0107672,2.3114061,2.135708,1.9561055,1.7804074,1.6008049,1.4251068,1.4602464,1.4953861,1.5305257,1.5656652,1.6008049,1.6125181,1.6242313,1.6359446,1.6515622,1.6632754,1.5969005,1.53443,1.4680552,1.4016805,1.33921,1.3001659,1.261122,1.2259823,1.1869383,1.1517987,1.1205635,1.0932326,1.0659018,1.038571,1.0112402,1.0268579,1.038571,1.0502841,1.0619974,1.0737107,1.2064602,1.3353056,1.4641509,1.5969005,1.7257458,1.7491722,1.7686942,1.7921207,1.815547,1.8389735,1.6867018,1.53443,1.3782539,1.2259823,1.0737107,1.1049459,1.1361811,1.1635119,1.1947471,1.2259823,1.6710842,2.1200905,2.5690966,3.0141985,3.4632049,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.44900626,0.39824903,0.3513962,0.30063897,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.21083772,0.23816854,0.26159495,0.28892577,0.31235218,0.5622339,0.81211567,1.0619974,1.3118792,1.5617609,2.3855898,3.213323,4.037152,4.860981,5.688714,4.9624953,4.2362766,3.513962,2.787743,2.0615244,3.0610514,4.0605783,5.0640097,6.0635366,7.0630636,7.5862536,8.113348,8.636538,9.163632,9.686822,10.862047,12.037272,13.212498,14.387722,15.562947,15.863586,16.164225,16.46096,16.761599,17.062239,17.073952,17.085665,17.101282,17.112995,17.124708,19.248703,21.376602,23.500597,25.624592,27.748587,28.849628,29.95067,31.051712,32.14885,33.24989,30.848682,28.45138,26.05017,23.648964,21.251661,18.499058,15.750359,13.001659,10.249056,7.5003567,16.36335,25.226343,34.089336,42.948425,51.811417,46.274975,40.738533,35.198185,29.661743,24.125301,24.113588,24.101875,24.086258,24.074545,24.062832,19.685997,15.313066,10.936231,6.5633,2.1864653,2.436347,2.6862288,2.9361105,3.1859922,3.435874,3.736513,4.037152,4.337791,4.6384296,4.939069,6.8483214,8.761478,10.674636,12.587793,14.50095,11.748346,8.999647,6.250948,3.4983444,0.74964523,1.4133936,2.0732377,2.736986,3.4007344,4.0605783,3.2640803,2.463678,1.6632754,0.8628729,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,1.1244678,1.8741131,2.6237583,3.3734035,4.123049,3.435874,2.7486992,2.0615244,1.3743496,0.6871748,0.63641757,0.58566034,0.5388075,0.48805028,0.43729305,0.7262188,1.0112402,1.3001659,1.5890918,1.8741131,2.1864653,2.4988174,2.8111696,3.1235218,3.435874,2.951728,2.463678,1.9756275,1.4875772,0.999527,0.8394465,0.6754616,0.5114767,0.3513962,0.18741131,0.21083772,0.23816854,0.26159495,0.28892577,0.31235218,0.39824903,0.48805028,0.57394713,0.6637484,0.74964523,0.6481308,0.5505207,0.44900626,0.3513962,0.24988174,2.4871042,4.7243266,6.9615493,9.198771,11.435994,9.187058,6.9381227,4.689187,2.436347,0.18741131,2.135708,4.087909,6.036206,7.988407,9.936704,8.960603,7.988407,7.012306,6.036206,5.0640097,5.4856853,5.911265,6.336845,6.7624245,7.1880045,7.211431,7.238762,7.262188,7.2856145,7.3129454,7.8751793,8.437413,8.999647,9.561881,10.124115,9.339331,8.550641,7.7619514,6.9732623,6.1884775,4.950782,3.7130866,2.475391,1.2376955,0.0,0.7106012,1.4251068,2.135708,2.8502135,3.5608149,2.8502135,2.135708,1.4251068,0.7106012,0.0,1.6749885,3.349977,5.024966,6.699954,8.374943,7.7892823,7.1997175,6.6140575,6.0244927,5.4388323,8.773191,12.111456,15.449719,18.787983,22.126247,17.698656,13.274967,8.85128,4.423688,0.0,3.310933,6.6257706,9.936704,13.251541,16.562475,13.911386,11.2642,8.6131115,5.9620223,3.310933,3.611572,3.912211,4.21285,4.513489,4.814128,5.899552,6.98888,8.074304,9.163632,10.249056,9.975748,9.698535,9.425227,9.151918,8.874706,9.073831,9.276859,9.475985,9.675109,9.874233,8.886419,7.898606,6.910792,5.9268827,4.939069,6.036206,7.137247,8.238289,9.339331,10.436467,10.174872,9.913278,9.651682,9.386183,9.124588,10.198298,11.275913,12.349625,13.423335,14.50095,30.37625,46.247646,62.12685,78.00215,93.87354,76.97529,60.077038,43.17488,26.276627,9.37447,11.912332,14.450192,16.988054,19.525915,22.063778,25.612879,29.16198,32.711082,36.264088,39.81319,33.074192,26.339098,19.6001,12.861101,6.126007,4.900025,3.6740425,2.4480603,1.2259823,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,1.9248703,3.5998588,5.2748475,6.949836,8.624825,8.273428,7.9259367,7.57454,7.223144,6.8756523,5.5013027,4.126953,2.7486992,1.3743496,0.0,5.1889505,10.373997,15.562947,20.751898,25.936945,21.911505,17.886066,13.860628,9.839094,5.813655,4.7243266,3.638903,2.5495746,1.4641509,0.37482262,3.076669,5.774611,8.476458,11.174399,13.8762455,11.849861,9.823476,7.800996,5.774611,3.7482262,2.998581,2.2489357,1.4992905,0.74964523,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.22645533,0.3240654,0.42557985,0.5231899,0.62470436,0.8511597,1.0737107,1.3001659,1.5266213,1.7491722,1.4485333,1.1517987,0.8511597,0.5505207,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.92534333,1.8506867,2.77603,3.7013733,4.6267166,4.3143644,3.998108,3.6857557,3.3734035,3.0610514,2.4480603,1.8389735,1.2259823,0.61299115,0.0,0.0,0.0,0.0,0.0,0.0,2.2996929,4.5993857,6.899079,9.198771,11.498465,11.088503,10.674636,10.260769,9.850807,9.43694,9.323712,9.21439,9.101162,8.987934,8.874706,7.812709,6.7507114,5.688714,4.6267166,3.5608149,3.1859922,2.8111696,2.436347,2.0615244,1.6867018,1.3509232,1.0112402,0.6754616,0.3357786,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,0.60127795,0.57394713,0.5505207,0.5231899,0.4997635,0.43729305,0.37482262,0.31235218,0.24988174,0.18741131,0.22645533,0.26159495,0.30063897,0.3357786,0.37482262,0.63641757,0.9019169,1.1635119,1.4251068,1.6867018,1.43682,1.1869383,0.93705654,0.6871748,0.43729305,0.39824903,0.3631094,0.3240654,0.28892577,0.24988174,0.58566034,0.92534333,1.261122,1.6008049,1.9365835,1.6359446,1.33921,1.038571,0.737932,0.43729305,0.42557985,0.41386664,0.39824903,0.38653582,0.37482262,0.43729305,0.4997635,0.5622339,0.62470436,0.6871748,0.92534333,1.1635119,1.4016805,1.6359446,1.8741131,1.7257458,1.5734742,1.4251068,1.2767396,1.1244678,1.0619974,0.999527,0.93705654,0.8745861,0.81211567,0.78868926,0.76135844,0.737932,0.7106012,0.6871748,0.78868926,0.8862993,0.9878138,1.0893283,1.1869383,1.1986516,1.2142692,1.2259823,1.2376955,1.2494087,1.2259823,1.1986516,1.175225,1.1517987,1.1244678,1.1517987,1.175225,1.1986516,1.2259823,1.2494087,1.4133936,1.5734742,1.737459,1.901444,2.0615244,2.0888553,2.1122816,2.135708,2.1630387,2.1864653,1.9639144,1.737459,1.5110037,1.2884527,1.0619974,1.0737107,1.0893283,1.1010414,1.1127546,1.1244678,1.4485333,1.7765031,2.1005683,2.4246337,2.7486992,1.6359446,1.4133936,1.1869383,0.96438736,0.737932,0.5114767,0.5192855,0.5231899,0.5270943,0.5309987,0.5388075,0.42948425,0.3240654,0.21474212,0.10932326,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.19131571,0.23035973,0.26940376,0.30844778,0.3513962,0.5309987,0.7106012,0.8902037,1.0698062,1.2494087,1.9404879,2.631567,3.3187418,4.009821,4.7009,4.5369153,4.376835,4.21285,4.0488653,3.8887846,4.3846436,4.884407,5.380266,5.8761253,6.375889,6.801469,7.223144,7.648724,8.074304,8.499884,9.999174,11.49456,12.993851,14.489237,15.988527,16.613232,17.237936,17.86264,18.487345,19.11205,19.194042,19.27213,19.354122,19.43221,19.514202,21.532778,23.551353,25.573835,27.592411,29.610987,29.575848,29.540707,29.509472,29.474333,29.439194,27.811058,26.182922,24.554787,22.926651,21.298513,19.533724,17.76503,15.996336,14.231546,12.4628525,18.272602,24.082354,29.892103,35.701855,41.511604,37.068394,32.62909,28.18588,23.74267,19.29946,19.43221,19.56496,19.69771,19.83046,19.96321,17.058334,14.157363,11.256392,8.351517,5.4505453,5.376362,5.3060827,5.2318993,5.1616197,5.087436,4.93126,4.7711797,4.6150036,4.4588275,4.298747,5.8487945,7.394938,8.941081,10.491129,12.037272,9.858616,7.676055,5.4973984,3.3187418,1.1361811,1.8663043,2.592523,3.3187418,4.0488653,4.775084,3.951255,3.1313305,2.3075018,1.4836729,0.6637484,0.8511597,1.0424755,1.2337911,1.4212024,1.6125181,1.5851873,1.5578566,1.5305257,1.5031948,1.475864,2.077142,2.67842,3.2836022,3.8848803,4.4861584,3.8770714,3.2679846,2.6588979,2.0459068,1.43682,1.2884527,1.1439898,0.9956226,0.8472553,0.698888,1.0659018,1.4290112,1.796025,2.1591344,2.5261483,2.5769055,2.6237583,2.6745155,2.7252727,2.77603,2.3933985,2.0146716,1.6359446,1.2533131,0.8745861,0.80040246,0.7262188,0.6481308,0.57394713,0.4997635,0.44900626,0.39824903,0.3513962,0.30063897,0.24988174,0.32016098,0.39044023,0.46071947,0.5309987,0.60127795,0.8316377,1.0659018,1.2962615,1.5305257,1.7608855,3.240654,4.716518,6.196286,7.6721506,9.151918,7.3519893,5.548156,3.7482262,1.9482968,0.14836729,1.7140326,3.279698,4.845363,6.4110284,7.9766936,7.1997175,6.426646,5.64967,4.8765984,4.0996222,4.4510183,4.7985106,5.1499066,5.5013027,5.8487945,5.852699,5.8566036,5.8566036,5.860508,5.8644123,6.3134184,6.7624245,7.211431,7.6643414,8.113348,7.660437,7.2075267,6.754616,6.3017054,5.8487945,4.9624953,4.0761957,3.1859922,2.2996929,1.4133936,1.698415,1.9873407,2.2762666,2.5612879,2.8502135,2.2918842,1.7335546,1.1791295,0.62079996,0.062470436,1.5890918,3.1157131,4.646239,6.17286,7.699481,7.6721506,7.6448197,7.617489,7.590158,7.562827,9.698535,11.834243,13.966047,16.101755,18.237463,14.707883,11.178304,7.648724,4.1191444,0.58566034,3.1196175,5.6535745,8.183627,10.717585,13.251541,11.412568,9.573594,7.7385254,5.899552,4.0605783,4.0761957,4.087909,4.0996222,4.1113358,4.126953,5.6262436,7.125534,8.624825,10.124115,11.623405,11.174399,10.721489,10.268578,9.815667,9.362757,9.846903,10.327144,10.81129,11.291532,11.775677,10.221725,8.663869,7.1099167,5.5559645,3.998108,5.1186714,6.2353306,7.3519893,8.468649,9.589212,9.163632,8.738052,8.312472,7.8868923,7.461313,8.308568,9.155824,10.006983,10.8542385,11.701493,24.882755,38.060112,51.241375,64.41873,77.6,64.77794,51.95588,39.133823,26.307863,13.4858055,15.7035055,17.921206,20.138906,22.356607,24.574308,27.080935,29.583656,32.090282,34.59691,37.09963,32.144943,27.190258,22.23557,17.280884,12.326198,10.155351,7.988407,5.8214636,3.6545205,1.4875772,1.2259823,0.96829176,0.7066968,0.44900626,0.18741131,0.1678893,0.14836729,0.12884527,0.10932326,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.21083772,1.6945106,3.174279,4.6540475,6.133816,7.6135845,7.445695,7.28171,7.1177254,6.9537406,6.785851,6.309514,5.833177,5.35684,4.8765984,4.4002614,8.749765,13.09927,17.448774,21.798277,26.151686,22.516687,18.88169,15.246691,11.611692,7.9766936,8.218767,8.464745,8.710721,8.956698,9.198771,10.865952,12.533132,14.204215,15.871395,17.538574,14.903104,12.271536,9.639969,7.008402,4.376835,3.4983444,2.6237583,1.7491722,0.8745861,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.22645533,0.3513962,0.47633708,0.60127795,0.7262188,1.0346665,1.3431144,1.6554666,1.9639144,2.2762666,2.2177005,2.1591344,2.1005683,2.0459068,1.9873407,1.5890918,1.1908426,0.79649806,0.39824903,0.0,0.05466163,0.10932326,0.1639849,0.21864653,0.27330816,0.96048295,1.6437533,2.330928,3.0141985,3.7013733,3.4514916,3.2016098,2.951728,2.7018464,2.4480603,1.9600099,1.4719596,0.98000497,0.48805028,0.0,0.13665408,0.27330816,0.41386664,0.5505207,0.6871748,2.5456703,4.40807,6.266566,8.128965,9.987461,10.377901,10.768341,11.158782,11.549222,11.935758,10.990892,10.046027,9.101162,8.156297,7.211431,7.016211,6.817086,6.621866,6.422742,6.223617,5.251421,4.2753205,3.2992198,2.3231194,1.3509232,1.0815194,0.80821127,0.5388075,0.26940376,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.5622339,0.62470436,0.6871748,0.74964523,0.81211567,0.7145056,0.61689556,0.5192855,0.42167544,0.3240654,0.3357786,0.3435874,0.3553006,0.3631094,0.37482262,0.58175594,0.78478485,0.9917182,1.1947471,1.4016805,1.2064602,1.0112402,0.8160201,0.62079996,0.42557985,0.38653582,0.3513962,0.31235218,0.27330816,0.23816854,0.5388075,0.8355421,1.1361811,1.43682,1.737459,1.4680552,1.1986516,0.92924774,0.6559396,0.38653582,0.37482262,0.3631094,0.3513962,0.3357786,0.3240654,0.39044023,0.45681506,0.5192855,0.58566034,0.6481308,0.8433509,1.038571,1.2337911,1.4290112,1.6242313,1.5383345,1.456342,1.3704453,1.2845483,1.1986516,1.1205635,1.0463798,0.96829176,0.8902037,0.81211567,0.78088045,0.74574083,0.7145056,0.6832704,0.6481308,0.7262188,0.80040246,0.8745861,0.94876975,1.0268579,1.0502841,1.0737107,1.1010414,1.1244678,1.1517987,1.1400855,1.1283722,1.1205635,1.1088502,1.1010414,1.1088502,1.116659,1.1205635,1.1283722,1.1361811,1.2689307,1.4016805,1.53443,1.6671798,1.7999294,1.8506867,1.901444,1.9482968,1.999054,2.0498111,1.8545911,1.6593709,1.4641509,1.2689307,1.0737107,1.1127546,1.1517987,1.1869383,1.2259823,1.261122,1.5578566,1.8506867,2.1474214,2.4441557,2.736986,3.2757936,2.7252727,2.174752,1.6242313,1.0737107,0.5231899,0.58566034,0.6442264,0.7066968,0.76526284,0.8238289,0.659844,0.4958591,0.3318742,0.1639849,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.1678893,0.22255093,0.27721256,0.3318742,0.38653582,0.4958591,0.60908675,0.71841,0.8277333,0.93705654,1.4914817,2.0459068,2.6042364,3.1586614,3.7130866,4.1113358,4.513489,4.911738,5.3138914,5.7121406,5.708236,5.704332,5.6965227,5.6926184,5.688714,6.012779,6.336845,6.66091,6.98888,7.3129454,9.132397,10.951848,12.771299,14.590752,16.414106,17.362877,18.311647,19.26432,20.21309,21.16186,21.310228,21.458595,21.606962,21.751425,21.899792,23.816854,25.730011,27.643167,29.56023,31.473387,30.305971,29.13465,27.96333,26.795912,25.624592,24.769527,23.914463,23.0594,22.204336,21.349272,20.564487,19.779701,18.994917,18.210133,17.425346,20.181856,22.938364,25.698776,28.455284,31.211792,27.865719,24.515741,21.169668,17.823597,14.473619,14.750832,15.028045,15.309161,15.586374,15.863586,14.430671,13.001659,11.572648,10.143637,8.710721,8.316377,7.9220324,7.5276875,7.1333427,6.7389984,6.1221027,5.5091114,4.892216,4.279225,3.6623292,4.845363,6.028397,7.211431,8.39056,9.573594,7.9649806,6.356367,4.743849,3.135235,1.5266213,2.3192148,3.1118085,3.9044023,4.6930914,5.4856853,4.6423345,3.7989833,2.951728,2.1083772,1.261122,1.6554666,2.0459068,2.4402514,2.8306916,3.2250361,3.096191,2.9634414,2.8345962,2.7057507,2.5769055,3.0298162,3.4866312,3.9395418,4.396357,4.8492675,4.318269,3.7833657,3.252367,2.7213683,2.1864653,1.9443923,1.698415,1.4524376,1.2064602,0.96438736,1.4055848,1.8467822,2.2918842,2.7330816,3.174279,2.9634414,2.7486992,2.5378613,2.3231194,2.1122816,1.8389735,1.5656652,1.2962615,1.0229534,0.74964523,0.76135844,0.77307165,0.78868926,0.80040246,0.81211567,0.6871748,0.5622339,0.43729305,0.31235218,0.18741131,0.23816854,0.29283017,0.3435874,0.39824903,0.44900626,1.0151446,1.5812829,2.1435168,2.7096553,3.2757936,3.9942036,4.7087092,5.4271193,6.1455293,6.8639393,5.5130157,4.1620927,2.8111696,1.4641509,0.113227665,1.2923572,2.4714866,3.6506162,4.83365,6.012779,5.4388323,4.860981,4.2870336,3.7130866,3.1391394,3.4124475,3.6857557,3.9629683,4.2362766,4.513489,4.493967,4.4705405,4.4510183,4.4314966,4.4119744,4.7516575,5.087436,5.423215,5.7628975,6.098676,5.9815445,5.8644123,5.74728,5.630148,5.5130157,4.9742084,4.4393053,3.900498,3.3616903,2.8267872,2.6862288,2.5495746,2.4129205,2.2762666,2.135708,1.7335546,1.3314011,0.92924774,0.5270943,0.12494087,1.5031948,2.8853533,4.263607,5.645766,7.0240197,7.558923,8.089922,8.62092,9.155824,9.686822,10.619974,11.553126,12.486279,13.419431,14.348679,11.713207,9.081639,6.446168,3.8106966,1.175225,2.9283018,4.6813784,6.434455,8.183627,9.936704,8.913751,7.8868923,6.8639393,5.8370814,4.814128,4.5369153,4.263607,3.9863946,3.7130866,3.435874,5.349031,7.262188,9.175345,11.088503,13.001659,12.369146,11.740538,11.111929,10.479416,9.850807,10.61607,11.381332,12.146595,12.911859,13.673217,11.553126,9.4291315,7.309041,5.185046,3.0610514,4.1972322,5.3334136,6.46569,7.601871,8.738052,8.148487,7.562827,6.9732623,6.387602,5.7980375,6.4188375,7.039637,7.660437,8.281238,8.898132,19.385357,29.868677,40.355904,50.839222,61.326447,52.580585,43.834724,35.088863,26.343002,17.601046,19.498585,21.396124,23.293663,25.191204,27.088743,28.548988,30.009235,31.469482,32.925823,34.38607,31.215696,28.041416,24.871042,21.696764,18.526388,15.41458,12.306676,9.194867,6.083059,2.9751544,2.455869,1.9365835,1.4133936,0.8941081,0.37482262,0.3357786,0.29673457,0.25378615,0.21474212,0.1756981,0.1756981,0.1756981,0.1756981,0.1756981,0.1756981,1.4602464,2.7447948,4.029343,5.3138914,6.5984397,6.621866,6.6413884,6.66091,6.6804323,6.699954,7.1216297,7.5394006,7.9610763,8.378847,8.800523,12.314485,15.824542,19.338505,22.848562,26.362524,23.117966,19.873407,16.628849,13.384291,10.135828,11.713207,13.2905855,14.871868,16.449247,18.026625,18.659138,19.295555,19.931974,20.564487,21.200905,17.96025,14.719597,11.478943,8.238289,5.001539,3.998108,2.998581,1.999054,0.999527,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.22645533,0.37482262,0.5231899,0.6754616,0.8238289,1.2181735,1.6164225,2.0107672,2.4051118,2.7994564,2.9868677,3.1703746,3.3538816,3.541293,3.7247996,2.979059,2.233318,1.4914817,0.74574083,0.0,0.10932326,0.21864653,0.3318742,0.44119745,0.5505207,0.9956226,1.4407244,1.8858263,2.330928,2.77603,2.5886188,2.4012074,2.2137961,2.0263848,1.8389735,1.4680552,1.1010414,0.7340276,0.3670138,0.0,0.27330816,0.5505207,0.8238289,1.1010414,1.3743496,2.795552,4.2167544,5.6340523,7.055255,8.476458,9.6673,10.858143,12.05289,13.243732,14.438479,12.658072,10.881569,9.105066,7.328563,5.548156,6.2158084,6.883461,7.551114,8.218767,8.886419,7.3129454,5.7394714,4.1620927,2.5886188,1.0112402,0.80821127,0.60908675,0.40605783,0.20302892,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.5231899,0.6754616,0.8238289,0.97610056,1.1244678,0.9917182,0.8589685,0.7262188,0.59346914,0.46071947,0.44510186,0.42557985,0.40996224,0.39434463,0.37482262,0.5231899,0.6715572,0.8160201,0.96438736,1.1127546,0.97219616,0.8316377,0.6910792,0.5544251,0.41386664,0.37482262,0.3357786,0.30063897,0.26159495,0.22645533,0.48805028,0.74964523,1.0112402,1.2767396,1.5383345,1.2962615,1.0580931,0.8160201,0.57785153,0.3357786,0.3240654,0.31235218,0.30063897,0.28892577,0.27330816,0.3435874,0.40996224,0.47633708,0.5466163,0.61299115,0.76526284,0.91753453,1.0698062,1.2220778,1.3743496,1.3548276,1.3353056,1.3157835,1.2962615,1.2767396,1.183034,1.0893283,0.9956226,0.9058213,0.81211567,0.77307165,0.7340276,0.6910792,0.6520352,0.61299115,0.6637484,0.7106012,0.76135844,0.81211567,0.8628729,0.9019169,0.93705654,0.97610056,1.0112402,1.0502841,1.0541886,1.0580931,1.0659018,1.0698062,1.0737107,1.0659018,1.0541886,1.0463798,1.0346665,1.0268579,1.1283722,1.2298868,1.3314011,1.43682,1.5383345,1.6125181,1.6867018,1.7608855,1.8389735,1.9131571,1.7491722,1.5812829,1.4172981,1.2533131,1.0893283,1.1517987,1.2142692,1.2767396,1.33921,1.4016805,1.6632754,1.9287747,2.194274,2.4597735,2.7252727,4.911738,4.037152,3.1625657,2.2879796,1.4133936,0.5388075,0.6520352,0.76916724,0.8823949,0.9956226,1.1127546,0.8902037,0.6676528,0.44510186,0.22255093,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.14446288,0.21474212,0.28502136,0.3553006,0.42557985,0.46462387,0.5036679,0.5466163,0.58566034,0.62470436,1.0463798,1.4641509,1.8858263,2.3035975,2.7252727,3.6857557,4.650143,5.610626,6.575013,7.5394006,7.0318284,6.524256,6.016684,5.5091114,5.001539,5.22409,5.4505453,5.6730967,5.899552,6.126007,8.265619,10.409137,12.552653,14.69617,16.835783,18.112522,19.389261,20.662096,21.938837,23.211672,23.426414,23.641155,23.855898,24.07064,24.289286,26.097025,27.908667,29.716406,31.528048,33.335785,31.032188,28.728592,26.42109,24.117493,21.813896,21.727999,21.646006,21.564014,21.482021,21.400028,21.599154,21.794373,21.993498,22.188719,22.387842,22.091108,21.798277,21.501543,21.208714,20.911978,18.659138,16.406298,14.153459,11.900618,9.651682,10.073358,10.495033,10.916709,11.338385,11.763964,11.803008,11.845957,11.888905,11.931853,11.974802,11.256392,10.541886,9.823476,9.105066,8.386656,7.3168497,6.2431393,5.169429,4.095718,3.0259118,3.8419318,4.661856,5.477876,6.2938967,7.113821,6.0713453,5.0327744,3.9942036,2.951728,1.9131571,2.7682211,3.6271896,4.4861584,5.3412223,6.2001905,5.3334136,4.466636,3.5959544,2.7291772,1.8623998,2.455869,3.0532427,3.6467118,4.2440853,4.8375545,4.60329,4.3729305,4.138666,3.9083066,3.6740425,3.9824903,4.290938,4.5993857,4.903929,5.212377,4.759466,4.3026514,3.8458362,3.3929255,2.9361105,2.5964274,2.25284,1.9092526,1.5656652,1.2259823,1.7452679,2.2645533,2.7838387,3.3031244,3.8263142,3.349977,2.87364,2.4012074,1.9248703,1.4485333,1.2845483,1.1205635,0.95657855,0.78868926,0.62470436,0.7262188,0.8238289,0.92534333,1.0268579,1.1244678,0.92534333,0.7262188,0.5231899,0.3240654,0.12494087,0.16008049,0.19522011,0.23035973,0.26549935,0.30063897,1.1986516,2.096664,2.9907722,3.8887846,4.786797,4.743849,4.7009,4.661856,4.618908,4.575959,3.6740425,2.77603,1.8741131,0.97610056,0.07418364,0.8706817,1.6632754,2.4597735,3.2562714,4.0488653,3.6740425,3.2992198,2.9243972,2.5495746,2.174752,2.3738766,2.5769055,2.77603,2.9751544,3.174279,3.1313305,3.0883822,3.049338,3.0063896,2.9634414,3.1859922,3.4124475,3.638903,3.8614538,4.087909,4.3065557,4.521298,4.7399445,4.958591,5.173333,4.985922,4.7985106,4.6110992,4.423688,4.2362766,3.6740425,3.1118085,2.5495746,1.9873407,1.4251068,1.1791295,0.92924774,0.6832704,0.43338865,0.18741131,1.4212024,2.6510892,3.8848803,5.1186714,6.348558,7.4417906,8.535024,9.628256,10.721489,11.810817,11.541413,11.272009,11.002605,10.733202,10.4637985,8.722435,6.9810715,5.2436123,3.5022488,1.7608855,2.7330816,3.7091823,4.6813784,5.6535745,6.6257706,6.4110284,6.2001905,5.989353,5.774611,5.563773,5.001539,4.4393053,3.873167,3.310933,2.7486992,5.0757227,7.3988423,9.725866,12.0489855,14.376009,13.567798,12.759586,11.951375,11.143164,10.338858,11.385237,12.431617,13.481901,14.528281,15.57466,12.884527,10.194394,7.504261,4.814128,2.1239948,3.2757936,4.4314966,5.5832953,6.735094,7.8868923,7.137247,6.387602,5.6379566,4.8883114,4.138666,4.5291066,4.9234514,5.3138914,5.708236,6.098676,13.891863,21.681147,29.470428,37.259712,45.048992,40.383232,35.713566,31.047806,26.378141,21.712381,23.289759,24.867138,26.444517,28.021894,29.599274,30.01314,30.430912,30.844778,31.258644,31.676416,30.286448,28.89648,27.506514,26.116547,24.72658,20.67381,16.62104,12.568271,8.515501,4.462732,3.6818514,2.900971,2.1239948,1.3431144,0.5622339,0.5036679,0.44119745,0.38263142,0.3240654,0.26159495,0.23816854,0.21083772,0.18741131,0.1639849,0.13665408,1.2259823,2.3192148,3.408543,4.4978714,5.5871997,5.794133,5.997162,6.2040954,6.407124,6.6140575,7.929841,9.245625,10.565312,11.881096,13.200784,15.875299,18.549814,21.22433,23.898846,26.573362,23.719244,20.865126,18.011007,15.15689,12.298867,15.211552,18.12033,21.02911,23.941795,26.850574,26.452326,26.054077,25.655827,25.261482,24.863234,21.013493,17.167656,13.32182,9.47208,5.6262436,4.5017757,3.3734035,2.2489357,1.1244678,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.22645533,0.39824903,0.57394713,0.74964523,0.92534333,1.4055848,1.8858263,2.366068,2.8463092,3.3265507,3.7521305,4.181615,4.607195,5.036679,5.462259,4.369026,3.2757936,2.1864653,1.0932326,0.0,0.1639849,0.3318742,0.4958591,0.659844,0.8238289,1.0307622,1.2337911,1.4407244,1.6437533,1.8506867,1.7257458,1.6008049,1.475864,1.3509232,1.2259823,0.98000497,0.7340276,0.48805028,0.24597734,0.0,0.41386664,0.8238289,1.2376955,1.6515622,2.0615244,3.0415294,4.0215344,5.001539,5.9815445,6.9615493,8.956698,10.951848,12.946998,14.942147,16.937298,14.329156,11.717112,9.108971,6.4969254,3.8887846,5.4193106,6.9537406,8.484266,10.018696,11.549222,9.37447,7.1997175,5.024966,2.8502135,0.6754616,0.5388075,0.40605783,0.26940376,0.13665408,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.48805028,0.7262188,0.96438736,1.1986516,1.43682,1.2689307,1.1010414,0.93315214,0.76916724,0.60127795,0.5544251,0.5114767,0.46462387,0.42167544,0.37482262,0.46462387,0.5544251,0.6442264,0.7340276,0.8238289,0.7418364,0.6559396,0.5700427,0.48414588,0.39824903,0.3631094,0.3240654,0.28892577,0.24988174,0.21083772,0.43729305,0.6637484,0.8862993,1.1127546,1.33921,1.1283722,0.91753453,0.7066968,0.4958591,0.28892577,0.27330816,0.26159495,0.24988174,0.23816854,0.22645533,0.29673457,0.3631094,0.43338865,0.5036679,0.57394713,0.6832704,0.79649806,0.9058213,1.0151446,1.1244678,1.1713207,1.2142692,1.261122,1.3040704,1.3509232,1.2415999,1.1361811,1.0268579,0.92143893,0.81211567,0.76526284,0.71841,0.6715572,0.62079996,0.57394713,0.60127795,0.62470436,0.6481308,0.6754616,0.698888,0.74964523,0.80040246,0.8511597,0.9019169,0.94876975,0.96829176,0.9917182,1.0112402,1.0307622,1.0502841,1.0229534,0.9956226,0.96829176,0.94096094,0.9136301,0.98390937,1.0580931,1.1283722,1.2025559,1.2767396,1.3743496,1.475864,1.5734742,1.6749885,1.7765031,1.639849,1.5031948,1.3704453,1.2337911,1.1010414,1.1869383,1.2767396,1.3626363,1.4485333,1.5383345,1.7725986,2.0068626,2.241127,2.4792955,2.7135596,6.551587,5.349031,4.1503797,2.951728,1.7491722,0.5505207,0.71841,0.8902037,1.0580931,1.2298868,1.4016805,1.1205635,0.8394465,0.5583295,0.28111696,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.12103647,0.20693332,0.29283017,0.37872702,0.46071947,0.43338865,0.40215343,0.3709182,0.3435874,0.31235218,0.59737355,0.8823949,1.1674163,1.4524376,1.737459,3.2640803,4.786797,6.3134184,7.8361354,9.362757,8.351517,7.3441806,6.3329406,5.3217,4.3143644,4.4393053,4.564246,4.689187,4.814128,4.939069,7.4027467,9.866425,12.334006,14.797685,17.261362,18.862167,20.462973,22.063778,23.660677,25.261482,25.546503,25.827621,26.108738,26.393759,26.674877,28.3811,30.08342,31.789642,33.49587,35.198185,31.758408,28.31863,24.87885,21.439074,17.999294,18.690374,19.381453,20.068628,20.759706,21.450787,22.629915,23.809046,24.988174,26.171207,27.350338,24.004265,20.654287,17.308216,13.958238,10.612165,9.456462,8.296855,7.141152,5.9815445,4.825841,5.3919797,5.958118,6.5281606,7.094299,7.6643414,9.17925,10.694158,12.209065,13.723974,15.238882,14.196406,13.157836,12.119265,11.076789,10.0382185,8.507692,6.9771667,5.446641,3.9161155,2.3855898,2.8385005,3.2914112,3.7443218,4.1972322,4.650143,4.181615,3.7091823,3.240654,2.7682211,2.2996929,3.2211318,4.1464753,5.067914,5.989353,6.910792,6.0205884,5.134289,4.2440853,3.3538816,2.463678,3.260176,4.056674,4.853172,5.6535745,6.4500723,6.114294,5.7785153,5.446641,5.1108627,4.775084,4.9351645,5.095245,5.2553253,5.4154058,5.575486,5.196759,4.8219366,4.4432096,4.0644827,3.6857557,3.2484627,2.8072653,2.366068,1.9287747,1.4875772,2.084951,2.6823244,3.279698,3.8770714,4.474445,3.736513,2.998581,2.260649,1.5266213,0.78868926,0.7301232,0.6715572,0.61689556,0.5583295,0.4997635,0.6871748,0.8745861,1.0619974,1.2494087,1.43682,1.1635119,0.8862993,0.61299115,0.3357786,0.062470436,0.078088045,0.09761006,0.113227665,0.13274968,0.14836729,1.3782539,2.6081407,3.8419318,5.0718184,6.3017054,5.4973984,4.6930914,3.892689,3.0883822,2.2879796,1.8389735,1.3860629,0.93705654,0.48805028,0.039044023,0.44900626,0.8589685,1.2689307,1.678893,2.0888553,1.9131571,1.737459,1.5617609,1.3860629,1.2142692,1.33921,1.4641509,1.5890918,1.7140326,1.8389735,1.7725986,1.7062237,1.6437533,1.5773785,1.5110037,1.6242313,1.737459,1.8506867,1.9639144,2.0732377,2.6276627,3.1781836,3.7326086,4.283129,4.8375545,5.001539,5.1616197,5.3256044,5.4856853,5.64967,4.661856,3.6740425,2.6862288,1.698415,0.7106012,0.62079996,0.5270943,0.43338865,0.3435874,0.24988174,1.3353056,2.4207294,3.506153,4.591577,5.6730967,7.328563,8.980125,10.631687,12.28325,13.938716,12.466757,10.990892,9.518932,8.046973,6.575013,5.7316628,4.884407,4.041056,3.193801,2.35045,2.541766,2.7330816,2.9283018,3.1196175,3.310933,3.912211,4.513489,5.1108627,5.7121406,6.3134184,5.462259,4.6110992,3.7638438,2.912684,2.0615244,4.7985106,7.535496,10.276386,13.013372,15.750359,14.766449,13.778636,12.794726,11.810817,10.826907,12.154405,13.4858055,14.813302,16.144703,17.476105,14.215929,10.959657,7.703386,4.4432096,1.1869383,2.358259,3.5256753,4.6969957,5.8683167,7.0357327,6.126007,5.212377,4.298747,3.3890212,2.475391,2.639376,2.803361,2.97125,3.135235,3.2992198,8.3944645,13.48971,18.584955,23.6802,28.775444,28.18588,27.596315,27.00675,26.41328,25.823717,27.080935,28.338152,29.599274,30.856491,32.11371,31.481195,30.852587,30.223978,29.591465,28.962856,29.353296,29.74764,30.141985,30.532425,30.926771,25.929136,20.935406,15.941674,10.944039,5.950309,4.911738,3.8692627,2.8306916,1.7882162,0.74964523,0.6715572,0.58956474,0.5114767,0.42948425,0.3513962,0.30063897,0.24988174,0.19912452,0.14836729,0.10151446,0.9956226,1.8897307,2.7838387,3.6818514,4.575959,4.9663997,5.35684,5.743376,6.133816,6.524256,8.741957,10.955752,13.169549,15.383345,17.601046,19.436115,21.275087,23.114061,24.949131,26.788103,24.320522,21.856844,19.393166,16.925583,14.461906,18.705992,22.946173,27.190258,31.434343,35.674522,34.245514,32.8165,31.383585,29.954575,28.525562,24.07064,19.615717,15.160794,10.705871,6.250948,5.001539,3.7482262,2.4988174,1.2494087,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.22645533,0.42557985,0.62470436,0.8238289,1.0268579,1.5890918,2.15523,2.7213683,3.2836022,3.8497405,4.521298,5.1889505,5.860508,6.5281606,7.1997175,5.758993,4.318269,2.8814487,1.4407244,0.0,0.21864653,0.44119745,0.659844,0.8784905,1.1010414,1.0659018,1.0307622,0.9956226,0.96048295,0.92534333,0.8628729,0.80040246,0.737932,0.6754616,0.61299115,0.48805028,0.3670138,0.24597734,0.12103647,0.0,0.5505207,1.1010414,1.6515622,2.1981785,2.7486992,3.2914112,3.8302186,4.369026,4.911738,5.4505453,8.246098,11.045554,13.841106,16.640562,19.436115,15.996336,12.552653,9.108971,5.6691923,2.2255092,4.6228123,7.0201154,9.4174185,11.814721,14.212025,11.435994,8.663869,5.8878384,3.1118085,0.3357786,0.26940376,0.20302892,0.13665408,0.06637484,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.44900626,0.77307165,1.1010414,1.4251068,1.7491722,1.5461433,1.3431144,1.1439898,0.94096094,0.737932,0.6637484,0.59346914,0.5192855,0.44900626,0.37482262,0.40605783,0.44119745,0.47243267,0.5036679,0.5388075,0.5075723,0.47633708,0.44900626,0.41777104,0.38653582,0.3513962,0.31235218,0.27330816,0.23816854,0.19912452,0.38653582,0.57394713,0.76135844,0.94876975,1.1361811,0.95657855,0.77697605,0.59737355,0.41777104,0.23816854,0.22645533,0.21083772,0.19912452,0.18741131,0.1756981,0.24597734,0.32016098,0.39434463,0.46462387,0.5388075,0.60518235,0.6715572,0.7418364,0.80821127,0.8745861,0.98390937,1.0932326,1.2064602,1.3157835,1.4251068,1.3040704,1.1791295,1.0580931,0.93315214,0.81211567,0.75745404,0.7027924,0.6481308,0.59346914,0.5388075,0.5388075,0.5388075,0.5388075,0.5388075,0.5388075,0.60127795,0.6637484,0.7262188,0.78868926,0.8511597,0.8862993,0.92143893,0.95657855,0.9917182,1.0268579,0.98000497,0.93315214,0.8902037,0.8433509,0.80040246,0.8433509,0.8862993,0.92924774,0.96829176,1.0112402,1.1361811,1.261122,1.3860629,1.5110037,1.6359446,1.53443,1.4290112,1.3235924,1.2181735,1.1127546,1.2259823,1.33921,1.4485333,1.5617609,1.6749885,1.8819219,2.084951,2.2918842,2.494913,2.7018464,8.187531,6.66091,5.138193,3.611572,2.0888553,0.5622339,0.78868926,1.0112402,1.2376955,1.4641509,1.6867018,1.3509232,1.0112402,0.6754616,0.3357786,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.14836729,0.30063897,0.44900626,0.60127795,0.74964523,2.8385005,4.9234514,7.012306,9.101162,11.186112,9.675109,8.164105,6.649197,5.138193,3.6232853,3.6506162,3.6740425,3.7013733,3.7247996,3.7482262,6.5359693,9.323712,12.111456,14.899199,17.686943,19.611813,21.536682,23.461554,25.386423,27.311295,27.66269,28.014086,28.361578,28.712975,29.064371,30.66127,32.262077,33.86288,35.463684,37.060585,32.488533,27.91257,23.336613,18.760653,14.188598,15.648844,17.112995,18.573242,20.037392,21.501543,23.660677,25.823717,27.986755,30.149794,32.31283,25.913517,19.514202,13.110983,6.7116675,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.7106012,1.4251068,2.135708,2.8502135,3.5608149,6.551587,9.538455,12.525322,15.51219,18.499058,17.136421,15.773785,14.411149,13.048512,11.685876,9.698535,7.7111945,5.7238536,3.736513,1.7491722,1.8389735,1.9248703,2.0107672,2.1005683,2.1864653,2.2879796,2.3855898,2.4871042,2.5886188,2.6862288,3.6740425,4.661856,5.64967,6.6374836,7.6252975,6.7116675,5.801942,4.8883114,3.9746814,3.0610514,4.0605783,5.0640097,6.0635366,7.0630636,8.062591,7.6252975,7.1880045,6.7507114,6.3134184,5.8761253,5.8878384,5.899552,5.911265,5.9268827,5.938596,5.6379566,5.337318,5.036679,4.73604,4.4393053,3.900498,3.3616903,2.8267872,2.2879796,1.7491722,2.4246337,3.1000953,3.775557,4.4510183,5.12648,4.126953,3.1235218,2.1239948,1.1244678,0.12494087,0.1756981,0.22645533,0.27330816,0.3240654,0.37482262,0.6481308,0.92534333,1.1986516,1.475864,1.7491722,1.4016805,1.0502841,0.698888,0.3513962,0.0,0.0,0.0,0.0,0.0,0.0,1.5617609,3.1235218,4.689187,6.250948,7.812709,6.250948,4.689187,3.1235218,1.5617609,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.1756981,0.19912452,0.22645533,0.24988174,0.30063897,0.3513962,0.39824903,0.44900626,0.4997635,0.41386664,0.3240654,0.23816854,0.14836729,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.94876975,1.8389735,2.7252727,3.611572,4.5017757,5.0132523,5.5247293,6.036206,6.551587,7.0630636,5.64967,4.2362766,2.8267872,1.4133936,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,1.2494087,2.1864653,3.1235218,4.0605783,5.001539,7.211431,9.425227,11.639023,13.848915,16.062712,13.388195,10.71368,8.039165,5.3607445,2.6862288,2.736986,2.787743,2.8385005,2.8892577,2.9361105,2.35045,1.7608855,1.175225,0.58566034,0.0,1.4133936,2.8267872,4.2362766,5.64967,7.0630636,5.9268827,4.786797,3.6506162,2.5105307,1.3743496,4.5252023,7.676055,10.826907,13.973856,17.124708,15.961197,14.801589,13.638077,12.4745655,11.311053,12.923572,14.53609,16.148607,17.761126,19.373644,15.551234,11.72492,7.898606,4.0761957,0.24988174,1.43682,2.6237583,3.8106966,5.001539,6.1884775,5.1108627,4.037152,2.9634414,1.8858263,0.81211567,0.74964523,0.6871748,0.62470436,0.5622339,0.4997635,2.900971,5.298274,7.699481,10.100689,12.501896,15.988527,19.475159,22.96179,26.448421,29.938957,30.876013,31.81307,32.750126,33.687183,34.62424,32.94925,31.274261,29.599274,27.924286,26.249296,28.42405,30.5988,32.773552,34.948303,37.12306,31.188366,25.24977,19.311174,13.376482,7.437886,6.13772,4.8375545,3.5373883,2.2372224,0.93705654,0.8355421,0.737932,0.63641757,0.5388075,0.43729305,0.3631094,0.28892577,0.21083772,0.13665408,0.062470436,0.76135844,1.4641509,2.1630387,2.8619268,3.5608149,4.138666,4.7126136,5.2865605,5.8644123,6.4383593,9.550168,12.661977,15.773785,18.889498,22.001307,23.000834,24.00036,24.999887,25.999414,26.998941,24.925705,22.848562,20.775324,18.698183,16.624945,22.200432,27.775917,33.351402,38.92689,44.498474,42.0387,39.57502,37.111343,34.65157,32.187893,27.123882,22.063778,16.999767,11.935758,6.8756523,5.5013027,4.126953,2.7486992,1.3743496,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22645533,0.44900626,0.6754616,0.9019169,1.1244678,1.7765031,2.4246337,3.076669,3.7247996,4.376835,5.2865605,6.2001905,7.113821,8.023546,8.937177,7.1489606,5.3607445,3.5764325,1.7882162,0.0,0.27330816,0.5505207,0.8238289,1.1010414,1.3743496,1.1010414,0.8238289,0.5505207,0.27330816,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6871748,1.3743496,2.0615244,2.7486992,3.435874,3.5373883,3.638903,3.736513,3.8380275,3.9356375,7.5394006,11.139259,14.739119,18.338978,21.938837,17.663515,13.388195,9.112875,4.8375545,0.5622339,3.8263142,7.08649,10.350571,13.610746,16.874826,13.501423,10.124115,6.7507114,3.3734035,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.41386664,0.8238289,1.2376955,1.6515622,2.0615244,1.8233559,1.5890918,1.3509232,1.1127546,0.8745861,0.77307165,0.6754616,0.57394713,0.47633708,0.37482262,0.3513962,0.3240654,0.30063897,0.27330816,0.24988174,0.27330816,0.30063897,0.3240654,0.3513962,0.37482262,0.3357786,0.30063897,0.26159495,0.22645533,0.18741131,0.3357786,0.48805028,0.63641757,0.78868926,0.93705654,0.78868926,0.63641757,0.48805028,0.3357786,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.19912452,0.27330816,0.3513962,0.42557985,0.4997635,0.5231899,0.5505207,0.57394713,0.60127795,0.62470436,0.80040246,0.97610056,1.1517987,1.3235924,1.4992905,1.3626363,1.2259823,1.0893283,0.94876975,0.81211567,0.74964523,0.6871748,0.62470436,0.5622339,0.4997635,0.47633708,0.44900626,0.42557985,0.39824903,0.37482262,0.44900626,0.5231899,0.60127795,0.6754616,0.74964523,0.80040246,0.8511597,0.9019169,0.94876975,0.999527,0.93705654,0.8745861,0.81211567,0.74964523,0.6871748,0.698888,0.7106012,0.7262188,0.737932,0.74964523,0.9019169,1.0502841,1.1986516,1.3509232,1.4992905,1.4251068,1.3509232,1.2767396,1.1986516,1.1244678,1.261122,1.4016805,1.5383345,1.6749885,1.8116426,1.9873407,2.1630387,2.338737,2.514435,2.6862288,8.125061,6.617962,5.1108627,3.6037633,2.096664,0.58566034,0.8980125,1.2064602,1.5188124,1.8272603,2.135708,1.8858263,1.6359446,1.3860629,1.1361811,0.8862993,0.7106012,0.5309987,0.3553006,0.1756981,0.0,0.0,0.0,0.0,0.0,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,0.3240654,0.24988174,0.1756981,0.10151446,0.023426414,0.24597734,0.46462387,0.6832704,0.9058213,1.1244678,3.0415294,4.9546866,6.871748,8.784905,10.698062,9.589212,8.476458,7.363703,6.250948,5.138193,5.009348,4.884407,4.755562,4.6267166,4.5017757,7.113821,9.729771,12.34572,14.96167,17.573715,19.330696,21.083773,22.840754,24.59383,26.350811,25.956467,25.558218,25.163872,24.769527,24.375183,25.608974,26.84667,28.080462,29.314253,30.551949,27.475279,24.39861,21.325846,18.249176,15.176412,16.43363,17.694752,18.955873,20.21309,21.474213,22.37613,23.274141,24.17606,25.074072,25.975988,20.8417,15.711315,10.577025,5.446641,0.31235218,1.678893,3.0415294,4.40807,5.7707067,7.137247,6.477403,5.8175592,5.1577153,4.4978714,3.8380275,6.0323014,8.226576,10.42085,12.619028,14.813302,13.856724,12.89624,11.939662,10.983084,10.0265045,8.421796,6.8209906,5.2162814,3.6154766,2.0107672,1.9834363,1.9561055,1.9287747,1.901444,1.8741131,2.7565079,3.638903,4.521298,5.4036927,6.2860875,6.688241,7.08649,7.4886436,7.8868923,8.289046,7.3910336,6.493021,5.5950084,4.6969957,3.7989833,4.6657605,5.5286336,6.395411,7.2582836,8.125061,7.519879,6.914696,6.309514,5.704332,5.099149,5.1186714,5.134289,5.153811,5.169429,5.1889505,5.794133,6.3993154,7.000593,7.605776,8.210958,8.468649,8.726339,8.98403,9.24172,9.499411,9.448653,9.393991,9.343235,9.288573,9.237816,8.140678,7.0474463,5.9542136,4.8570766,3.7638438,3.310933,2.8580225,2.4051118,1.9522011,1.4992905,1.5812829,1.6593709,1.7413634,1.8194515,1.901444,1.756981,1.6164225,1.4719596,1.3314011,1.1869383,1.1088502,1.0268579,0.94876975,0.8667773,0.78868926,1.8819219,2.97125,4.0644827,5.1577153,6.250948,5.0718184,3.8965936,2.717464,1.5383345,0.3631094,0.29283017,0.22255093,0.15227169,0.08199245,0.011713207,0.031235218,0.05075723,0.07418364,0.093705654,0.113227665,0.15617609,0.20302892,0.24597734,0.29283017,0.3357786,0.3553006,0.3709182,0.39044023,0.40605783,0.42557985,0.359205,0.28892577,0.22255093,0.15617609,0.08589685,0.13274968,0.1756981,0.22255093,0.26940376,0.31235218,0.96829176,1.6281357,2.2840753,2.9439192,3.5998588,4.1035266,4.6110992,5.114767,5.618435,6.126007,5.0132523,3.9044023,2.795552,1.6867018,0.57394713,0.6832704,0.79649806,0.9058213,1.0151446,1.1244678,2.6823244,4.240181,5.7980375,7.355894,8.913751,9.698535,10.487225,11.275913,12.0606985,12.849388,11.490656,10.135828,8.777096,7.4183645,6.0635366,5.388075,4.716518,4.044961,3.3734035,2.7018464,2.2020829,1.7062237,1.2064602,0.7106012,0.21083772,1.4836729,2.7565079,4.029343,5.3021784,6.575013,5.55206,4.5291066,3.506153,2.4831998,1.4641509,4.650143,7.8361354,11.0260315,14.212025,17.40192,16.378967,15.356014,14.33306,13.310107,12.287154,13.005564,13.727879,14.446288,15.168603,15.8870125,12.767395,9.647778,6.5281606,3.408543,0.28892577,1.261122,2.233318,3.2055142,4.1777105,5.1499066,4.251894,3.349977,2.4480603,1.5500476,0.6481308,0.679366,0.7106012,0.7418364,0.76916724,0.80040246,2.8306916,4.8648853,6.899079,8.929368,10.963562,14.348679,17.7377,21.12672,24.511837,27.900858,29.177599,30.454338,31.731077,33.011723,34.28846,33.04686,31.801357,30.559757,29.318157,28.076557,29.6227,31.168842,32.71889,34.265034,35.811176,30.57147,25.327858,20.084246,14.840633,9.600925,7.9766936,6.356367,4.732136,3.1118085,1.4875772,1.397776,1.3079748,1.2181735,1.1283722,1.038571,1.0580931,1.0815194,1.1049459,1.1283722,1.1517987,1.678893,2.2098918,2.7408905,3.2718892,3.7989833,4.0761957,4.3534083,4.630621,4.911738,5.1889505,7.7970915,10.401327,13.009468,15.617609,18.22575,19.846077,21.470308,23.090635,24.714867,26.339098,24.351757,22.364416,20.37317,18.38583,16.398489,20.240421,24.07845,27.92038,31.758408,35.600338,33.82774,32.05514,30.282543,28.509945,26.737347,23.207767,19.678188,16.148607,12.619028,9.085544,7.269997,5.45445,3.6349986,1.815547,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.25378615,0.43338865,0.61689556,0.79649806,0.97610056,1.6945106,2.416825,3.135235,3.853645,4.575959,5.2084727,5.840986,6.473499,7.1060123,7.7385254,6.364176,4.9937305,3.619381,2.2489357,0.8745861,0.92143893,0.96438736,1.0112402,1.0541886,1.1010414,0.97610056,0.8550641,0.7340276,0.60908675,0.48805028,0.39044023,0.29283017,0.19522011,0.09761006,0.0,0.0,0.0,0.0,0.0,0.0,0.5505207,1.1010414,1.6515622,2.1981785,2.7486992,2.8345962,2.920493,3.0063896,3.0883822,3.174279,6.211904,9.245625,12.2793455,15.31697,18.35069,15.1061325,11.8654785,8.62092,5.380266,2.135708,4.4119744,6.6843367,8.956698,11.229061,13.501423,11.268105,9.034787,6.801469,4.5681505,2.338737,1.8702087,1.4016805,0.93315214,0.46852827,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.058566034,0.06637484,0.07418364,0.078088045,0.08589685,0.40996224,0.7340276,1.0541886,1.3782539,1.698415,1.5461433,1.3899672,1.2337911,1.0815194,0.92534333,0.8628729,0.80040246,0.737932,0.6754616,0.61299115,0.57394713,0.5388075,0.4997635,0.46071947,0.42557985,0.41777104,0.40996224,0.40215343,0.39434463,0.38653582,0.3513962,0.31235218,0.27330816,0.23816854,0.19912452,0.31235218,0.42557985,0.5388075,0.6481308,0.76135844,0.6637484,0.5661383,0.46852827,0.3709182,0.27330816,0.24597734,0.21864653,0.19131571,0.1639849,0.13665408,0.21474212,0.29283017,0.3709182,0.44900626,0.5231899,0.5544251,0.58175594,0.60908675,0.63641757,0.6637484,0.8238289,0.98390937,1.1439898,1.3040704,1.4641509,1.3509232,1.2415999,1.1322767,1.0229534,0.9136301,0.8316377,0.74574083,0.6637484,0.58175594,0.4997635,0.46852827,0.44119745,0.40996224,0.37872702,0.3513962,0.41386664,0.47633708,0.5388075,0.60127795,0.6637484,0.7027924,0.7418364,0.78088045,0.8238289,0.8628729,0.8160201,0.76916724,0.71841,0.6715572,0.62470436,0.63641757,0.6442264,0.6559396,0.6637484,0.6754616,0.80430686,0.92924774,1.0580931,1.1869383,1.3118792,1.2572175,1.2025559,1.1478943,1.0932326,1.038571,1.1439898,1.2494087,1.3509232,1.456342,1.5617609,1.6945106,1.8272603,1.9600099,2.0927596,2.2255092,8.062591,6.571109,5.083532,3.59205,2.1005683,0.61299115,1.0073358,1.4016805,1.796025,2.194274,2.5886188,2.4246337,2.260649,2.1005683,1.9365835,1.7765031,1.4212024,1.0659018,0.7106012,0.3553006,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.339683,0.62860876,0.92143893,1.2103647,1.4992905,3.240654,4.985922,6.727285,8.468649,10.213917,9.499411,8.78881,8.074304,7.363703,6.649197,6.36808,6.0908675,5.8097506,5.5286336,5.251421,7.6916723,10.135828,12.576079,15.020235,17.464392,19.045673,20.630861,22.21605,23.801235,25.386423,24.246338,23.106253,21.966167,20.826082,19.685997,20.556679,21.42736,22.29804,23.168722,24.0355,22.462027,20.888552,19.311174,17.7377,16.164225,17.218414,18.276506,19.3346,20.392693,21.450787,21.087677,20.724567,20.361458,19.998348,19.639143,15.773785,11.908427,8.043069,4.1777105,0.31235218,3.1039999,5.8956475,8.691199,11.482847,14.274494,12.244205,10.2100115,8.175818,6.1455293,4.1113358,5.5169206,6.918601,8.320281,9.721962,11.123642,10.573121,10.018696,9.468176,8.913751,8.36323,7.1450562,5.9268827,4.7087092,3.4905357,2.2762666,2.1318035,1.9912452,1.8467822,1.7062237,1.5617609,3.2289407,4.892216,6.559396,8.2226715,9.885946,9.698535,9.511124,9.323712,9.136301,8.94889,8.066495,7.1841,6.3017054,5.4193106,4.5369153,5.267039,5.997162,6.727285,7.4574084,8.187531,7.4144597,6.6413884,5.8683167,5.099149,4.3260775,4.3455997,4.369026,4.3924527,4.415879,4.4393053,5.9464045,7.4574084,8.968412,10.479416,11.986515,13.040704,14.090988,15.145176,16.199366,17.24965,16.46877,15.6917925,14.9109125,14.130032,13.349152,12.158309,10.971371,9.780528,8.589685,7.3988423,6.446168,5.4895897,4.5369153,3.5803368,2.6237583,2.5105307,2.3933985,2.280171,2.1669433,2.0498111,2.1161861,2.1786566,2.2450314,2.3114061,2.3738766,2.2137961,2.0537157,1.893635,1.7335546,1.5734742,2.1981785,2.8189783,3.4436827,4.0644827,4.689187,3.8965936,3.1039999,2.3114061,1.5188124,0.7262188,0.58566034,0.44510186,0.30454338,0.1639849,0.023426414,0.039044023,0.05466163,0.07027924,0.08589685,0.10151446,0.1639849,0.23035973,0.29673457,0.359205,0.42557985,0.40996224,0.39434463,0.37872702,0.3631094,0.3513962,0.30063897,0.25378615,0.20693332,0.16008049,0.113227665,0.20302892,0.29283017,0.38263142,0.47243267,0.5622339,0.9917182,1.4172981,1.8467822,2.2723622,2.7018464,3.1977055,3.6935644,4.193328,4.689187,5.1889505,4.380739,3.5725281,2.7643168,1.9561055,1.1517987,1.3079748,1.4641509,1.6242313,1.7804074,1.9365835,4.11524,6.2938967,8.468649,10.647305,12.825961,12.185639,11.549222,10.912805,10.276386,9.636065,9.597021,9.557977,9.518932,9.475985,9.43694,8.043069,6.649197,5.251421,3.8575494,2.463678,2.0537157,1.6476578,1.2415999,0.8316377,0.42557985,1.5578566,2.690133,3.8224099,4.9546866,6.086963,5.181142,4.271416,3.3655949,2.455869,1.5500476,4.775084,8.00012,11.225157,14.450192,17.675228,16.792833,15.9104395,15.028045,14.145649,13.263254,13.091461,12.915763,12.743969,12.572175,12.400381,9.983557,7.570636,5.153811,2.7408905,0.3240654,1.0815194,1.8389735,2.5964274,3.3538816,4.1113358,3.3890212,2.6628022,1.9365835,1.2142692,0.48805028,0.60908675,0.7340276,0.8550641,0.97610056,1.1010414,2.7643168,4.4314966,6.094772,7.7619514,9.425227,12.712734,16.00024,19.287746,22.575254,25.86276,27.479183,29.095606,30.715933,32.332355,33.948776,33.140568,32.32845,31.520239,30.708124,29.899912,30.821352,31.738886,32.660324,33.581764,34.4993,29.95067,25.405945,20.857317,16.30869,11.763964,9.815667,7.871275,5.9268827,3.9824903,2.0380979,1.9561055,1.8780174,1.796025,1.717937,1.6359446,1.756981,1.8780174,1.999054,2.1161861,2.2372224,2.5964274,2.9556324,3.3187418,3.677947,4.037152,4.01763,3.998108,3.978586,3.959064,3.9356375,6.04011,8.140678,10.2451515,12.34572,14.450192,16.695225,18.940256,21.185287,23.430319,25.67535,23.773905,21.876366,19.974922,18.073479,16.175938,18.28041,20.384884,22.489357,24.59383,26.698303,25.616783,24.535263,23.453745,22.36832,21.2868,19.29165,17.292597,15.293544,13.298394,11.29934,9.0386915,6.7819467,4.521298,2.260649,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.28502136,0.42167544,0.5544251,0.6910792,0.8238289,1.6164225,2.4051118,3.193801,3.9863946,4.775084,5.12648,5.481781,5.833177,6.184573,6.5359693,5.579391,4.6228123,3.6662338,2.7057507,1.7491722,1.5656652,1.3782539,1.1947471,1.0112402,0.8238289,0.8550641,0.8862993,0.9136301,0.94486535,0.97610056,0.78088045,0.58566034,0.39044023,0.19522011,0.0,0.0,0.0,0.0,0.0,0.0,0.41386664,0.8238289,1.2376955,1.6515622,2.0615244,2.1318035,2.2020829,2.2723622,2.3426414,2.4129205,4.884407,7.3519893,9.823476,12.291059,14.762545,12.552653,10.342762,8.13287,5.9229784,3.7130866,4.9937305,6.278279,7.558923,8.843472,10.124115,9.034787,7.9454584,6.8561306,5.7668023,4.6735697,3.7404175,2.803361,1.8702087,0.93315214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.113227665,0.12884527,0.14446288,0.16008049,0.1756981,0.40605783,0.64032197,0.8706817,1.1049459,1.33921,1.2650263,1.1908426,1.1205635,1.0463798,0.97610056,0.94876975,0.92534333,0.9019169,0.8745861,0.8511597,0.80040246,0.74964523,0.698888,0.6481308,0.60127795,0.5583295,0.5192855,0.48024148,0.44119745,0.39824903,0.3631094,0.3240654,0.28892577,0.24988174,0.21083772,0.28892577,0.3631094,0.43729305,0.5114767,0.58566034,0.5427119,0.4958591,0.45291066,0.40605783,0.3631094,0.32016098,0.27721256,0.23426414,0.19131571,0.14836729,0.23035973,0.30844778,0.39044023,0.46852827,0.5505207,0.58175594,0.60908675,0.64032197,0.6715572,0.698888,0.8433509,0.9917182,1.1361811,1.2806439,1.4251068,1.3431144,1.261122,1.1791295,1.0932326,1.0112402,0.9097257,0.80821127,0.7066968,0.60127795,0.4997635,0.46462387,0.42948425,0.39434463,0.359205,0.3240654,0.37482262,0.42557985,0.47633708,0.5231899,0.57394713,0.60518235,0.63641757,0.6637484,0.6949836,0.7262188,0.6910792,0.659844,0.62860876,0.59346914,0.5622339,0.5700427,0.57785153,0.58566034,0.59346914,0.60127795,0.7066968,0.80821127,0.9136301,1.0190489,1.1244678,1.0893283,1.0541886,1.0190489,0.98390937,0.94876975,1.0229534,1.0932326,1.1674163,1.2415999,1.3118792,1.4016805,1.4914817,1.5812829,1.6710842,1.7608855,8.00012,6.5281606,5.056201,3.5842414,2.1083772,0.63641757,1.116659,1.5969005,2.077142,2.5573835,3.0376248,2.9634414,2.8892577,2.8111696,2.736986,2.6628022,2.1318035,1.5969005,1.0659018,0.5309987,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.1756981,0.14836729,0.12494087,0.10151446,0.07418364,0.43338865,0.79649806,1.1557031,1.5149081,1.8741131,3.4436827,5.0132523,6.5867267,8.156297,9.725866,9.413514,9.101162,8.78881,8.476458,8.164105,7.7307167,7.297328,6.8639393,6.434455,6.001066,8.269524,10.541886,12.810344,15.078801,17.351164,18.764557,20.181856,21.59525,23.008642,24.425941,22.540113,20.654287,18.768461,16.88654,15.000713,15.504381,16.008049,16.515621,17.019289,17.522957,17.448774,17.37459,17.300406,17.226223,17.148134,18.003199,18.858263,19.713327,20.568392,21.423454,19.799223,18.174992,16.55076,14.92653,13.298394,10.701966,8.105539,5.5091114,2.9087796,0.31235218,4.533011,8.75367,12.974329,17.191084,21.411741,18.007103,14.602465,11.197825,7.793187,4.388548,4.997635,5.606722,6.2158084,6.8287997,7.437886,7.289519,7.141152,6.996689,6.8483214,6.699954,5.8683167,5.036679,4.2011366,3.3694992,2.5378613,2.280171,2.0224805,1.7647898,1.5070993,1.2494087,3.697469,6.1455293,8.59359,11.04165,13.4858055,12.712734,11.935758,11.162686,10.38571,9.612638,8.745861,7.8790836,7.008402,6.141625,5.2748475,5.8683167,6.46569,7.0591593,7.656533,8.250002,7.309041,6.36808,5.4310236,4.4900627,3.5491016,3.5764325,3.6037633,3.631094,3.6584249,3.6857557,6.1025805,8.519405,10.932326,13.349152,15.762072,17.608854,19.459541,21.306324,23.153105,24.999887,23.492788,21.98569,20.47859,18.97149,17.464392,16.175938,14.89139,13.606842,12.322293,11.037745,9.581403,8.121157,6.6648145,5.2084727,3.7482262,3.4397783,3.1313305,2.8189783,2.5105307,2.1981785,2.4714866,2.7447948,3.018103,3.2914112,3.5608149,3.3226464,3.084478,2.8424048,2.6042364,2.3621633,2.514435,2.6667068,2.8189783,2.97125,3.1235218,2.717464,2.3114061,1.901444,1.4953861,1.0893283,0.8784905,0.6676528,0.45681506,0.24597734,0.039044023,0.046852827,0.058566034,0.06637484,0.078088045,0.08589685,0.1717937,0.25769055,0.3435874,0.42557985,0.5114767,0.46462387,0.41777104,0.3709182,0.3240654,0.27330816,0.24597734,0.21864653,0.19131571,0.1639849,0.13665408,0.27330816,0.40605783,0.5427119,0.679366,0.81211567,1.0112402,1.2064602,1.4055848,1.6008049,1.7999294,2.2918842,2.7799344,3.2718892,3.7599394,4.251894,3.7443218,3.240654,2.7330816,2.2294137,1.7257458,1.9287747,2.135708,2.338737,2.5456703,2.7486992,5.548156,8.343708,11.143164,13.938716,16.738173,14.676648,12.611219,10.549695,8.488171,6.426646,7.703386,8.980125,10.256865,11.533605,12.814248,10.694158,8.577971,6.461786,4.3416953,2.2255092,1.9092526,1.5890918,1.2728351,0.95657855,0.63641757,1.6281357,2.6237583,3.6154766,4.607195,5.5989127,4.806319,4.0137253,3.2211318,2.4285383,1.6359446,4.900025,8.164105,11.424281,14.688361,17.948538,17.206701,16.464865,15.723028,14.981192,14.239355,13.173453,12.107552,11.04165,9.975748,8.913751,7.2036223,5.493494,3.7833657,2.0732377,0.3631094,0.9058213,1.4485333,1.9912452,2.533957,3.076669,2.5261483,1.9756275,1.4251068,0.8745861,0.3240654,0.5388075,0.75354964,0.96829176,1.1869383,1.4016805,2.697942,3.9942036,5.2943697,6.590631,7.8868923,11.076789,14.262781,17.448774,20.63867,23.824663,25.780767,27.740778,29.696884,31.656893,33.613,33.234272,32.85945,32.48072,32.101994,31.723269,32.016098,32.30893,32.601757,32.89459,33.18742,29.333775,25.484034,21.630388,17.776743,13.927003,11.6585455,9.390087,7.1216297,4.853172,2.5886188,2.5183394,2.4480603,2.377781,2.3075018,2.2372224,2.455869,2.6706111,2.8892577,3.1079042,3.3265507,3.513962,3.7052777,3.8965936,4.084005,4.2753205,3.959064,3.638903,3.3226464,3.0063896,2.6862288,4.283129,5.883934,7.480835,9.077735,10.674636,13.544372,16.410202,19.276033,22.14577,25.0116,23.199959,21.388315,19.576674,17.761126,15.949483,16.320402,16.69132,17.058334,17.429253,17.800169,17.405825,17.015385,16.62104,16.2306,15.836256,15.371632,14.907008,14.442384,13.97776,13.513136,10.81129,8.109444,5.4036927,2.7018464,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.08980125,0.13665408,0.1796025,0.22645533,0.31625658,0.40605783,0.4958591,0.58566034,0.6754616,1.53443,2.3933985,3.2562714,4.11524,4.9742084,5.0483923,5.1186714,5.192855,5.263134,5.337318,4.794606,4.251894,3.7091823,3.1664703,2.6237583,2.2098918,1.796025,1.3782539,0.96438736,0.5505207,0.7340276,0.9136301,1.097137,1.2806439,1.4641509,1.1713207,0.8784905,0.58566034,0.29283017,0.0,0.0,0.0,0.0,0.0,0.0,0.27330816,0.5505207,0.8238289,1.1010414,1.3743496,1.4290112,1.4836729,1.5383345,1.5969005,1.6515622,3.5569105,5.4583545,7.363703,9.269051,11.174399,9.999174,8.8200445,7.6409154,6.46569,5.2865605,5.579391,5.872221,6.165051,6.4578815,6.7507114,6.801469,6.8561306,6.9068875,6.9615493,7.012306,5.610626,4.2089458,2.803361,1.4016805,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.1717937,0.19522011,0.21864653,0.23816854,0.26159495,0.40605783,0.5466163,0.6910792,0.8316377,0.97610056,0.98390937,0.9956226,1.0034313,1.0151446,1.0268579,1.038571,1.0502841,1.0619974,1.0737107,1.0893283,1.0268579,0.96438736,0.9019169,0.8394465,0.77307165,0.7027924,0.62860876,0.5583295,0.48414588,0.41386664,0.37482262,0.3357786,0.30063897,0.26159495,0.22645533,0.26159495,0.30063897,0.3357786,0.37482262,0.41386664,0.42167544,0.42557985,0.43338865,0.44119745,0.44900626,0.39434463,0.3357786,0.27721256,0.21864653,0.1639849,0.24597734,0.3279698,0.40996224,0.49195468,0.57394713,0.60908675,0.64032197,0.6715572,0.7066968,0.737932,0.8667773,0.9956226,1.1283722,1.2572175,1.3860629,1.3314011,1.2767396,1.2220778,1.1674163,1.1127546,0.9917182,0.8667773,0.74574083,0.62079996,0.4997635,0.46071947,0.42167544,0.37872702,0.339683,0.30063897,0.3357786,0.37482262,0.41386664,0.44900626,0.48805028,0.5075723,0.5270943,0.5466163,0.5661383,0.58566034,0.5700427,0.5544251,0.5349031,0.5192855,0.4997635,0.5036679,0.5114767,0.5153811,0.5192855,0.5231899,0.60908675,0.6910792,0.77307165,0.8550641,0.93705654,0.92143893,0.9058213,0.8941081,0.8784905,0.8628729,0.9019169,0.94096094,0.98390937,1.0229534,1.0619974,1.1088502,1.1557031,1.2064602,1.2533131,1.3001659,7.9376497,6.481308,5.02887,3.5725281,2.1161861,0.6637484,1.2259823,1.7921207,2.358259,2.9243972,3.4866312,3.4983444,3.513962,3.5256753,3.5373883,3.5491016,2.8385005,2.1318035,1.4212024,0.7106012,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.5309987,0.96048295,1.3899672,1.8194515,2.2489357,3.6467118,5.044488,6.4422636,7.8400397,9.237816,9.323712,9.413514,9.499411,9.589212,9.675109,9.089449,8.503788,7.918128,7.336372,6.7507114,8.847376,10.944039,13.040704,15.141272,17.237936,18.48344,19.728945,20.97445,22.21605,23.461554,20.83389,18.202324,15.570756,12.943093,10.311526,10.452085,10.592644,10.733202,10.87376,11.014318,12.435521,13.860628,15.285735,16.710842,18.135948,18.791887,19.443924,20.095959,20.747993,21.400028,18.51077,15.625418,12.73616,9.850807,6.9615493,5.6340523,4.3026514,2.97125,1.6437533,0.31235218,5.958118,11.607788,17.253553,22.903223,28.548988,23.773905,18.994917,14.215929,9.440845,4.661856,4.478349,4.298747,4.11524,3.9317331,3.7482262,4.0059166,4.263607,4.521298,4.7789884,5.036679,4.591577,4.142571,3.6935644,3.2484627,2.7994564,2.4285383,2.0537157,1.6827974,1.3118792,0.93705654,4.165997,7.3988423,10.627783,13.856724,17.085665,15.726933,14.364296,13.001659,11.639023,10.276386,9.421323,8.570163,7.719003,6.8639393,6.012779,6.473499,6.9342184,7.3910336,7.8517528,8.312472,7.2036223,6.098676,4.989826,3.8809757,2.77603,2.8072653,2.8385005,2.87364,2.9048753,2.9361105,6.2587566,9.577498,12.89624,16.218887,19.537628,22.18091,24.82419,27.463566,30.106846,32.750126,30.516808,28.279585,26.046267,23.809046,21.575727,20.19357,18.815315,17.433157,16.054901,14.676648,12.716639,10.756628,8.796618,6.8366084,4.8765984,4.369026,3.8653584,3.3616903,2.854118,2.35045,2.8306916,3.310933,3.7911747,4.271416,4.7516575,4.4314966,4.1113358,3.7911747,3.4710135,3.1508527,2.8306916,2.514435,2.1981785,1.8819219,1.5617609,1.5383345,1.5188124,1.4953861,1.4719596,1.4485333,1.1713207,0.8902037,0.60908675,0.3318742,0.05075723,0.05466163,0.058566034,0.06637484,0.07027924,0.07418364,0.1796025,0.28502136,0.39044023,0.4958591,0.60127795,0.5192855,0.44119745,0.359205,0.28111696,0.19912452,0.19131571,0.1835069,0.1756981,0.1717937,0.1639849,0.3435874,0.5231899,0.7027924,0.8823949,1.0619974,1.0307622,0.9956226,0.96438736,0.93315214,0.9019169,1.3821584,1.8663043,2.3465457,2.8306916,3.310933,3.1118085,2.9087796,2.7057507,2.5027218,2.2996929,2.5534792,2.803361,3.057147,3.310933,3.5608149,6.9810715,10.397423,13.813775,17.234032,20.650383,17.163752,13.673217,10.186585,6.699954,3.213323,5.805846,8.402273,10.998701,13.591225,16.187653,13.349152,10.506746,7.6682463,4.825841,1.9873407,1.7608855,1.53443,1.3040704,1.077615,0.8511597,1.7023194,2.5534792,3.408543,4.2597027,5.1108627,4.435401,3.7560349,3.0805733,2.4012074,1.7257458,5.024966,8.324185,11.623405,14.92653,18.22575,17.620567,17.019289,16.41801,15.816733,15.211552,13.2554455,11.29934,9.339331,7.3832245,5.423215,4.4197836,3.416352,2.4090161,1.4055848,0.39824903,0.7262188,1.0541886,1.3821584,1.7101282,2.0380979,1.6632754,1.2884527,0.9136301,0.5388075,0.1639849,0.46852827,0.77697605,1.0854238,1.3938715,1.698415,2.631567,3.5608149,4.4900627,5.4193106,6.348558,9.43694,12.525322,15.613705,18.698183,21.786564,24.086258,26.382046,28.68174,30.977528,33.273315,33.331882,33.386543,33.441204,33.49587,33.55053,33.21475,32.87897,32.543194,32.21132,31.87554,28.716879,25.558218,22.40346,19.244799,16.086138,13.497519,10.9089,8.316377,5.727758,3.1391394,3.076669,3.018103,2.9556324,2.8970666,2.8385005,3.1508527,3.4671092,3.7833657,4.095718,4.4119744,4.4314966,4.4510183,4.474445,4.493967,4.513489,3.8965936,3.2836022,2.6667068,2.0537157,1.43682,2.5300527,3.6232853,4.716518,5.805846,6.899079,10.389614,13.88015,17.370686,20.861221,24.351757,22.62601,20.900265,19.174519,17.448774,15.726933,14.360392,12.993851,11.631214,10.264673,8.898132,9.198771,9.495506,9.792241,10.088976,10.38571,11.455516,12.521418,13.591225,14.657126,15.726933,12.579984,9.43694,6.289992,3.1430438,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.3435874,0.39044023,0.43338865,0.48024148,0.5231899,1.456342,2.3855898,3.3148375,4.2440853,5.173333,4.9663997,4.759466,4.552533,4.3455997,4.138666,4.009821,3.8809757,3.7560349,3.6271896,3.4983444,2.854118,2.2098918,1.5656652,0.92143893,0.27330816,0.60908675,0.94486535,1.2806439,1.6164225,1.9482968,1.5617609,1.1713207,0.78088045,0.39044023,0.0,0.0,0.0,0.0,0.0,0.0,0.13665408,0.27330816,0.41386664,0.5505207,0.6871748,0.7262188,0.76916724,0.80821127,0.8472553,0.8862993,2.2294137,3.5686235,4.9078336,6.2470436,7.5862536,7.4417906,7.297328,7.152865,7.008402,6.8639393,6.165051,5.466163,4.7711797,4.0722914,3.3734035,4.5681505,5.7668023,6.9615493,8.156297,9.351044,7.480835,5.610626,3.7404175,1.8702087,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.23035973,0.26159495,0.28892577,0.32016098,0.3513962,0.40215343,0.45681506,0.5075723,0.5583295,0.61299115,0.7066968,0.79649806,0.8902037,0.98390937,1.0737107,1.1244678,1.175225,1.2259823,1.2767396,1.3235924,1.2494087,1.175225,1.1010414,1.0268579,0.94876975,0.8433509,0.7418364,0.63641757,0.5309987,0.42557985,0.38653582,0.3513962,0.31235218,0.27330816,0.23816854,0.23816854,0.23816854,0.23816854,0.23816854,0.23816854,0.29673457,0.359205,0.41777104,0.47633708,0.5388075,0.46462387,0.39434463,0.32016098,0.24597734,0.1756981,0.26159495,0.3435874,0.42948425,0.5153811,0.60127795,0.63641757,0.6715572,0.7066968,0.7418364,0.77307165,0.8902037,1.0034313,1.1205635,1.2337911,1.3509232,1.3235924,1.2962615,1.2689307,1.2415999,1.2142692,1.0698062,0.92924774,0.78478485,0.6442264,0.4997635,0.45681506,0.40996224,0.3631094,0.32016098,0.27330816,0.30063897,0.3240654,0.3513962,0.37482262,0.39824903,0.40996224,0.42167544,0.42948425,0.44119745,0.44900626,0.44900626,0.44510186,0.44119745,0.44119745,0.43729305,0.44119745,0.44119745,0.44510186,0.44900626,0.44900626,0.5114767,0.5700427,0.62860876,0.6910792,0.74964523,0.75354964,0.76135844,0.76526284,0.76916724,0.77307165,0.78088045,0.78868926,0.79649806,0.80430686,0.81211567,0.8160201,0.8238289,0.8277333,0.8316377,0.8355421,7.8751793,6.4383593,5.001539,3.5608149,2.1239948,0.6871748,1.33921,1.9873407,2.639376,3.2875066,3.9356375,4.037152,4.138666,4.2362766,4.337791,4.4393053,3.5491016,2.6628022,1.7765031,0.8862993,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.62470436,1.1244678,1.6242313,2.1239948,2.6237583,3.8497405,5.0757227,6.3017054,7.523783,8.749765,9.237816,9.725866,10.213917,10.698062,11.186112,10.44818,9.714153,8.976221,8.238289,7.5003567,9.425227,11.350098,13.274967,15.199838,17.124708,18.19842,19.276033,20.349745,21.423454,22.50107,19.123762,15.750359,12.373051,8.999647,5.6262436,5.3997884,5.173333,4.950782,4.7243266,4.5017757,7.426173,10.350571,13.274967,16.199366,19.123762,19.576674,20.025679,20.474686,20.92369,21.376602,17.226223,13.075843,8.925464,4.775084,0.62470436,0.5622339,0.4997635,0.43729305,0.37482262,0.31235218,7.387129,14.461906,21.536682,28.61146,35.686237,29.536802,23.38737,17.237936,11.088503,4.939069,3.9629683,2.9868677,2.0107672,1.038571,0.062470436,0.7262188,1.3860629,2.0498111,2.7135596,3.3734035,3.310933,3.2484627,3.1859922,3.1235218,3.0610514,2.5769055,2.0888553,1.6008049,1.1127546,0.62470436,4.6384296,8.648251,12.661977,16.675701,20.689428,18.737226,16.788929,14.836729,12.888432,10.936231,10.100689,9.261242,8.4257,7.5862536,6.7507114,7.0747766,7.3988423,7.726812,8.050878,8.374943,7.098203,5.825368,4.548629,3.2757936,1.999054,2.0380979,2.0732377,2.1122816,2.1513257,2.1864653,6.4110284,10.6355915,14.864059,19.088623,23.313187,26.74906,30.188839,33.624714,37.06449,40.500366,37.536922,34.573483,31.613945,28.650503,25.687063,24.211199,22.739239,21.263374,19.78751,18.311647,15.851873,13.388195,10.924518,8.460839,6.001066,5.298274,4.5993857,3.900498,3.2016098,2.4988174,3.1859922,3.873167,4.564246,5.251421,5.938596,5.5364423,5.138193,4.73604,4.337791,3.9356375,3.1508527,2.3621633,1.5734742,0.78868926,0.0,0.3631094,0.7262188,1.0893283,1.4485333,1.8116426,1.4641509,1.1127546,0.76135844,0.41386664,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.18741131,0.31235218,0.43729305,0.5622339,0.6871748,0.57394713,0.46071947,0.3513962,0.23816854,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.41386664,0.63641757,0.8628729,1.0893283,1.3118792,1.0502841,0.78868926,0.5231899,0.26159495,0.0,0.47633708,0.94876975,1.4251068,1.901444,2.3738766,2.475391,2.5769055,2.6745155,2.77603,2.87364,3.174279,3.474918,3.775557,4.0761957,4.376835,8.413987,12.4511385,16.48829,20.525442,24.562595,19.650856,14.739119,9.823476,4.911738,0.0,3.912211,7.824422,11.736633,15.648844,19.561056,16.00024,12.439425,8.874706,5.3138914,1.7491722,1.6125181,1.475864,1.33921,1.1986516,1.0619974,1.7765031,2.4871042,3.2016098,3.912211,4.6267166,4.0605783,3.4983444,2.9361105,2.3738766,1.8116426,5.1499066,8.488171,11.826434,15.160794,18.499058,18.038338,17.573715,17.112995,16.64837,16.187653,13.337439,10.487225,7.6370106,4.786797,1.9365835,1.6359446,1.33921,1.038571,0.737932,0.43729305,0.5505207,0.6637484,0.77307165,0.8862993,0.999527,0.80040246,0.60127795,0.39824903,0.19912452,0.0,0.39824903,0.80040246,1.1986516,1.6008049,1.999054,2.5612879,3.1235218,3.6857557,4.251894,4.814128,7.800996,10.787864,13.774731,16.761599,19.748466,22.387842,25.023314,27.66269,30.29816,32.93754,33.425587,33.91364,34.401688,34.885834,35.373886,34.413403,33.449013,32.488533,31.524143,30.563662,28.099983,25.636305,23.176533,20.712854,18.249176,15.336493,12.423808,9.511124,6.5984397,3.6857557,3.638903,3.5881457,3.5373883,3.4866312,3.435874,3.8497405,4.263607,4.6735697,5.087436,5.5013027,5.349031,5.2006636,5.0483923,4.900025,4.7516575,3.8380275,2.9243972,2.0107672,1.1010414,0.18741131,0.77697605,1.3626363,1.9482968,2.5378613,3.1235218,7.238762,11.350098,15.461433,19.576674,23.68801,22.048159,20.412214,18.77627,17.136421,15.500477,12.400381,9.300286,6.2001905,3.1000953,0.0,0.9878138,1.9756275,2.9634414,3.951255,4.939069,7.5394006,10.135828,12.73616,15.336493,17.936825,14.348679,10.764437,7.1762915,3.5881457,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,1.3743496,2.3738766,3.3734035,4.376835,5.376362,4.8883114,4.4002614,3.912211,3.4241607,2.9361105,3.2250361,3.513962,3.7989833,4.087909,4.376835,3.4983444,2.6237583,1.7491722,0.8745861,0.0,0.48805028,0.97610056,1.4641509,1.9482968,2.436347,1.9482968,1.4641509,0.97610056,0.48805028,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.9019169,1.6749885,2.4519646,3.2250361,3.998108,4.8883114,5.774611,6.66091,7.551114,8.437413,6.7507114,5.0640097,3.3734035,1.6867018,0.0,2.338737,4.6735697,7.012306,9.351044,11.685876,9.351044,7.012306,4.6735697,2.338737,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.28892577,0.3240654,0.3631094,0.39824903,0.43729305,0.39824903,0.3631094,0.3240654,0.28892577,0.24988174,0.42557985,0.60127795,0.77307165,0.94876975,1.1244678,1.2142692,1.3001659,1.3860629,1.475864,1.5617609,1.475864,1.3860629,1.3001659,1.2142692,1.1244678,0.9878138,0.8511597,0.7106012,0.57394713,0.43729305,0.39824903,0.3631094,0.3240654,0.28892577,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,0.1756981,0.28892577,0.39824903,0.5114767,0.62470436,0.5388075,0.44900626,0.3631094,0.27330816,0.18741131,0.27330816,0.3631094,0.44900626,0.5388075,0.62470436,0.6637484,0.698888,0.737932,0.77307165,0.81211567,0.9136301,1.0112402,1.1127546,1.2142692,1.3118792,1.3118792,1.3118792,1.3118792,1.3118792,1.3118792,1.1517987,0.9878138,0.8238289,0.6637484,0.4997635,0.44900626,0.39824903,0.3513962,0.30063897,0.24988174,0.26159495,0.27330816,0.28892577,0.30063897,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.3240654,0.3357786,0.3513962,0.3631094,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.41386664,0.44900626,0.48805028,0.5231899,0.5622339,0.58566034,0.61299115,0.63641757,0.6637484,0.6871748,0.6637484,0.63641757,0.61299115,0.58566034,0.5622339,0.5231899,0.48805028,0.44900626,0.41386664,0.37482262,6.524256,5.7980375,5.0718184,4.3416953,3.6154766,2.8892577,3.5530062,4.220659,4.8883114,5.5559645,6.223617,6.001066,5.774611,5.548156,5.3256044,5.099149,4.2167544,3.3343596,2.4519646,1.5695697,0.6871748,0.5505207,0.41386664,0.27330816,0.13665408,0.0,0.046852827,0.093705654,0.14055848,0.19131571,0.23816854,0.21083772,0.18741131,0.1639849,0.13665408,0.113227665,0.57785153,1.0424755,1.5070993,1.9717231,2.436347,3.4436827,4.447114,5.45445,6.4578815,7.461313,8.628729,9.796145,10.963562,12.130978,13.298394,13.376482,13.45457,13.532659,13.610746,13.688834,14.957765,16.226696,17.495626,18.768461,20.037392,19.814842,19.59229,19.36974,19.147188,18.924637,17.26917,15.613705,13.958238,12.306676,10.651209,11.990419,13.329629,14.668839,16.008049,17.351164,16.976341,16.605423,16.2306,15.859682,15.488764,16.69913,17.905588,19.115953,20.326319,21.536682,17.476105,13.411622,9.351044,5.2865605,1.2259823,1.3314011,1.43682,1.5383345,1.6437533,1.7491722,7.1216297,12.494087,17.866545,23.239002,28.61146,23.703627,18.795792,13.887959,8.98403,4.0761957,3.2757936,2.475391,1.6749885,0.8745861,0.07418364,0.62470436,1.175225,1.7257458,2.2762666,2.8267872,2.7643168,2.7018464,2.639376,2.5769055,2.514435,2.6081407,2.7018464,2.795552,2.893162,2.9868677,6.282183,9.577498,12.872814,16.168129,19.463446,18.014912,16.56638,15.12175,13.673217,12.224684,10.869856,9.515028,8.160201,6.805373,5.4505453,5.840986,6.2353306,6.6257706,7.0201154,7.4144597,6.4110284,5.4115014,4.4119744,3.4124475,2.4129205,2.3035975,2.194274,2.0810463,1.9717231,1.8623998,5.860508,9.858616,13.856724,17.850927,21.849035,24.183868,26.5187,28.853533,31.188366,33.523197,31.000954,28.47871,25.956467,23.434223,20.911978,19.678188,18.448301,17.21451,15.980719,14.750832,13.048512,11.350098,9.651682,7.9493628,6.250948,5.446641,4.646239,3.8419318,3.0415294,2.2372224,3.349977,4.462732,5.575486,6.688241,7.800996,7.1606736,6.524256,5.8878384,5.251421,4.6110992,3.68966,2.7682211,1.8467822,0.92143893,0.0,0.28892577,0.58175594,0.8706817,1.1596074,1.4485333,1.1713207,0.8902037,0.60908675,0.3318742,0.05075723,0.08589685,0.12103647,0.15617609,0.19131571,0.22645533,0.37872702,0.5309987,0.6832704,0.8355421,0.9878138,1.0034313,1.0229534,1.038571,1.0580931,1.0737107,1.0190489,0.96438736,0.9097257,0.8550641,0.80040246,0.8628729,0.92534333,0.9878138,1.0502841,1.1127546,1.0346665,0.95657855,0.8784905,0.80430686,0.7262188,1.097137,1.4680552,1.8428779,2.2137961,2.5886188,2.533957,2.4792955,2.4207294,2.366068,2.3114061,2.6081407,2.9087796,3.2055142,3.5022488,3.7989833,7.355894,10.9089,14.465811,18.018816,21.575727,18.499058,15.418485,12.341816,9.265146,6.1884775,8.484266,10.77615,13.0719385,15.367727,17.663515,14.4970455,11.334479,8.16801,5.001539,1.8389735,1.8467822,1.8506867,1.8584955,1.8663043,1.8741131,2.2567444,2.639376,3.0220075,3.4046388,3.78727,3.3538816,2.9243972,2.4910088,2.05762,1.6242313,4.560342,7.4964523,10.4286585,13.364769,16.300879,16.46877,16.640562,16.808453,16.980246,17.148134,14.59856,12.0489855,9.499411,6.949836,4.4002614,3.6584249,2.9165885,2.1708477,1.4290112,0.6871748,1.0073358,1.3274968,1.6476578,1.9678187,2.2879796,1.8311646,1.3743496,0.9136301,0.45681506,0.0,0.32016098,0.64032197,0.96048295,1.2806439,1.6008049,2.1630387,2.7252727,3.2875066,3.8497405,4.4119744,6.6960497,8.976221,11.260296,13.544372,15.824542,18.436588,21.044727,23.656773,26.264914,28.876959,31.336733,33.80041,36.264088,38.72386,41.18754,39.92642,38.6692,37.408077,36.146957,34.885834,32.340164,29.790588,27.244919,24.69925,22.149673,18.90121,15.648844,12.400381,9.148014,5.899552,5.6223392,5.3451266,5.067914,4.7907014,4.513489,4.755562,5.001539,5.2475166,5.493494,5.735567,5.794133,5.8487945,5.903456,5.958118,6.012779,5.0132523,4.0137253,3.0141985,2.0107672,1.0112402,1.815547,2.6159496,3.4202564,4.220659,5.024966,8.296855,11.568744,14.844538,18.116426,21.388315,19.596195,17.804073,16.008049,14.215929,12.423808,9.940608,7.461313,4.9781127,2.494913,0.011713207,0.80040246,1.5890918,2.3738766,3.1625657,3.951255,7.2192397,10.491129,13.759113,17.031002,20.298986,17.456583,14.610273,11.763964,8.921559,6.0752497,5.7316628,5.388075,5.0483923,4.704805,4.3612175,3.5491016,2.736986,1.9248703,1.1127546,0.30063897,0.30844778,0.31625658,0.3240654,0.3318742,0.3357786,1.1283722,1.9209659,2.7135596,3.506153,4.298747,4.1777105,4.056674,3.9317331,3.8106966,3.6857557,3.873167,4.056674,4.2440853,4.4275923,4.6110992,3.892689,3.174279,2.4519646,1.7335546,1.0112402,1.2064602,1.4016805,1.5969005,1.7921207,1.9873407,2.6823244,3.377308,4.0722914,4.7672753,5.462259,6.094772,6.727285,7.3597984,7.9923115,8.624825,6.902983,5.181142,3.4593005,1.7335546,0.011713207,0.7418364,1.4680552,2.194274,2.9243972,3.6506162,3.9356375,4.220659,4.50568,4.7907014,5.0757227,5.74728,6.4188375,7.094299,7.7658563,8.437413,7.277806,6.1181984,4.958591,3.7989833,2.639376,4.009821,5.3841705,6.754616,8.128965,9.499411,7.5979667,5.700427,3.7989833,1.901444,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.47633708,0.57394713,0.6754616,0.77307165,0.8745861,0.80430686,0.7340276,0.6637484,0.59346914,0.5231899,0.61689556,0.7106012,0.80430686,0.8941081,0.9878138,1.1049459,1.2220778,1.33921,1.456342,1.5734742,1.5031948,1.43682,1.3665408,1.2962615,1.2259823,1.0619974,0.9019169,0.737932,0.57394713,0.41386664,0.37872702,0.3474918,0.31625658,0.28111696,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,0.15227169,0.24207294,0.3318742,0.42167544,0.5114767,0.44119745,0.3709182,0.30063897,0.23426414,0.1639849,0.23035973,0.29673457,0.3631094,0.43338865,0.4997635,0.5466163,0.58956474,0.63641757,0.679366,0.7262188,0.8433509,0.96438736,1.0854238,1.2064602,1.3235924,1.4172981,1.5110037,1.6008049,1.6945106,1.7882162,1.6281357,1.4719596,1.3157835,1.1557031,0.999527,0.8433509,0.6910792,0.5349031,0.37872702,0.22645533,0.23816854,0.24988174,0.26159495,0.27330816,0.28892577,0.28892577,0.29283017,0.29673457,0.29673457,0.30063897,0.31625658,0.3318742,0.3435874,0.359205,0.37482262,0.37872702,0.37872702,0.38263142,0.38653582,0.38653582,0.41386664,0.44119745,0.46852827,0.4958591,0.5231899,0.5427119,0.5583295,0.57785153,0.59346914,0.61299115,0.59346914,0.57394713,0.5544251,0.5309987,0.5114767,0.48024148,0.44900626,0.41386664,0.38263142,0.3513962,5.173333,5.1577153,5.138193,5.1225758,5.1069584,5.087436,5.7707067,6.4578815,7.141152,7.8283267,8.511597,7.9610763,7.4144597,6.8639393,6.3134184,5.7628975,4.884407,4.0059166,3.1313305,2.25284,1.3743496,1.1010414,0.8238289,0.5505207,0.27330816,0.0,0.093705654,0.19131571,0.28502136,0.37872702,0.47633708,0.39824903,0.3240654,0.24988174,0.1756981,0.10151446,0.5309987,0.96048295,1.3899672,1.8194515,2.2489357,3.0337205,3.8185053,4.60329,5.388075,6.1767645,8.023546,9.870329,11.717112,13.563893,15.410676,16.304783,17.198893,18.089096,18.983204,19.873407,20.490303,21.103294,21.72019,22.333181,22.950077,21.431265,19.908546,18.389734,16.870922,15.348206,15.41458,15.480955,15.543426,15.6098,15.676175,18.58105,21.485926,24.3908,27.295675,30.200552,26.530413,22.860275,19.190138,15.519999,11.849861,13.821584,15.789403,17.761126,19.728945,21.700668,17.725986,13.751305,9.776623,5.7980375,1.8233559,2.096664,2.3699722,2.6432803,2.9165885,3.1859922,6.8561306,10.526268,14.196406,17.866545,21.536682,17.874353,14.208119,10.541886,6.8756523,3.213323,2.5886188,1.9639144,1.33921,0.7106012,0.08589685,0.5231899,0.96438736,1.4016805,1.8389735,2.2762666,2.2137961,2.1513257,2.0888553,2.0263848,1.9639144,2.639376,3.3187418,3.9942036,4.6735697,5.349031,7.9259367,10.506746,13.083652,15.660558,18.237463,17.292597,16.347733,15.402867,14.458001,13.513136,11.639023,9.768814,7.8947015,6.0205884,4.1503797,4.6110992,5.0718184,5.5286336,5.989353,6.4500723,5.7238536,5.001539,4.2753205,3.5491016,2.8267872,2.5690966,2.3114061,2.0537157,1.796025,1.5383345,5.3060827,9.077735,12.849388,16.617136,20.388788,21.618675,22.852467,24.086258,25.316145,26.549934,24.46889,22.383938,20.30289,18.221846,16.136894,15.14908,14.157363,13.165645,12.177831,11.186112,10.249056,9.311999,8.374943,7.437886,6.5008297,5.5950084,4.689187,3.7833657,2.8814487,1.9756275,3.513962,5.0483923,6.5867267,8.125061,9.663396,8.78881,7.914223,7.0357327,6.1611466,5.2865605,4.2284675,3.174279,2.1161861,1.0580931,0.0,0.21864653,0.43338865,0.6520352,0.8706817,1.0893283,0.8784905,0.6676528,0.45681506,0.24597734,0.039044023,0.10932326,0.1756981,0.24597734,0.31625658,0.38653582,0.5661383,0.74574083,0.92924774,1.1088502,1.2884527,1.43682,1.5812829,1.7296503,1.8780174,2.0263848,1.901444,1.7804074,1.6593709,1.53443,1.4133936,1.3118792,1.2142692,1.1127546,1.0112402,0.9136301,1.0190489,1.1283722,1.2337911,1.3431144,1.4485333,1.7218413,1.9912452,2.260649,2.5300527,2.7994564,2.5886188,2.3816853,2.1708477,1.9600099,1.7491722,2.0459068,2.338737,2.6354716,2.9283018,3.2250361,6.297801,9.370565,12.44333,15.516094,18.58886,17.343355,16.101755,14.860155,13.618555,12.376955,13.052417,13.731783,14.407245,15.086611,15.762072,12.993851,10.22563,7.461313,4.6930914,1.9248703,2.077142,2.2294137,2.3816853,2.533957,2.6862288,2.7408905,2.7916477,2.8463092,2.8970666,2.951728,2.6471848,2.3465457,2.0420024,1.7413634,1.43682,3.970777,6.5008297,9.034787,11.568744,14.098797,14.903104,15.7035055,16.507812,17.308216,18.112522,15.863586,13.610746,11.361811,9.112875,6.8639393,5.677001,4.493967,3.3070288,2.1239948,0.93705654,1.4641509,1.9912452,2.5183394,3.049338,3.5764325,2.8619268,2.1435168,1.4290112,0.7145056,0.0,0.23816854,0.48024148,0.71841,0.96048295,1.1986516,1.7608855,2.3231194,2.8892577,3.4514916,4.0137253,5.591104,7.168483,8.745861,10.323239,11.900618,14.481428,17.066143,19.646952,22.231667,24.812477,29.251781,33.687183,38.126488,42.56189,47.001194,45.443336,43.885483,42.327625,40.769768,39.21191,36.580345,33.948776,31.313307,28.68174,26.05017,22.462027,18.87388,15.285735,11.701493,8.113348,7.605776,7.1021075,6.5984397,6.0908675,5.5871997,5.6652875,5.743376,5.8214636,5.8956475,5.9737353,6.2353306,6.4969254,6.754616,7.016211,7.2739015,6.1884775,5.099149,4.0137253,2.9243972,1.8389735,2.854118,3.873167,4.8883114,5.9073606,6.9264097,9.358852,11.791295,14.223738,16.65618,19.088623,17.140326,15.192029,13.243732,11.29934,9.351044,7.4847393,5.618435,3.7560349,1.8897307,0.023426414,0.61299115,1.1986516,1.7882162,2.3738766,2.9634414,6.902983,10.8425255,14.782067,18.72161,22.66115,20.560583,18.45611,16.355541,14.251068,12.150499,11.4633255,10.780055,10.096785,9.40961,8.726339,7.0240197,5.3256044,3.6232853,1.9248703,0.22645533,0.23816854,0.25378615,0.26940376,0.28502136,0.30063897,0.8862993,1.4680552,2.0537157,2.639376,3.2250361,3.4671092,3.7091823,3.951255,4.193328,4.4393053,4.521298,4.60329,4.6852827,4.7672753,4.8492675,4.283129,3.7208953,3.154757,2.5886188,2.0263848,1.9287747,1.8311646,1.7335546,1.6359446,1.5383345,3.416352,5.2943697,7.168483,9.0465,10.924518,12.189544,13.45457,14.719597,15.984623,17.24965,13.805966,10.358379,6.914696,3.4710135,0.023426414,1.456342,2.8853533,4.3143644,5.743376,7.1762915,6.969358,6.7663293,6.559396,6.356367,6.1494336,6.606249,7.0630636,7.523783,7.9805984,8.437413,7.8049,7.172387,6.5398736,5.9073606,5.2748475,5.6809053,6.0908675,6.4969254,6.9068875,7.3129454,5.8487945,4.388548,2.9243972,1.4641509,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.6637484,0.8238289,0.9878138,1.1517987,1.3118792,1.2103647,1.1088502,1.0034313,0.9019169,0.80040246,0.80821127,0.8199245,0.8316377,0.8394465,0.8511597,0.9956226,1.1439898,1.2923572,1.4407244,1.5890918,1.53443,1.4836729,1.4290112,1.3782539,1.3235924,1.1361811,0.94876975,0.76135844,0.57394713,0.38653582,0.359205,0.3318742,0.30454338,0.27721256,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,0.12884527,0.19912452,0.26549935,0.3318742,0.39824903,0.3474918,0.29673457,0.24207294,0.19131571,0.13665408,0.1835069,0.23426414,0.28111696,0.3279698,0.37482262,0.42557985,0.48024148,0.5309987,0.58566034,0.63641757,0.77697605,0.91753453,1.0580931,1.1986516,1.33921,1.5227169,1.7062237,1.893635,2.077142,2.260649,2.1083772,1.9561055,1.8038338,1.6515622,1.4992905,1.2415999,0.98000497,0.71841,0.46071947,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,0.26159495,0.26940376,0.27330816,0.27721256,0.28111696,0.28892577,0.30454338,0.3240654,0.339683,0.359205,0.37482262,0.37872702,0.38653582,0.39044023,0.39434463,0.39824903,0.41777104,0.43338865,0.45291066,0.46852827,0.48805028,0.4958591,0.5075723,0.5192855,0.5270943,0.5388075,0.5231899,0.5075723,0.49195468,0.47633708,0.46071947,0.43338865,0.40605783,0.37872702,0.3513962,0.3240654,3.8263142,4.5173936,5.2084727,5.903456,6.5945354,7.289519,7.988407,8.691199,9.393991,10.096785,10.799577,9.924991,9.050405,8.175818,7.3012323,6.426646,5.55206,4.6813784,3.8067923,2.9361105,2.0615244,1.6515622,1.2376955,0.8238289,0.41386664,0.0,0.14055848,0.28502136,0.42557985,0.5700427,0.7106012,0.58566034,0.46071947,0.3357786,0.21083772,0.08589685,0.48414588,0.8784905,1.2728351,1.6671798,2.0615244,2.6276627,3.193801,3.7560349,4.322173,4.8883114,7.4144597,9.940608,12.470661,14.996809,17.526861,19.233086,20.93931,22.649437,24.355661,26.061886,26.02284,25.983797,25.94085,25.901804,25.86276,23.043781,20.228708,17.409729,14.590752,11.775677,13.559989,15.344301,17.128613,18.916828,20.701141,25.17168,29.638317,34.108856,38.5794,43.04994,36.084484,29.115128,22.14577,15.180316,8.210958,10.944039,13.673217,16.402393,19.13157,21.860748,17.975868,14.087084,10.198298,6.3134184,2.4246337,2.8658314,3.3031244,3.7443218,4.185519,4.6267166,6.590631,8.55845,10.526268,12.494087,14.461906,12.041177,9.616543,7.195813,4.7711797,2.35045,1.901444,1.4485333,0.999527,0.5505207,0.10151446,0.42557985,0.74964523,1.0737107,1.4016805,1.7257458,1.6632754,1.6008049,1.5383345,1.475864,1.4133936,2.6706111,3.9317331,5.192855,6.453977,7.7111945,9.573594,11.43209,13.29449,15.152986,17.01148,16.570284,16.129086,15.683984,15.242786,14.801589,12.408191,10.018696,7.629202,5.239708,2.8502135,3.377308,3.9044023,4.4314966,4.958591,5.4856853,5.036679,4.5876727,4.138666,3.6857557,3.2367494,2.8306916,2.4285383,2.0224805,1.6164225,1.2142692,4.755562,8.296855,11.838148,15.383345,18.924637,19.053482,19.186234,19.315079,19.443924,19.576674,17.93292,16.289165,14.645412,13.005564,11.361811,10.61607,9.866425,9.120684,8.371038,7.6252975,7.4495993,7.2739015,7.098203,6.9264097,6.7507114,5.743376,4.73604,3.7287042,2.7213683,1.7140326,3.6740425,5.6379566,7.601871,9.561881,11.525795,10.413041,9.300286,8.187531,7.0747766,5.9620223,4.7711797,3.5764325,2.3855898,1.1908426,0.0,0.14446288,0.28892577,0.43338865,0.58175594,0.7262188,0.58566034,0.44510186,0.30454338,0.1639849,0.023426414,0.12884527,0.23426414,0.339683,0.44510186,0.5505207,0.75745404,0.96438736,1.1713207,1.3782539,1.5890918,1.8663043,2.1435168,2.4207294,2.697942,2.9751544,2.7838387,2.5964274,2.4051118,2.2137961,2.0263848,1.7608855,1.4992905,1.2376955,0.97610056,0.7106012,1.0034313,1.2962615,1.5890918,1.8819219,2.174752,2.3426414,2.5105307,2.67842,2.8463092,3.0141985,2.6471848,2.2840753,1.9170616,1.5539521,1.1869383,1.4797685,1.7725986,2.0654287,2.358259,2.6510892,5.239708,7.8283267,10.42085,13.009468,15.598087,16.191557,16.785025,17.378494,17.971964,18.56153,17.624472,16.683512,15.74255,14.801589,13.860628,11.490656,9.120684,6.7507114,4.380739,2.0107672,2.3114061,2.6081407,2.9048753,3.2016098,3.4983444,3.2211318,2.9439192,2.6667068,2.3894942,2.1122816,1.9404879,1.7686942,1.5969005,1.4212024,1.2494087,3.3812122,5.5091114,7.6409154,9.768814,11.900618,13.333533,14.770353,16.20327,17.640089,19.07691,17.124708,15.176412,13.224211,11.275913,9.323712,7.699481,6.0713453,4.4432096,2.815074,1.1869383,1.9209659,2.6588979,3.3929255,4.126953,4.860981,3.8887846,2.9165885,1.9443923,0.97219616,0.0,0.16008049,0.32016098,0.48024148,0.64032197,0.80040246,1.3626363,1.9248703,2.4871042,3.049338,3.611572,4.4861584,5.35684,6.2314262,7.1021075,7.9766936,10.530173,13.083652,15.641035,18.194515,20.747993,27.162926,33.573956,39.988888,46.399918,52.810944,50.956352,49.10176,47.247173,45.392582,43.53799,40.820526,38.10306,35.385597,32.668133,29.95067,26.026745,22.098917,18.174992,14.251068,10.323239,9.593117,8.859089,8.128965,7.394938,6.66091,6.571109,6.481308,6.3915067,6.3017054,6.211904,6.676528,7.141152,7.605776,8.074304,8.538928,7.363703,6.1884775,5.0132523,3.8380275,2.6628022,3.8965936,5.12648,6.3602715,7.5940623,8.823949,10.416945,12.009941,13.602938,15.195933,16.788929,14.684457,12.583888,10.479416,8.378847,6.2743745,5.02887,3.7794614,2.533957,1.2845483,0.039044023,0.42557985,0.81211567,1.1986516,1.5890918,1.9756275,6.5867267,11.193921,15.80502,20.416119,25.023314,23.664581,22.305851,20.943214,19.584482,18.22575,17.198893,16.172033,15.141272,14.114414,13.087557,10.498938,7.914223,5.3256044,2.736986,0.14836729,0.1717937,0.19522011,0.21864653,0.23816854,0.26159495,0.64032197,1.0190489,1.3938715,1.7725986,2.1513257,2.7565079,3.3655949,3.970777,4.579864,5.1889505,5.169429,5.1460023,5.12648,5.1069584,5.087436,4.677474,4.267512,3.8575494,3.4475873,3.0376248,2.6471848,2.2567444,1.8663043,1.475864,1.0893283,4.1464753,7.2075267,10.268578,13.329629,16.386776,18.284315,20.181856,22.079395,23.976934,25.874474,20.70895,15.539521,10.373997,5.2045684,0.039044023,2.1708477,4.3026514,6.434455,8.566258,10.701966,10.006983,9.311999,8.6131115,7.918128,7.223144,7.4691215,7.7111945,7.9532676,8.19534,8.437413,8.331994,8.226576,8.121157,8.015738,7.914223,7.355894,6.7975645,6.239235,5.6809053,5.12648,4.0996222,3.076669,2.0498111,1.0268579,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,0.8511597,1.0737107,1.3001659,1.5266213,1.7491722,1.6164225,1.4797685,1.3431144,1.2103647,1.0737107,1.0034313,0.92924774,0.8589685,0.78478485,0.7106012,0.8902037,1.0659018,1.2455044,1.4212024,1.6008049,1.5656652,1.5305257,1.4953861,1.4602464,1.4251068,1.2142692,0.999527,0.78868926,0.57394713,0.3631094,0.339683,0.31625658,0.29673457,0.27330816,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,0.10932326,0.15227169,0.19912452,0.24207294,0.28892577,0.25378615,0.21864653,0.1835069,0.14836729,0.113227665,0.14055848,0.1678893,0.19522011,0.22255093,0.24988174,0.30844778,0.3709182,0.42948425,0.48805028,0.5505207,0.7106012,0.8706817,1.0307622,1.1908426,1.3509232,1.6281357,1.9053483,2.182561,2.4597735,2.736986,2.5886188,2.4441557,2.2957885,2.1474214,1.999054,1.6359446,1.2689307,0.9058213,0.5388075,0.1756981,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24597734,0.25378615,0.26159495,0.26940376,0.27330816,0.29673457,0.31625658,0.3357786,0.3553006,0.37482262,0.38263142,0.39044023,0.39824903,0.40605783,0.41386664,0.42167544,0.42557985,0.43338865,0.44119745,0.44900626,0.45291066,0.45681506,0.45681506,0.46071947,0.46071947,0.45291066,0.44119745,0.43338865,0.42167544,0.41386664,0.39044023,0.3670138,0.3435874,0.3240654,0.30063897,2.475391,3.8770714,5.278752,6.6843367,8.086017,9.487698,10.206107,10.928422,11.6468315,12.369146,13.087557,11.888905,10.686349,9.487698,8.289046,7.08649,6.2197127,5.3529353,4.4861584,3.619381,2.7486992,2.1981785,1.6515622,1.1010414,0.5505207,0.0,0.19131571,0.37872702,0.5700427,0.76135844,0.94876975,0.77307165,0.60127795,0.42557985,0.24988174,0.07418364,0.43338865,0.79649806,1.1557031,1.5149081,1.8741131,2.2216048,2.5651922,2.9087796,3.2562714,3.5998588,6.8092775,10.0147915,13.224211,16.429726,19.639143,22.161386,24.683632,27.205875,29.728119,32.250362,31.55538,30.860395,30.165411,29.470428,28.775444,24.660204,20.544964,16.429726,12.314485,8.1992445,11.705398,15.211552,18.7138,22.219954,25.726107,31.758408,37.794613,43.83082,49.867027,55.899326,45.634655,35.36998,25.105307,14.840633,4.575959,8.066495,11.553126,15.043662,18.534197,22.024733,18.22575,14.426766,10.6238785,6.824895,3.0259118,3.631094,4.240181,4.8492675,5.45445,6.0635366,6.329036,6.590631,6.8561306,7.1216297,7.387129,6.2079997,5.02887,3.8458362,2.6667068,1.4875772,1.2142692,0.93705654,0.6637484,0.38653582,0.113227665,0.3240654,0.5388075,0.74964523,0.96438736,1.175225,1.1127546,1.0502841,0.9878138,0.92534333,0.8628729,2.7057507,4.548629,6.3915067,8.234385,10.073358,11.217348,12.361338,13.501423,14.645412,15.789403,15.847969,15.906535,15.969006,16.02757,16.086138,13.181262,10.272482,7.363703,4.4588275,1.5500476,2.1435168,2.7408905,3.3343596,3.9317331,4.5252023,4.349504,4.173806,3.998108,3.8263142,3.6506162,3.096191,2.5456703,1.9912452,1.4407244,0.8862993,4.2011366,7.5159745,10.8308115,14.145649,17.464392,16.48829,15.516094,14.543899,13.571702,12.599506,11.39695,10.194394,8.991838,7.7892823,6.5867267,6.083059,5.579391,5.0718184,4.5681505,4.0605783,4.650143,5.2358036,5.825368,6.4110284,7.000593,5.891743,4.7789884,3.6701381,2.5612879,1.4485333,3.8380275,6.223617,8.6131115,10.998701,13.388195,12.037272,10.686349,9.339331,7.988407,6.6374836,5.309987,3.9824903,2.6549935,1.3274968,0.0,0.07418364,0.14446288,0.21864653,0.28892577,0.3631094,0.29283017,0.22255093,0.15227169,0.08199245,0.011713207,0.15227169,0.29283017,0.43338865,0.57394713,0.7106012,0.94876975,1.183034,1.4172981,1.6515622,1.8858263,2.2957885,2.7018464,3.1118085,3.5178664,3.9239242,3.6662338,3.408543,3.1508527,2.893162,2.639376,2.2137961,1.7882162,1.3626363,0.93705654,0.5114767,0.9917182,1.4680552,1.9443923,2.4207294,2.900971,2.9634414,3.0298162,3.096191,3.1586614,3.2250361,2.7057507,2.1864653,1.6632754,1.1439898,0.62470436,0.9136301,1.2064602,1.4953861,1.7843118,2.0732377,4.181615,6.289992,8.398369,10.506746,12.611219,15.039758,17.468296,19.896833,22.321468,24.750006,22.192623,19.635239,17.077856,14.520472,11.963089,9.991365,8.015738,6.044015,4.0722914,2.1005683,2.541766,2.9868677,3.4280653,3.8692627,4.3143644,3.7052777,3.096191,2.4910088,1.8819219,1.2767396,1.2337911,1.1908426,1.1478943,1.1049459,1.0619974,2.7916477,4.5173936,6.2431393,7.9727893,9.698535,11.767868,13.833297,15.902631,17.971964,20.037392,18.38583,16.738173,15.086611,13.438952,11.787391,9.718058,7.648724,5.579391,3.506153,1.43682,2.3816853,3.3226464,4.263607,5.2084727,6.1494336,4.919547,3.68966,2.4597735,1.2298868,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,0.96438736,1.5266213,2.0888553,2.6510892,3.213323,3.3812122,3.5491016,3.7130866,3.8809757,4.0488653,6.578918,9.105066,11.631214,14.161267,16.687416,25.074072,33.460728,41.851288,50.237946,58.6246,56.473274,54.32195,52.166718,50.015392,47.864067,45.060707,42.257347,39.453983,36.650623,33.851166,29.58756,25.323954,21.06425,16.800642,12.537036,11.576552,10.61607,9.655587,8.699008,7.7385254,7.480835,7.223144,6.9654536,6.707763,6.4500723,7.1216297,7.7892823,8.460839,9.128492,9.80005,8.538928,7.2739015,6.012779,4.7516575,3.4866312,4.9351645,6.3836975,7.8283267,9.276859,10.725393,11.478943,12.228588,12.982138,13.735687,14.489237,12.228588,9.971844,7.715099,5.4583545,3.2016098,2.5690966,1.9404879,1.3118792,0.679366,0.05075723,0.23816854,0.42557985,0.61299115,0.80040246,0.9878138,6.266566,11.549222,16.827974,22.106726,27.389381,26.768581,26.151686,25.53479,24.917894,24.300999,22.930555,21.56011,20.189665,18.81922,17.448774,13.973856,10.498938,7.0240197,3.5491016,0.07418364,0.10541886,0.13665408,0.1639849,0.19522011,0.22645533,0.39434463,0.5661383,0.7340276,0.9058213,1.0737107,2.0459068,3.018103,3.9942036,4.9663997,5.938596,5.813655,5.6926184,5.571582,5.446641,5.3256044,5.0718184,4.814128,4.560342,4.3065557,4.0488653,3.3655949,2.6862288,2.0029583,1.319688,0.63641757,4.8805027,9.120684,13.364769,17.608854,21.849035,24.379087,26.90914,29.439194,31.969246,34.4993,27.608028,20.720663,13.829392,6.9381227,0.05075723,2.8853533,5.7199492,8.554545,11.389141,14.223738,13.040704,11.8537655,10.670732,9.483793,8.300759,8.32809,8.355421,8.382751,8.410083,8.437413,8.859089,9.280765,9.706344,10.128019,10.549695,9.026978,7.504261,5.9815445,4.4588275,2.9361105,2.35045,1.7608855,1.175225,0.58566034,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14836729,0.30063897,0.44900626,0.60127795,0.74964523,1.038571,1.3235924,1.6125181,1.901444,2.1864653,2.018576,1.8506867,1.6867018,1.5188124,1.3509232,1.1947471,1.038571,0.8862993,0.7301232,0.57394713,0.78088045,0.9917182,1.1986516,1.4055848,1.6125181,1.5969005,1.5773785,1.5617609,1.542239,1.5266213,1.2884527,1.0502841,0.81211567,0.57394713,0.3357786,0.32016098,0.30063897,0.28502136,0.26940376,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,0.08589685,0.10932326,0.12884527,0.15227169,0.1756981,0.15617609,0.14055848,0.12103647,0.10541886,0.08589685,0.093705654,0.10151446,0.10932326,0.11713207,0.12494087,0.19131571,0.26159495,0.3279698,0.39434463,0.46071947,0.6442264,0.8238289,1.0034313,1.183034,1.3626363,1.7335546,2.1044729,2.4714866,2.8424048,3.213323,3.06886,2.9283018,2.7838387,2.6432803,2.4988174,2.0302892,1.5617609,1.0893283,0.62079996,0.14836729,0.1639849,0.1756981,0.18741131,0.19912452,0.21083772,0.22255093,0.23426414,0.24207294,0.25378615,0.26159495,0.28502136,0.30844778,0.3318742,0.3513962,0.37482262,0.38653582,0.39434463,0.40605783,0.41386664,0.42557985,0.42167544,0.42167544,0.41777104,0.41386664,0.41386664,0.40605783,0.40215343,0.39824903,0.39434463,0.38653582,0.38263142,0.37872702,0.3709182,0.3670138,0.3631094,0.3435874,0.3279698,0.30844778,0.29283017,0.27330816,1.1244678,3.2367494,5.349031,7.461313,9.573594,11.685876,12.423808,13.16174,13.899672,14.637604,15.375536,13.848915,12.326198,10.799577,9.276859,7.7502384,6.8873653,6.0244927,5.1616197,4.298747,3.435874,2.7486992,2.0615244,1.3743496,0.6871748,0.0,0.23816854,0.47633708,0.7106012,0.94876975,1.1869383,0.96438736,0.737932,0.5114767,0.28892577,0.062470436,0.38653582,0.7106012,1.038571,1.3626363,1.6867018,1.8116426,1.9365835,2.0615244,2.1864653,2.3114061,6.2001905,10.088976,13.973856,17.86264,21.751425,25.085785,28.42405,31.762312,35.100574,38.43884,37.087917,35.736996,34.38607,33.03905,31.68813,26.276627,20.861221,15.449719,10.0382185,4.6267166,9.850807,15.074897,20.298986,25.526981,30.751072,38.349037,45.95091,53.548878,61.15075,68.74872,55.188725,41.624832,28.06094,14.50095,0.93705654,5.1889505,9.43694,13.688834,17.936825,22.188719,18.475632,14.762545,11.0494585,7.336372,3.6232853,4.4002614,5.173333,5.950309,6.7233806,7.5003567,6.0635366,4.6267166,3.1859922,1.7491722,0.31235218,0.37482262,0.43729305,0.4997635,0.5622339,0.62470436,0.5231899,0.42557985,0.3240654,0.22645533,0.12494087,0.22645533,0.3240654,0.42557985,0.5231899,0.62470436,0.5622339,0.4997635,0.43729305,0.37482262,0.31235218,2.736986,5.1616197,7.5862536,10.010887,12.439425,12.861101,13.286681,13.712261,14.13784,14.56342,15.125654,15.687888,16.250122,16.812357,17.37459,13.950429,10.526268,7.098203,3.6740425,0.24988174,0.9136301,1.5734742,2.2372224,2.900971,3.5608149,3.6623292,3.7638438,3.8614538,3.9629683,4.0605783,3.3616903,2.6628022,1.9639144,1.261122,0.5622339,3.6506162,6.7389984,9.823476,12.911859,16.00024,13.923099,11.849861,9.776623,7.699481,5.6262436,4.860981,4.0996222,3.338264,2.5769055,1.8116426,1.5500476,1.2884527,1.0268579,0.76135844,0.4997635,1.8506867,3.2016098,4.548629,5.899552,7.250475,6.036206,4.825841,3.611572,2.4012074,1.1869383,3.998108,6.813182,9.6243515,12.439425,15.250595,13.661504,12.076316,10.487225,8.898132,7.3129454,5.8487945,4.388548,2.9243972,1.4641509,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1756981,0.3513962,0.5231899,0.698888,0.8745861,1.1361811,1.4016805,1.6632754,1.9248703,2.1864653,2.7252727,3.2640803,3.7989833,4.337791,4.8765984,4.548629,4.224563,3.900498,3.5764325,3.2484627,2.6628022,2.0732377,1.4875772,0.9019169,0.31235218,0.97610056,1.6359446,2.2996929,2.9634414,3.6232853,3.5881457,3.5491016,3.513962,3.474918,3.435874,2.7643168,2.0888553,1.4133936,0.737932,0.062470436,0.3513962,0.63641757,0.92534333,1.2142692,1.4992905,3.1235218,4.7516575,6.375889,8.00012,9.6243515,13.887959,18.151566,22.411268,26.674877,30.938484,26.760773,22.586967,18.41316,14.239355,10.061645,8.488171,6.910792,5.337318,3.7638438,2.1864653,2.77603,3.3616903,3.951255,4.5369153,5.12648,4.1894236,3.2484627,2.3114061,1.3743496,0.43729305,0.5231899,0.61299115,0.698888,0.78868926,0.8745861,2.1981785,3.5256753,4.8492675,6.1767645,7.5003567,10.198298,12.900145,15.601992,18.299932,21.00178,19.650856,18.299932,16.94901,15.598087,14.251068,11.736633,9.226103,6.7116675,4.2011366,1.6867018,2.8385005,3.9863946,5.138193,6.2860875,7.437886,5.950309,4.462732,2.9751544,1.4875772,0.0,0.0,0.0,0.0,0.0,0.0,0.5622339,1.1244678,1.6867018,2.2489357,2.8111696,2.2762666,1.737459,1.1986516,0.6637484,0.12494087,2.6237583,5.12648,7.6252975,10.124115,12.626837,22.98912,33.351402,43.713688,54.07597,64.438255,61.98629,59.53823,57.086266,54.638206,52.18624,49.300888,46.41163,43.526276,40.63702,37.751667,33.148376,28.548988,23.949604,19.350218,14.750832,13.563893,12.376955,11.186112,9.999174,8.812236,8.386656,7.9610763,7.5394006,7.113821,6.688241,7.562827,8.437413,9.311999,10.186585,11.061172,9.714153,8.36323,7.012306,5.661383,4.3143644,5.9737353,7.6370106,9.300286,10.963562,12.626837,12.537036,12.4511385,12.361338,12.27544,12.185639,9.776623,7.363703,4.950782,2.5378613,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,5.950309,11.900618,17.850927,23.801235,29.751545,29.876486,30.001427,30.126368,30.251308,30.37625,28.662216,26.948185,25.238056,23.524023,21.813896,17.448774,13.087557,8.726339,4.3612175,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,1.33921,2.6745155,4.0137253,5.349031,6.688241,6.461786,6.239235,6.012779,5.786324,5.563773,5.462259,5.3607445,5.263134,5.1616197,5.0640097,4.087909,3.1118085,2.135708,1.1635119,0.18741131,5.6145306,11.037745,16.46096,21.888079,27.311295,30.47386,33.636425,36.798992,39.961555,43.124123,34.511013,25.901804,17.288692,8.675582,0.062470436,3.5998588,7.137247,10.674636,14.212025,17.749413,16.074425,14.399435,12.724447,11.0494585,9.37447,9.187058,8.999647,8.812236,8.624825,8.437413,9.386183,10.338858,11.287627,12.236397,13.189071,10.698062,8.210958,5.7238536,3.2367494,0.74964523,0.60127795,0.44900626,0.30063897,0.14836729,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1756981,0.3513962,0.5231899,0.698888,0.8745861,1.2259823,1.5734742,1.9248703,2.2762666,2.6237583,2.4246337,2.2255092,2.0263848,1.8233559,1.6242313,1.3860629,1.1517987,0.9136301,0.6754616,0.43729305,0.6754616,0.9136301,1.1517987,1.3860629,1.6242313,1.6242313,1.6242313,1.6242313,1.6242313,1.6242313,1.3626363,1.1010414,0.8355421,0.57394713,0.31235218,0.30063897,0.28892577,0.27330816,0.26159495,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.57394713,0.77697605,0.97610056,1.175225,1.3743496,1.8389735,2.2996929,2.7643168,3.2250361,3.6857557,3.5491016,3.4124475,3.2757936,3.1391394,2.998581,2.4246337,1.8506867,1.2767396,0.698888,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,0.27330816,0.30063897,0.3240654,0.3513962,0.37482262,0.38653582,0.39824903,0.41386664,0.42557985,0.43729305,0.42557985,0.41386664,0.39824903,0.38653582,0.37482262,0.3631094,0.3513962,0.3357786,0.3240654,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.30063897,0.28892577,0.27330816,0.26159495,0.24988174,7.250475,8.097731,8.944985,9.792241,10.639496,11.486752,11.799104,12.107552,12.415999,12.728352,13.036799,11.795199,10.553599,9.308095,8.066495,6.824895,6.0908675,5.35684,4.618908,3.8848803,3.1508527,2.5534792,1.9561055,1.358732,0.76135844,0.1639849,0.37872702,0.59737355,0.8160201,1.0307622,1.2494087,1.0151446,0.78088045,0.5466163,0.30844778,0.07418364,0.3709182,0.6715572,0.96829176,1.2650263,1.5617609,1.9717231,2.377781,2.7838387,3.193801,3.5998588,6.7780423,9.96013,13.138313,16.320402,19.498585,23.37956,27.260536,31.141512,35.018585,38.89956,37.876606,36.849747,35.826794,34.79994,33.77308,29.16198,24.55088,19.935879,15.324779,10.71368,14.989,19.260416,23.535736,27.811058,32.086376,36.935646,41.78882,46.638084,51.487354,56.33662,45.396484,34.45635,23.516214,12.576079,1.6359446,5.1303844,8.62092,12.11536,15.605896,19.100336,15.918248,12.73616,9.554072,6.36808,3.1859922,3.7482262,4.3143644,4.8765984,5.4388323,6.001066,4.9820175,3.9668727,2.9478238,1.9287747,0.9136301,0.8316377,0.74574083,0.6637484,0.58175594,0.4997635,0.44510186,0.39044023,0.3357786,0.28111696,0.22645533,0.31625658,0.40996224,0.5036679,0.59346914,0.6871748,0.8862993,1.0815194,1.2806439,1.475864,1.6749885,3.4671092,5.2592297,7.0513506,8.843472,10.6355915,11.111929,11.584361,12.056794,12.529227,13.001659,13.6693125,14.34087,15.008522,15.680079,16.351637,13.153932,9.96013,6.7663293,3.5686235,0.37482262,0.8980125,1.4212024,1.9443923,2.463678,2.9868677,3.541293,4.0918136,4.646239,5.196759,5.7511845,5.083532,4.4197836,3.7560349,3.0883822,2.4246337,4.853172,7.28171,9.706344,12.134882,14.56342,13.528754,12.497992,11.4633255,10.432563,9.4018,8.695104,7.988407,7.2856145,6.578918,5.8761253,4.9078336,3.9395418,2.97125,2.0068626,1.038571,2.069333,3.096191,4.126953,5.1577153,6.1884775,5.298274,4.4119744,3.5256753,2.639376,1.7491722,3.8614538,5.9737353,8.086017,10.198298,12.314485,11.029937,9.749292,8.464745,7.1841,5.899552,4.747753,3.5959544,2.4441557,1.2884527,0.13665408,0.12103647,0.10151446,0.08589685,0.06637484,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.14055848,0.28502136,0.42557985,0.5700427,0.7106012,0.92143893,1.1283722,1.3353056,1.542239,1.7491722,2.1864653,2.6237583,3.0610514,3.4983444,3.9356375,3.6701381,3.4007344,3.135235,2.8658314,2.6003318,2.1318035,1.6632754,1.1986516,0.7301232,0.26159495,0.78868926,1.3157835,1.8467822,2.3738766,2.900971,2.87364,2.8463092,2.8189783,2.7916477,2.7643168,2.3621633,1.9639144,1.5617609,1.1635119,0.76135844,0.8589685,0.95657855,1.0541886,1.1517987,1.2494087,2.97125,4.689187,6.4110284,8.128965,9.850807,13.423335,16.995863,20.568392,24.140919,27.713448,23.891037,20.068628,16.246218,12.423808,8.601398,7.4417906,6.278279,5.1186714,3.959064,2.7994564,3.310933,3.8185053,4.3299823,4.841459,5.349031,4.349504,3.349977,2.35045,1.3509232,0.3513962,0.48414588,0.62079996,0.75354964,0.8902037,1.0268579,2.5183394,4.009821,5.5013027,6.996689,8.488171,10.373997,12.263727,14.149553,16.039284,17.92511,16.769407,15.6098,14.454097,13.29449,12.138786,10.518459,8.898132,7.277806,5.657479,4.037152,4.9546866,5.872221,6.7897553,7.70729,8.624825,6.899079,5.173333,3.4514916,1.7257458,0.0,0.23426414,0.46462387,0.698888,0.92924774,1.1635119,1.4290112,1.698415,1.9639144,2.233318,2.4988174,2.0420024,1.5851873,1.1283722,0.6715572,0.21083772,3.2640803,6.3173227,9.370565,12.423808,15.473146,22.977407,30.47386,37.974216,45.47457,52.97493,52.533733,52.08863,51.647434,51.206234,50.761135,48.465343,46.165653,43.869865,41.574074,39.274384,34.401688,29.528994,24.6563,19.783606,14.9109125,14.176885,13.442857,12.708829,11.970898,11.23687,10.979179,10.721489,10.4637985,10.206107,9.948417,10.393518,10.834716,11.275913,11.721016,12.162213,11.510178,10.858143,10.206107,9.554072,8.898132,9.823476,10.748819,11.674163,12.599506,13.524849,14.606369,15.683984,16.765503,17.843119,18.924637,15.160794,11.39695,7.629202,3.8653584,0.10151446,0.9136301,1.7257458,2.5378613,3.349977,4.1620927,3.8419318,3.521771,3.2016098,2.8814487,2.5612879,6.942027,11.322766,15.7035055,20.084246,24.46108,25.456703,26.448421,27.44014,28.431858,29.423576,27.084839,24.746101,22.40346,20.064724,17.725986,14.219833,10.71368,7.211431,3.7052777,0.19912452,0.29673457,0.39044023,0.48414588,0.58175594,0.6754616,0.58175594,0.48414588,0.39044023,0.29673457,0.19912452,1.4133936,2.631567,3.8458362,5.0601053,6.2743745,6.1611466,6.0518236,5.938596,5.825368,5.7121406,5.7121406,5.7121406,5.7121406,5.7121406,5.7121406,4.618908,3.5256753,2.436347,1.3431144,0.24988174,4.6423345,9.034787,13.427239,17.819693,22.212145,24.72658,27.241014,29.759354,32.27379,34.788223,27.842293,20.89636,13.950429,7.008402,0.062470436,3.1586614,6.250948,9.347139,12.44333,15.535617,14.208119,12.880623,11.553126,10.22563,8.898132,8.85128,8.804427,8.757574,8.710721,8.663869,9.339331,10.018696,10.694158,11.373524,12.0489855,9.839094,7.629202,5.4193106,3.2094188,0.999527,0.8394465,0.679366,0.5192855,0.359205,0.19912452,0.1796025,0.16008049,0.14055848,0.12103647,0.10151446,0.41386664,0.7262188,1.038571,1.3509232,1.6632754,1.3314011,0.9956226,0.6637484,0.3318742,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14055848,0.28111696,0.42167544,0.5583295,0.698888,1.0112402,1.3235924,1.6359446,1.9482968,2.260649,2.1396124,2.018576,1.893635,1.7725986,1.6515622,1.3938715,1.1361811,0.8784905,0.62079996,0.3631094,0.57785153,0.79259366,1.0073358,1.2220778,1.43682,1.8272603,2.2177005,2.6081407,2.998581,3.3890212,2.8072653,2.2294137,1.6476578,1.0659018,0.48805028,0.42948425,0.3709182,0.31625658,0.25769055,0.19912452,0.1717937,0.14446288,0.11713207,0.08980125,0.062470436,0.13665408,0.20693332,0.28111696,0.3513962,0.42557985,0.40215343,0.37872702,0.359205,0.3357786,0.31235218,0.28892577,0.26159495,0.23816854,0.21083772,0.18741131,0.28892577,0.39434463,0.4958591,0.59737355,0.698888,1.0541886,1.4094892,1.7647898,2.1200905,2.475391,2.7135596,2.9556324,3.193801,3.435874,3.6740425,3.5842414,3.4905357,3.39683,3.3031244,3.213323,2.7526035,2.2918842,1.8311646,1.3743496,0.9136301,0.78478485,0.6559396,0.5309987,0.40215343,0.27330816,0.3279698,0.37872702,0.43338865,0.48414588,0.5388075,0.5192855,0.5036679,0.48414588,0.46852827,0.44900626,0.45681506,0.46462387,0.47243267,0.48024148,0.48805028,0.46071947,0.43729305,0.41386664,0.38653582,0.3631094,0.3513962,0.3357786,0.3240654,0.31235218,0.30063897,0.30063897,0.30063897,0.30063897,0.30063897,0.30063897,0.28892577,0.27330816,0.26159495,0.24988174,0.23816854,13.376482,12.958711,12.54094,12.123169,11.705398,11.287627,11.170495,11.053363,10.936231,10.819098,10.698062,9.741484,8.781001,7.8205175,6.860035,5.899552,5.2943697,4.6852827,4.0761957,3.4710135,2.8619268,2.3543546,1.8467822,1.33921,0.8316377,0.3240654,0.5231899,0.71841,0.91753453,1.116659,1.3118792,1.0659018,0.8238289,0.57785153,0.3318742,0.08589685,0.359205,0.62860876,0.8980125,1.1674163,1.43682,2.1278992,2.8189783,3.506153,4.1972322,4.8883114,7.3597984,9.8312845,12.306676,14.778163,17.24965,21.673336,26.09312,30.516808,34.940495,39.364185,38.661392,37.9625,37.263615,36.56082,35.861935,32.05124,28.236637,24.425941,20.61134,16.800642,20.12329,23.44984,26.77639,30.099037,33.425587,35.526157,37.626724,39.72339,41.823956,43.924526,35.608147,27.29177,18.97149,10.655114,2.338737,5.0718184,7.8088045,10.541886,13.2788725,16.011953,13.360865,10.705871,8.054782,5.4036927,2.7486992,3.1000953,3.4514916,3.7989833,4.1503797,4.5017757,3.9044023,3.3031244,2.7057507,2.1083772,1.5110037,1.2845483,1.0580931,0.8316377,0.60127795,0.37482262,0.3631094,0.3553006,0.3435874,0.3357786,0.3240654,0.40996224,0.4958591,0.58175594,0.6637484,0.74964523,1.2064602,1.6632754,2.1239948,2.5808098,3.0376248,4.1972322,5.35684,6.5164475,7.676055,8.835662,9.358852,9.878138,10.397423,10.916709,11.435994,12.216875,12.993851,13.770826,14.547803,15.324779,12.361338,9.393991,6.4305506,3.4632049,0.4997635,0.8823949,1.2650263,1.6476578,2.0302892,2.4129205,3.416352,4.423688,5.4271193,6.434455,7.437886,6.8092775,6.1767645,5.548156,4.9156423,4.2870336,6.055728,7.8205175,9.589212,11.357906,13.1266,13.134409,13.146122,13.153932,13.165645,13.173453,12.529227,11.881096,11.232965,10.584834,9.936704,8.265619,6.590631,4.919547,3.2484627,1.5734742,2.2840753,2.9946766,3.7052777,4.415879,5.12648,4.564246,3.998108,3.435874,2.87364,2.3114061,3.7247996,5.138193,6.551587,7.9610763,9.37447,8.398369,7.4183645,6.4422636,5.466163,4.4861584,3.6467118,2.803361,1.9600099,1.116659,0.27330816,0.23816854,0.20693332,0.1717937,0.13665408,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.10932326,0.21864653,0.3318742,0.44119745,0.5505207,0.7027924,0.8550641,1.0073358,1.1596074,1.3118792,1.6515622,1.9873407,2.3231194,2.6628022,2.998581,2.7916477,2.5808098,2.3699722,2.1591344,1.9482968,1.6008049,1.2533131,0.9058213,0.5583295,0.21083772,0.60518235,0.9956226,1.3899672,1.7843118,2.174752,2.1591344,2.1396124,2.1239948,2.1044729,2.0888553,1.9639144,1.8389735,1.7140326,1.5890918,1.4641509,1.3704453,1.2767396,1.1869383,1.0932326,0.999527,2.815074,4.630621,6.446168,8.261715,10.073358,12.958711,15.84016,18.72161,21.606962,24.48841,21.017397,17.546383,14.079274,10.608261,7.137247,6.3915067,5.645766,4.903929,4.1581883,3.4124475,3.8458362,4.279225,4.7087092,5.142098,5.575486,4.513489,3.4514916,2.3855898,1.3235924,0.26159495,0.44510186,0.62860876,0.80821127,0.9917182,1.175225,2.8345962,4.493967,6.153338,7.816613,9.475985,10.549695,11.623405,12.70102,13.774731,14.848442,13.884054,12.919667,11.955279,10.990892,10.0265045,9.296382,8.570163,7.843944,7.113821,6.387602,7.0708723,7.758047,8.441318,9.128492,9.811763,7.8517528,5.8878384,3.9239242,1.9639144,0.0,0.46462387,0.92924774,1.3938715,1.8584955,2.3231194,2.2957885,2.2684577,2.241127,2.2137961,2.1864653,1.8116426,1.4329157,1.0541886,0.679366,0.30063897,3.9044023,7.5081654,11.115833,14.719597,18.32336,22.96179,27.60022,32.23865,36.873177,41.511604,43.07727,44.642937,46.2086,47.774265,49.336025,47.629803,45.92358,44.21345,42.50723,40.801003,35.655003,30.508999,25.362997,20.2209,15.074897,14.79378,14.508759,14.227642,13.946525,13.661504,13.571702,13.481901,13.392099,13.302299,13.212498,13.224211,13.232019,13.243732,13.251541,13.263254,13.306203,13.353056,13.396004,13.442857,13.4858055,13.673217,13.860628,14.051944,14.239355,14.426766,16.671797,18.920732,21.165764,23.4147,25.663635,20.544964,15.426293,10.311526,5.192855,0.07418364,1.7140326,3.349977,4.985922,6.6257706,8.261715,7.633106,7.008402,6.379793,5.7511845,5.12648,7.9337454,10.744915,13.556085,16.36335,19.174519,21.036919,22.895414,24.75391,26.61631,28.474806,25.50746,22.540113,19.57277,16.605423,13.638077,10.990892,8.343708,5.6965227,3.049338,0.39824903,0.5544251,0.7066968,0.8589685,1.0112402,1.1635119,1.0112402,0.8589685,0.7066968,0.5544251,0.39824903,1.4914817,2.5847144,3.677947,4.7711797,5.8644123,5.8644123,5.8644123,5.8644123,5.8644123,5.8644123,5.9620223,6.0635366,6.1611466,6.262661,6.364176,5.153811,3.9434462,2.7330816,1.5227169,0.31235218,3.6740425,7.0318284,10.393518,13.751305,17.112995,18.9793,20.845604,22.715813,24.582117,26.448421,21.173573,15.894821,10.61607,5.3412223,0.062470436,2.7135596,5.368553,8.019642,10.670732,13.325725,12.34572,11.365715,10.38571,9.405705,8.4257,8.519405,8.609207,8.702912,8.796618,8.886419,9.292478,9.698535,10.100689,10.506746,10.912805,8.980125,7.0474463,5.114767,3.182088,1.2494087,1.0815194,0.9097257,0.7418364,0.5700427,0.39824903,0.359205,0.32016098,0.28111696,0.23816854,0.19912452,0.8238289,1.4485333,2.0732377,2.7018464,3.3265507,2.6588979,1.9951496,1.3314011,0.6637484,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10541886,0.21083772,0.31625658,0.42167544,0.5231899,0.80040246,1.0737107,1.3509232,1.6242313,1.901444,1.8545911,1.8116426,1.7647898,1.7218413,1.6749885,1.397776,1.1205635,0.8433509,0.5661383,0.28892577,0.48024148,0.6715572,0.8667773,1.0580931,1.2494087,2.0302892,2.8111696,3.5881457,4.369026,5.1499066,4.251894,3.3538816,2.455869,1.5617609,0.6637484,0.5583295,0.45681506,0.3553006,0.25378615,0.14836729,0.13274968,0.113227665,0.09761006,0.078088045,0.062470436,0.20693332,0.3513962,0.4958591,0.6442264,0.78868926,0.7418364,0.698888,0.6520352,0.60908675,0.5622339,0.5231899,0.48805028,0.44900626,0.41386664,0.37482262,0.5036679,0.63641757,0.76526284,0.8941081,1.0268579,1.53443,2.0459068,2.5534792,3.0649557,3.5764325,3.59205,3.611572,3.6271896,3.6467118,3.6623292,3.6154766,3.5686235,3.521771,3.4710135,3.4241607,3.0805733,2.7330816,2.3894942,2.0459068,1.698415,1.4329157,1.1635119,0.8980125,0.62860876,0.3631094,0.45681506,0.5466163,0.64032197,0.7340276,0.8238289,0.76526284,0.7066968,0.6442264,0.58566034,0.5231899,0.5270943,0.5309987,0.5309987,0.5349031,0.5388075,0.4997635,0.46071947,0.42557985,0.38653582,0.3513962,0.3357786,0.3240654,0.31235218,0.30063897,0.28892577,0.28892577,0.28892577,0.28892577,0.28892577,0.28892577,0.27330816,0.26159495,0.24988174,0.23816854,0.22645533,19.498585,17.815788,16.136894,14.454097,12.771299,11.088503,10.541886,9.999174,9.452558,8.905942,8.36323,7.6838636,7.008402,6.329036,5.6535745,4.9742084,4.493967,4.0137253,3.533484,3.0532427,2.5769055,2.1591344,1.7413634,1.3235924,0.9058213,0.48805028,0.6637484,0.8433509,1.0190489,1.1986516,1.3743496,1.1205635,0.8667773,0.60908675,0.3553006,0.10151446,0.3435874,0.58566034,0.8277333,1.0698062,1.3118792,2.2840753,3.2562714,4.2284675,5.2006636,6.1767645,7.941554,9.706344,11.471134,13.235924,15.000713,19.96321,24.92961,29.896008,34.858505,39.8249,39.45008,39.075256,38.700436,38.32561,37.95079,34.936592,31.926298,28.912098,25.901804,22.887606,25.261482,27.639263,30.01314,32.387016,34.760895,34.112762,33.460728,32.812595,32.16056,31.51243,25.815908,20.12329,14.426766,8.734148,3.0376248,5.0132523,6.9927845,8.968412,10.947944,12.923572,10.803481,8.679486,6.5554914,4.435401,2.3114061,2.4480603,2.5886188,2.7252727,2.8619268,2.998581,2.822883,2.6432803,2.4675822,2.2918842,2.1122816,1.7413634,1.3665408,0.9956226,0.62079996,0.24988174,0.28502136,0.32016098,0.3553006,0.39044023,0.42557985,0.5036679,0.58175594,0.6559396,0.7340276,0.81211567,1.5305257,2.2489357,2.9634414,3.6818514,4.4002614,4.927356,5.45445,5.9815445,6.5086384,7.0357327,7.605776,8.171914,8.738052,9.308095,9.874233,10.760532,11.6468315,12.529227,13.415526,14.301826,11.564839,8.831758,6.094772,3.3616903,0.62470436,0.8667773,1.1088502,1.3509232,1.5969005,1.8389735,3.2953155,4.7516575,6.211904,7.6682463,9.124588,8.531119,7.9337454,7.3402762,6.746807,6.1494336,7.2582836,8.36323,9.47208,10.58093,11.685876,12.740065,13.794253,14.844538,15.8987255,16.94901,16.359446,15.76988,15.180316,14.590752,14.001186,11.623405,9.245625,6.8678436,4.4900627,2.1122816,2.5027218,2.893162,3.2836022,3.6740425,4.0605783,3.8263142,3.5881457,3.349977,3.1118085,2.87364,3.5881457,4.298747,5.0132523,5.7238536,6.4383593,5.7668023,5.0913405,4.4197836,3.7482262,3.076669,2.541766,2.0107672,1.475864,0.94486535,0.41386664,0.359205,0.30844778,0.25378615,0.20302892,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.078088045,0.15617609,0.23426414,0.30844778,0.38653582,0.48414588,0.58175594,0.679366,0.77697605,0.8745861,1.1127546,1.3509232,1.5890918,1.8233559,2.0615244,1.9092526,1.756981,1.6047094,1.4524376,1.3001659,1.0737107,0.8433509,0.61689556,0.39044023,0.1639849,0.42167544,0.679366,0.93315214,1.1908426,1.4485333,1.4407244,1.43682,1.4290112,1.4212024,1.4133936,1.5617609,1.7140326,1.8623998,2.0107672,2.1630387,1.8819219,1.5969005,1.3157835,1.0307622,0.74964523,2.6588979,4.5681505,6.481308,8.39056,10.299813,12.494087,14.684457,16.87873,19.069101,21.263374,18.143757,15.028045,11.908427,8.792714,5.6730967,5.3451266,5.0132523,4.6852827,4.3534083,4.025439,4.380739,4.73604,5.0913405,5.446641,5.801942,4.6735697,3.5491016,2.4246337,1.3001659,0.1756981,0.40605783,0.63641757,0.8667773,1.0932326,1.3235924,3.1508527,4.9781127,6.8092775,8.636538,10.4637985,10.725393,10.986988,11.248583,11.514082,11.775677,11.002605,10.229534,9.456462,8.683391,7.914223,8.078208,8.242193,8.406178,8.574067,8.738052,9.190963,9.643873,10.096785,10.545791,10.998701,8.800523,6.5984397,4.4002614,2.1981785,0.0,0.698888,1.3938715,2.0927596,2.7916477,3.4866312,3.1664703,2.8424048,2.5183394,2.1981785,1.8741131,1.5773785,1.2806439,0.98390937,0.6832704,0.38653582,4.5447245,8.702912,12.861101,17.019289,21.173573,22.950077,24.72658,26.499178,28.27568,30.048279,33.620808,37.193336,40.765865,44.33839,47.91092,46.794262,45.6776,44.560944,43.444283,42.32372,36.908314,31.489004,26.073599,20.654287,15.238882,15.406772,15.578565,15.746454,15.918248,16.086138,16.164225,16.242313,16.320402,16.398489,16.476578,16.050997,15.629322,15.207646,14.785972,14.364296,15.1061325,15.847969,16.589806,17.331642,18.073479,17.526861,16.976341,16.42582,15.875299,15.324779,18.74113,22.153578,25.569931,28.986282,32.39873,25.929136,19.459541,12.989946,6.520352,0.05075723,2.514435,4.9742084,7.437886,9.901564,12.361338,11.428185,10.491129,9.557977,8.62092,7.687768,8.929368,10.167064,11.408664,12.6463585,13.887959,16.613232,19.34241,22.071587,24.796858,27.526035,23.930082,20.334127,16.738173,13.146122,9.550168,7.758047,5.969831,4.181615,2.3894942,0.60127795,0.80821127,1.0190489,1.2298868,1.4407244,1.6515622,1.4407244,1.2298868,1.0190489,0.80821127,0.60127795,1.5695697,2.541766,3.5100577,4.478349,5.4505453,5.563773,5.6730967,5.786324,5.899552,6.012779,6.211904,6.4110284,6.6140575,6.813182,7.012306,5.6848097,4.357313,3.0298162,1.7023194,0.37482262,2.7018464,5.02887,7.355894,9.686822,12.013845,13.232019,14.454097,15.672271,16.890444,18.112522,14.50095,10.893282,7.28171,3.6740425,0.062470436,2.2723622,4.482254,6.6921453,8.902037,11.111929,10.479416,9.846903,9.21439,8.581876,7.9493628,8.183627,8.413987,8.648251,8.878611,9.112875,9.245625,9.378374,9.511124,9.643873,9.776623,8.121157,6.46569,4.8102236,3.154757,1.4992905,1.319688,1.1400855,0.96048295,0.78088045,0.60127795,0.5388075,0.48024148,0.42167544,0.359205,0.30063897,1.2376955,2.174752,3.1118085,4.0488653,4.985922,3.9902992,2.9907722,1.9951496,0.9956226,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07027924,0.14055848,0.21083772,0.28111696,0.3513962,0.58566034,0.8238289,1.0619974,1.3001659,1.5383345,1.5695697,1.6008049,1.6359446,1.6671798,1.698415,1.4016805,1.1049459,0.80821127,0.5114767,0.21083772,0.38263142,0.5544251,0.7223144,0.8941081,1.0619974,2.233318,3.4007344,4.572055,5.743376,6.910792,5.6965227,4.482254,3.2679846,2.0537157,0.8394465,0.6910792,0.5427119,0.39434463,0.24597734,0.10151446,0.093705654,0.08589685,0.078088045,0.07027924,0.062470436,0.28111696,0.4958591,0.7145056,0.93315214,1.1517987,1.0815194,1.0151446,0.94876975,0.8784905,0.81211567,0.76135844,0.7106012,0.6637484,0.61299115,0.5622339,0.71841,0.8784905,1.0346665,1.1908426,1.3509232,2.0146716,2.67842,3.3460727,4.009821,4.6735697,4.4705405,4.263607,4.0605783,3.853645,3.6506162,3.6467118,3.6467118,3.6428072,3.638903,3.638903,3.408543,3.1781836,2.9478238,2.717464,2.4871042,2.0810463,1.6710842,1.2650263,0.8589685,0.44900626,0.58175594,0.7145056,0.8472553,0.98000497,1.1127546,1.0112402,0.9058213,0.80430686,0.7027924,0.60127795,0.59737355,0.59346914,0.59346914,0.58956474,0.58566034,0.5388075,0.48805028,0.43729305,0.38653582,0.3357786,0.3240654,0.31235218,0.30063897,0.28892577,0.27330816,0.27330816,0.27330816,0.27330816,0.27330816,0.27330816,0.26159495,0.24988174,0.23816854,0.22645533,0.21083772,25.624592,22.67677,19.728945,16.78112,13.833297,10.889378,9.913278,8.941081,7.968885,6.996689,6.0244927,5.630148,5.2358036,4.841459,4.4432096,4.0488653,3.697469,3.3460727,2.9907722,2.639376,2.2879796,1.9600099,1.6320401,1.3040704,0.97610056,0.6481308,0.80821127,0.96438736,1.1205635,1.2806439,1.43682,1.1713207,0.9058213,0.6442264,0.37872702,0.113227665,0.3279698,0.5427119,0.75745404,0.97219616,1.1869383,2.4441557,3.697469,4.950782,6.2079997,7.461313,8.519405,9.577498,10.6355915,11.693685,12.751778,18.256985,23.766096,29.271303,34.780415,40.28562,40.23877,40.18801,40.137257,40.0865,40.03574,37.825848,35.612053,33.39826,31.188366,28.97457,30.399675,31.824783,33.24989,34.674995,36.1001,32.699368,29.298634,25.8979,22.50107,19.100336,16.02757,12.954806,9.882042,6.8092775,3.736513,4.958591,6.1767645,7.3988423,8.617016,9.839094,8.246098,6.6531014,5.0601053,3.4671092,1.8741131,1.7999294,1.7257458,1.6515622,1.5734742,1.4992905,1.7413634,1.9834363,2.2294137,2.4714866,2.7135596,2.194274,1.678893,1.1596074,0.6442264,0.12494087,0.20693332,0.28502136,0.3631094,0.44510186,0.5231899,0.59346914,0.6637484,0.7340276,0.80430686,0.8745861,1.8506867,2.8306916,3.8067923,4.786797,5.7628975,5.657479,5.55206,5.446641,5.3412223,5.2358036,5.852699,6.46569,7.082586,7.6955767,8.312472,9.304191,10.295909,11.291532,12.28325,13.274967,10.768341,8.265619,5.758993,3.2562714,0.74964523,0.8511597,0.95657855,1.0580931,1.1596074,1.261122,3.174279,5.083532,6.9927845,8.902037,10.81129,10.25296,9.690726,9.132397,8.574067,8.011833,8.460839,8.905942,9.354948,9.803954,10.249056,12.34572,14.438479,16.535143,18.631807,20.724567,20.19357,19.658665,19.127666,18.596668,18.061766,14.981192,11.896713,8.81614,5.7316628,2.6510892,2.7213683,2.7916477,2.8619268,2.9283018,2.998581,3.0883822,3.174279,3.2640803,3.349977,3.435874,3.4514916,3.4632049,3.474918,3.4866312,3.4983444,3.1313305,2.7643168,2.397303,2.0302892,1.6632754,1.4407244,1.2181735,0.9956226,0.77307165,0.5505207,0.48024148,0.40996224,0.339683,0.26940376,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.046852827,0.08980125,0.13665408,0.1796025,0.22645533,0.26940376,0.30844778,0.3513962,0.39434463,0.43729305,0.57394713,0.7106012,0.8511597,0.9878138,1.1244678,1.0307622,0.93315214,0.8394465,0.74574083,0.6481308,0.5427119,0.43338865,0.3279698,0.21864653,0.113227665,0.23426414,0.359205,0.48024148,0.60127795,0.7262188,0.7262188,0.7301232,0.7340276,0.7340276,0.737932,1.1635119,1.5890918,2.0107672,2.436347,2.8619268,2.3894942,1.9170616,1.4446288,0.97219616,0.4997635,2.5066261,4.5095844,6.5164475,8.519405,10.526268,12.025558,13.528754,15.031949,16.535143,18.038338,15.274021,12.5058,9.741484,6.9771667,4.21285,4.298747,4.380739,4.466636,4.552533,4.6384296,4.9156423,5.192855,5.4700675,5.74728,6.0244927,4.8375545,3.6506162,2.463678,1.2767396,0.08589685,0.3631094,0.6442264,0.92143893,1.1986516,1.475864,3.4710135,5.466163,7.461313,9.456462,11.4516115,10.901091,10.350571,9.80005,9.249529,8.699008,8.121157,7.5394006,6.9615493,6.379793,5.7980375,6.8561306,7.914223,8.972317,10.03041,11.088503,11.307149,11.525795,11.748346,11.966993,12.185639,9.749292,7.3129454,4.8765984,2.436347,0.0,0.92924774,1.8584955,2.7916477,3.7208953,4.650143,4.0332475,3.416352,2.795552,2.1786566,1.5617609,1.3431144,1.1283722,0.9097257,0.6910792,0.47633708,5.185046,9.893755,14.606369,19.315079,24.023787,22.938364,21.849035,20.76361,19.674282,18.58886,24.16825,29.74764,35.32703,40.90642,46.485813,45.958717,45.431625,44.90453,44.377438,43.85034,38.157722,32.46901,26.780294,21.091581,15.398962,16.023666,16.644466,17.26917,17.88997,18.51077,18.756748,19.002726,19.248703,19.490776,19.736753,18.88169,18.026625,17.17156,16.316498,15.461433,16.902157,18.342882,19.783606,21.22433,22.66115,21.376602,20.08815,18.799696,17.511244,16.226696,20.80656,25.390327,29.974096,34.55396,39.13773,31.313307,23.492788,15.668366,7.8478484,0.023426414,3.310933,6.5984397,9.885946,13.173453,16.46096,15.21936,13.97776,12.73616,11.490656,10.249056,9.921086,9.589212,9.261242,8.929368,8.601398,12.193448,15.789403,19.385357,22.981312,26.573362,22.352703,18.132044,13.907481,9.686822,5.462259,4.5291066,3.5959544,2.6667068,1.7335546,0.80040246,1.0659018,1.3353056,1.6008049,1.8702087,2.135708,1.8702087,1.6008049,1.3353056,1.0659018,0.80040246,1.6476578,2.494913,3.3421683,4.1894236,5.036679,5.263134,5.4856853,5.7121406,5.938596,6.1611466,6.461786,6.7624245,7.0630636,7.363703,7.6643414,6.2158084,4.7711797,3.3265507,1.8819219,0.43729305,1.7335546,3.0259118,4.322173,5.618435,6.910792,7.4847393,8.058686,8.628729,9.202676,9.776623,7.832231,5.891743,3.9473507,2.0068626,0.062470436,1.8311646,3.5959544,5.364649,7.1333427,8.898132,8.6131115,8.32809,8.043069,7.758047,7.47693,7.8478484,8.218767,8.59359,8.964508,9.339331,9.198771,9.058213,8.917655,8.777096,8.636538,7.2582836,5.883934,4.50568,3.1274261,1.7491722,1.5617609,1.3704453,1.1791295,0.9917182,0.80040246,0.71841,0.64032197,0.5583295,0.48024148,0.39824903,1.6515622,2.900971,4.1503797,5.3997884,6.649197,5.3217,3.9902992,2.6588979,1.3314011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.37482262,0.57394713,0.77307165,0.97610056,1.175225,1.2845483,1.3938715,1.5031948,1.6164225,1.7257458,1.4055848,1.0893283,0.77307165,0.45681506,0.13665408,0.28502136,0.43338865,0.58175594,0.7262188,0.8745861,2.436347,3.9942036,5.5559645,7.113821,8.675582,7.141152,5.610626,4.0761957,2.5456703,1.0112402,0.8199245,0.62860876,0.43338865,0.24207294,0.05075723,0.05075723,0.05466163,0.058566034,0.058566034,0.062470436,0.3513962,0.6442264,0.93315214,1.2220778,1.5110037,1.4212024,1.3314011,1.2415999,1.1517987,1.0619974,0.999527,0.93705654,0.8745861,0.81211567,0.74964523,0.93315214,1.1205635,1.3040704,1.4914817,1.6749885,2.494913,3.3148375,4.134762,4.9546866,5.774611,5.349031,4.919547,4.493967,4.0644827,3.638903,3.6818514,3.7208953,3.7638438,3.8067923,3.8497405,3.736513,3.619381,3.506153,3.3890212,3.2757936,2.7291772,2.1786566,1.6320401,1.0854238,0.5388075,0.7106012,0.8823949,1.0541886,1.2259823,1.4016805,1.2533131,1.1088502,0.96438736,0.8199245,0.6754616,0.6676528,0.659844,0.6520352,0.6442264,0.63641757,0.57394713,0.5114767,0.44900626,0.38653582,0.3240654,0.31235218,0.30063897,0.28892577,0.27330816,0.26159495,0.26159495,0.26159495,0.26159495,0.26159495,0.26159495,0.24988174,0.23816854,0.22645533,0.21083772,0.19912452,31.750599,27.537748,23.3249,19.11205,14.899199,10.686349,9.288573,7.8868923,6.4891167,5.087436,3.6857557,3.5764325,3.4632049,3.349977,3.2367494,3.1235218,2.900971,2.6745155,2.4480603,2.2255092,1.999054,1.7608855,1.5266213,1.2884527,1.0502841,0.81211567,0.94876975,1.0893283,1.2259823,1.3626363,1.4992905,1.2259823,0.94876975,0.6754616,0.39824903,0.12494087,0.31235218,0.4997635,0.6871748,0.8745861,1.0619974,2.6003318,4.138666,5.6730967,7.211431,8.749765,9.101162,9.448653,9.80005,10.151445,10.498938,16.55076,22.59868,28.650503,34.69842,40.750248,41.023556,41.300766,41.574074,41.851288,42.124596,40.7112,39.301712,37.88832,36.474926,35.06153,35.53787,36.014206,36.48664,36.962975,37.439312,31.285975,25.136541,18.987108,12.837675,6.688241,6.239235,5.786324,5.337318,4.8883114,4.4393053,4.900025,5.3607445,5.825368,6.2860875,6.7507114,5.688714,4.6267166,3.5608149,2.4988174,1.43682,1.1517987,0.8628729,0.57394713,0.28892577,0.0,0.6637484,1.3235924,1.9873407,2.6510892,3.310933,2.6510892,1.9873407,1.3235924,0.6637484,0.0,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,0.6871748,0.74964523,0.81211567,0.8745861,0.93705654,2.174752,3.4124475,4.650143,5.8878384,7.125534,6.387602,5.64967,4.911738,4.173806,3.435874,4.0996222,4.7633705,5.423215,6.086963,6.7507114,7.8517528,8.94889,10.049932,11.150972,12.24811,9.975748,7.699481,5.423215,3.1508527,0.8745861,0.8394465,0.80040246,0.76135844,0.7262188,0.6871748,3.049338,5.4115014,7.773665,10.135828,12.501896,11.974802,11.4516115,10.924518,10.401327,9.874233,9.663396,9.448653,9.237816,9.023073,8.812236,11.951375,15.086611,18.22575,21.360985,24.500124,24.023787,23.551353,23.075018,22.59868,22.126247,18.338978,14.551707,10.760532,6.9732623,3.1859922,2.9361105,2.6862288,2.436347,2.1864653,1.9365835,2.35045,2.7643168,3.174279,3.5881457,3.998108,3.310933,2.6237583,1.9365835,1.2494087,0.5622339,0.4997635,0.43729305,0.37482262,0.31235218,0.24988174,0.3357786,0.42557985,0.5114767,0.60127795,0.6871748,0.60127795,0.5114767,0.42557985,0.3357786,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.76135844,1.4641509,2.1630387,2.8619268,3.5608149,2.900971,2.2372224,1.5734742,0.9136301,0.24988174,2.35045,4.4510183,6.551587,8.648251,10.748819,11.560935,12.373051,13.189071,14.001186,14.813302,12.400381,9.987461,7.57454,5.1616197,2.7486992,3.2484627,3.7482262,4.251894,4.7516575,5.251421,5.4505453,5.64967,5.8487945,6.0518236,6.250948,5.001539,3.7482262,2.4988174,1.2494087,0.0,0.3240654,0.6481308,0.97610056,1.3001659,1.6242313,3.78727,5.950309,8.113348,10.276386,12.439425,11.076789,9.714153,8.351517,6.98888,5.6262436,5.2358036,4.8492675,4.462732,4.0761957,3.6857557,5.6379566,7.5862536,9.538455,11.486752,13.438952,13.423335,13.411622,13.399908,13.388195,13.376482,10.701966,8.023546,5.349031,2.6745155,0.0,1.1635119,2.3231194,3.4866312,4.650143,5.813655,4.900025,3.9863946,3.076669,2.1630387,1.2494087,1.1127546,0.97610056,0.8394465,0.698888,0.5622339,5.825368,11.088503,16.351637,21.610867,26.874,22.926651,18.975395,15.024139,11.076789,7.125534,14.711788,22.29804,29.888199,37.474453,45.060707,45.123177,45.185646,45.24812,45.31059,45.37306,39.411037,33.449013,27.486992,21.52497,15.562947,16.636658,17.714273,18.787983,19.861694,20.93931,21.349272,21.763138,22.1731,22.586967,23.000834,21.712381,20.423927,19.13938,17.850927,16.562475,18.698183,20.837795,22.973503,25.113115,27.248823,25.226343,23.199959,21.173573,19.151093,17.124708,22.875893,28.623173,34.37436,40.12554,45.876728,36.70138,27.526035,18.35069,9.175345,0.0,4.1113358,8.226576,12.337912,16.449247,20.560583,19.010534,17.464392,15.914344,14.364296,12.814248,10.912805,9.01136,7.113821,5.212377,3.310933,7.773665,12.236397,16.69913,21.16186,25.624592,20.775324,15.926057,11.076789,6.223617,1.3743496,1.3001659,1.2259823,1.1517987,1.0737107,0.999527,1.3235924,1.6515622,1.9756275,2.2996929,2.6237583,2.2996929,1.9756275,1.6515622,1.3235924,0.999527,1.7257458,2.4480603,3.174279,3.900498,4.6267166,4.9624953,5.298274,5.6379566,5.9737353,6.3134184,6.7116675,7.113821,7.5120697,7.914223,8.312472,6.7507114,5.1889505,3.6232853,2.0615244,0.4997635,0.76135844,1.0268579,1.2884527,1.5500476,1.8116426,1.737459,1.6632754,1.5890918,1.5110037,1.43682,1.1635119,0.8862993,0.61299115,0.3357786,0.062470436,1.3860629,2.7135596,4.037152,5.3607445,6.688241,6.7507114,6.813182,6.8756523,6.9381227,7.000593,7.5120697,8.023546,8.538928,9.050405,9.561881,9.151918,8.738052,8.324185,7.914223,7.5003567,6.3993154,5.298274,4.2011366,3.1000953,1.999054,1.7999294,1.6008049,1.4016805,1.1986516,0.999527,0.9019169,0.80040246,0.698888,0.60127795,0.4997635,2.0615244,3.6232853,5.1889505,6.7507114,8.312472,6.649197,4.985922,3.3265507,1.6632754,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1639849,0.3240654,0.48805028,0.6481308,0.81211567,0.999527,1.1869383,1.3743496,1.5617609,1.7491722,1.4133936,1.0737107,0.737932,0.39824903,0.062470436,0.18741131,0.31235218,0.43729305,0.5622339,0.6871748,2.639376,4.5876727,6.5359693,8.488171,10.436467,8.58578,6.7389984,4.8883114,3.0376248,1.1869383,0.94876975,0.7106012,0.47633708,0.23816854,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.42557985,0.78868926,1.1517987,1.5110037,1.8741131,1.7608855,1.6515622,1.5383345,1.4251068,1.3118792,1.2376955,1.1635119,1.0893283,1.0112402,0.93705654,1.1517987,1.3626363,1.5734742,1.7882162,1.999054,2.9751544,3.951255,4.9234514,5.899552,6.8756523,6.223617,5.575486,4.9234514,4.2753205,3.6232853,3.7130866,3.7989833,3.8887846,3.9746814,4.0605783,4.0605783,4.0605783,4.0605783,4.0605783,4.0605783,3.3734035,2.6862288,1.999054,1.3118792,0.62470436,0.8394465,1.0502841,1.261122,1.475864,1.6867018,1.4992905,1.3118792,1.1244678,0.93705654,0.74964523,0.737932,0.7262188,0.7106012,0.698888,0.6871748,0.61299115,0.5388075,0.46071947,0.38653582,0.31235218,0.30063897,0.28892577,0.27330816,0.26159495,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.23816854,0.22645533,0.21083772,0.19912452,0.18741131,25.987701,22.739239,19.486872,16.238409,12.986042,9.737579,8.503788,7.2739015,6.04011,4.806319,3.5764325,3.3890212,3.2055142,3.018103,2.8345962,2.6510892,2.475391,2.2996929,2.1239948,1.9482968,1.7765031,1.5539521,1.3353056,1.116659,0.8941081,0.6754616,0.9136301,1.1517987,1.3860629,1.6242313,1.8623998,2.67842,3.4905357,4.3065557,5.1225758,5.938596,6.899079,7.8634663,8.823949,9.788337,10.748819,11.549222,12.34572,13.142218,13.938716,14.739119,13.903577,13.0719385,12.240301,11.408664,10.573121,15.781594,20.986162,26.190731,31.395298,36.599865,36.38903,36.178192,35.971256,35.76042,35.549583,34.089336,32.62909,31.168842,29.708597,28.24835,29.111223,29.974096,30.83697,31.699842,32.562714,27.436235,22.305851,17.17937,12.05289,6.9264097,6.4149327,5.903456,5.395884,4.884407,4.376835,4.591577,4.8102236,5.02887,5.2436123,5.462259,4.743849,4.029343,3.310933,2.592523,1.8741131,1.4992905,1.1244678,0.74964523,0.37482262,0.0,0.6871748,1.3743496,2.0615244,2.7486992,3.435874,3.3538816,3.2679846,3.182088,3.096191,3.0141985,2.5105307,2.0107672,1.5110037,1.0112402,0.5114767,0.5700427,0.62860876,0.6832704,0.7418364,0.80040246,1.7843118,2.7643168,3.7482262,4.728231,5.7121406,5.606722,5.5013027,5.395884,5.2943697,5.1889505,5.883934,6.578918,7.2739015,7.968885,8.663869,9.433036,10.202203,10.971371,11.744442,12.513609,10.436467,8.359325,6.278279,4.2011366,2.1239948,2.15523,2.1864653,2.2137961,2.2450314,2.2762666,3.8692627,5.4583545,7.0513506,8.644346,10.237343,9.858616,9.483793,9.105066,8.726339,8.351517,8.171914,7.996216,7.816613,7.6409154,7.461313,9.897659,12.334006,14.766449,17.202797,19.639143,19.303364,18.967587,18.631807,18.296028,17.964155,15.223265,12.486279,9.749292,7.012306,4.2753205,3.8263142,3.3812122,2.9322062,2.4831998,2.0380979,2.3699722,2.7018464,3.0337205,3.3655949,3.7013733,3.049338,2.4012074,1.7491722,1.1010414,0.44900626,0.39824903,0.3513962,0.30063897,0.24988174,0.19912452,0.28111696,0.359205,0.44119745,0.5192855,0.60127795,0.5231899,0.44510186,0.3670138,0.28892577,0.21083772,0.1756981,0.14055848,0.10932326,0.07418364,0.039044023,0.039044023,0.042948425,0.046852827,0.046852827,0.05075723,0.14055848,0.23426414,0.3279698,0.42167544,0.5114767,0.45291066,0.39434463,0.3318742,0.27330816,0.21083772,0.1717937,0.12884527,0.08589685,0.042948425,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.80821127,1.4290112,2.0459068,2.6667068,3.2875066,3.06886,2.854118,2.6354716,2.416825,2.1981785,3.5022488,4.806319,6.1064854,7.4105554,8.710721,9.483793,10.25296,11.022127,11.791295,12.564366,10.491129,8.4178915,6.3446536,4.271416,2.1981785,2.6276627,3.0532427,3.4827268,3.9083066,4.337791,4.806319,5.270943,5.7394714,6.2079997,6.676528,5.6535745,4.630621,3.6076677,2.5847144,1.5617609,1.7725986,1.9834363,2.194274,2.4012074,2.612045,4.126953,5.6418614,7.1567693,8.671678,10.186585,9.253433,8.324185,7.3910336,6.4578815,5.5247293,5.278752,5.036679,4.7907014,4.5447245,4.298747,5.7316628,7.1606736,8.589685,10.018696,11.4516115,11.607788,11.763964,11.924045,12.08022,12.236397,9.792241,7.348085,4.903929,2.455869,0.011713207,1.3001659,2.5886188,3.873167,5.1616197,6.4500723,5.4427366,4.435401,3.4280653,2.4207294,1.4133936,1.3665408,1.3235924,1.2767396,1.2337911,1.1869383,5.3217,9.452558,13.583415,17.718178,21.849035,19.318983,16.788929,14.258877,11.728825,9.198771,15.012426,20.826082,26.635832,32.449486,38.26314,38.911274,39.559402,40.20363,40.85176,41.499893,37.310467,33.121044,28.931622,24.738293,20.548868,20.77142,20.990067,21.208714,21.431265,21.64991,22.34099,23.035973,23.727053,24.41813,25.113115,23.625538,22.141865,20.658192,19.170614,17.686943,19.276033,20.861221,22.450314,24.039404,25.624592,23.418604,21.208714,19.002726,16.796738,14.586847,19.596195,24.605543,29.618795,34.628143,39.637493,32.476818,25.316145,18.15547,10.998701,3.8380275,6.3915067,8.941081,11.49456,14.048039,16.601519,15.336493,14.0714655,12.806439,11.541413,10.276386,8.749765,7.223144,5.700427,4.173806,2.6510892,6.98888,11.326671,15.664462,19.998348,24.33614,19.689901,15.043662,10.393518,5.74728,1.1010414,1.0580931,1.0190489,0.98000497,0.94096094,0.9019169,1.1400855,1.3782539,1.620327,1.8584955,2.1005683,1.8389735,1.5812829,1.319688,1.0580931,0.80040246,1.5969005,2.3933985,3.193801,3.9902992,4.786797,4.845363,4.903929,4.958591,5.017157,5.0757227,5.3919797,5.708236,6.028397,6.3446536,6.66091,5.5442514,4.4275923,3.310933,2.194274,1.0737107,1.678893,2.2840753,2.8892577,3.49444,4.0996222,3.533484,2.9634414,2.397303,1.8311646,1.261122,1.0190489,0.77697605,0.5349031,0.29283017,0.05075723,1.1244678,2.194274,3.2679846,4.3416953,5.4115014,5.5832953,5.7511845,5.9229784,6.0908675,6.262661,6.7429028,7.223144,7.703386,8.183627,8.663869,8.62092,8.577971,8.535024,8.492075,8.449126,7.5159745,6.5867267,5.6535745,4.7204223,3.78727,3.349977,2.912684,2.475391,2.0380979,1.6008049,1.698415,1.796025,1.893635,1.9912452,2.0888553,3.3890212,4.689187,5.989353,7.2856145,8.58578,7.008402,5.4310236,3.853645,2.2762666,0.698888,0.5583295,0.42167544,0.28111696,0.14055848,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12884527,0.26159495,0.39044023,0.5192855,0.6481308,0.80040246,0.94876975,1.1010414,1.2494087,1.4016805,1.1361811,0.8745861,0.61299115,0.3513962,0.08589685,0.21474212,0.3435874,0.46852827,0.59737355,0.7262188,3.182088,5.6379566,8.097731,10.553599,13.013372,10.869856,8.726339,6.5867267,4.4432096,2.2996929,1.8389735,1.3782539,0.92143893,0.46071947,0.0,0.10932326,0.21864653,0.3318742,0.44119745,0.5505207,0.81211567,1.0737107,1.33921,1.6008049,1.8623998,1.9756275,2.0927596,2.2059872,2.3231194,2.436347,2.1864653,1.9326792,1.678893,1.4290112,1.175225,1.4055848,1.639849,1.8741131,2.1044729,2.338737,3.174279,4.0137253,4.8492675,5.688714,6.524256,6.3134184,6.098676,5.8878384,5.6730967,5.462259,5.173333,4.8883114,4.5993857,4.3143644,4.025439,4.0761957,4.126953,4.173806,4.224563,4.2753205,3.6701381,3.0649557,2.4597735,1.8545911,1.2494087,1.3665408,1.4836729,1.6008049,1.7218413,1.8389735,1.6320401,1.4290112,1.2220778,1.0190489,0.81211567,0.8316377,0.8511597,0.8706817,0.8941081,0.9136301,0.94096094,0.96829176,0.9956226,1.0229534,1.0502841,0.8941081,0.7340276,0.57785153,0.42167544,0.26159495,0.25378615,0.24207294,0.23426414,0.22255093,0.21083772,0.20302892,0.19131571,0.1835069,0.1717937,0.1639849,20.224804,17.936825,15.648844,13.360865,11.076789,8.78881,7.7229075,6.657006,5.591104,4.5291066,3.4632049,3.2055142,2.9478238,2.690133,2.4324427,2.174752,2.0498111,1.9248703,1.7999294,1.6749885,1.5500476,1.3470187,1.1439898,0.94096094,0.7418364,0.5388075,0.8745861,1.2142692,1.5500476,1.8858263,2.2255092,4.1308575,6.036206,7.941554,9.846903,11.748346,13.4858055,15.223265,16.960724,18.698183,20.435642,20.494207,20.552773,20.61134,20.666,20.724567,18.709896,16.695225,14.6805525,12.665881,10.651209,15.008522,19.36974,23.730957,28.08827,32.449486,31.754503,31.05952,30.364536,29.669552,28.97457,27.46747,25.960371,24.453272,22.946173,21.439074,22.688482,23.937891,25.1873,26.436708,27.686117,23.58259,19.479063,15.371632,11.268105,7.1606736,6.590631,6.0205884,5.4505453,4.884407,4.3143644,4.283129,4.2557983,4.2284675,4.2011366,4.173806,3.802888,3.4280653,3.057147,2.6862288,2.3114061,1.8506867,1.3860629,0.92534333,0.46071947,0.0,0.7106012,1.4251068,2.135708,2.8502135,3.5608149,4.056674,4.548629,5.040583,5.532538,6.0244927,4.900025,3.775557,2.6510892,1.5266213,0.39824903,0.45291066,0.5036679,0.5583295,0.60908675,0.6637484,1.3899672,2.1161861,2.8463092,3.5725281,4.298747,4.825841,5.35684,5.883934,6.4110284,6.9381227,7.6643414,8.39056,9.120684,9.846903,10.573121,11.014318,11.455516,11.896713,12.334006,12.775204,10.893282,9.0152645,7.1333427,5.2553253,3.3734035,3.4710135,3.5686235,3.6662338,3.7638438,3.8614538,4.6852827,5.5091114,6.329036,7.152865,7.9766936,7.746334,7.5159745,7.2856145,7.055255,6.824895,6.6843367,6.5398736,6.3993154,6.2548523,6.114294,7.843944,9.577498,11.311053,13.040704,14.774258,14.579038,14.383818,14.188598,13.993378,13.798158,12.111456,10.424754,8.738052,7.0513506,5.3607445,4.716518,4.0722914,3.4280653,2.7838387,2.135708,2.3894942,2.6432803,2.893162,3.1469483,3.4007344,2.787743,2.174752,1.5617609,0.94876975,0.3357786,0.30063897,0.26159495,0.22645533,0.18741131,0.14836729,0.22255093,0.29673457,0.3670138,0.44119745,0.5114767,0.44510186,0.37872702,0.30844778,0.24207294,0.1756981,0.15617609,0.13665408,0.113227665,0.093705654,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.23426414,0.43338865,0.62860876,0.8277333,1.0268579,0.8667773,0.7106012,0.5544251,0.39434463,0.23816854,0.19131571,0.14055848,0.093705654,0.046852827,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.37482262,0.31235218,0.24988174,0.18741131,0.12494087,0.1639849,0.19912452,0.23816854,0.27330816,0.31235218,0.8511597,1.3938715,1.9326792,2.4714866,3.0141985,3.240654,3.4671092,3.6935644,3.9239242,4.1503797,4.6540475,5.1616197,5.6652875,6.168956,6.676528,7.4027467,8.128965,8.859089,9.585307,10.311526,8.581876,6.8483214,5.114767,3.3812122,1.6515622,2.0068626,2.358259,2.7135596,3.06886,3.4241607,4.1581883,4.8961205,5.630148,6.364176,7.098203,6.3056097,5.5091114,4.716518,3.9200199,3.1235218,3.2211318,3.3148375,3.408543,3.506153,3.5998588,4.466636,5.3334136,6.2040954,7.0708723,7.9376497,7.433982,6.9342184,6.4305506,5.9268827,5.423215,5.3217,5.2201858,5.1186714,5.0132523,4.911738,5.8214636,6.7311897,7.6409154,8.550641,9.464272,9.788337,10.116306,10.444276,10.772245,11.100216,8.886419,6.6687193,4.454923,2.241127,0.023426414,1.43682,2.8502135,4.263607,5.6730967,7.08649,5.985449,4.884407,3.7794614,2.67842,1.5734742,1.6242313,1.6710842,1.717937,1.7647898,1.8116426,4.814128,7.816613,10.819098,13.821584,16.82407,15.7152195,14.606369,13.493614,12.384764,11.275913,15.313066,19.350218,23.38737,27.424522,31.461674,32.695465,33.929256,35.15914,36.392933,37.626724,35.205994,32.78917,30.372345,27.95552,25.538694,24.902277,24.26586,23.633347,22.99693,22.364416,23.336613,24.30881,25.281004,26.2532,27.225397,25.542599,23.859802,22.177006,20.494207,18.81141,19.849981,20.888552,21.923218,22.96179,24.00036,21.610867,19.221373,16.827974,14.438479,12.0489855,16.320402,20.587914,24.85933,29.130745,33.39826,28.256159,23.110157,17.964155,12.818152,7.676055,8.667773,9.659492,10.651209,11.6468315,12.63855,11.6585455,10.67854,9.698535,8.718531,7.7385254,6.5867267,5.4388323,4.2870336,3.1391394,1.9873407,6.2001905,10.413041,14.625891,18.838741,23.05159,18.604477,14.161267,9.714153,5.270943,0.8238289,0.8199245,0.8160201,0.80821127,0.80430686,0.80040246,0.95657855,1.1088502,1.2650263,1.4212024,1.5734742,1.3782539,1.1869383,0.9917182,0.79649806,0.60127795,1.4719596,2.338737,3.2094188,4.0801005,4.950782,4.728231,4.50568,4.283129,4.0605783,3.8380275,4.0722914,4.3065557,4.5408196,4.7789884,5.0132523,4.3416953,3.6662338,2.9946766,2.3231194,1.6515622,2.5964274,3.5451972,4.493967,5.4388323,6.387602,5.3256044,4.267512,3.2094188,2.1474214,1.0893283,0.8784905,0.6676528,0.45681506,0.24597734,0.039044023,0.8589685,1.678893,2.4988174,3.3187418,4.138666,4.415879,4.6930914,4.970304,5.2475166,5.5247293,5.9737353,6.4188375,6.8678436,7.3168497,7.7619514,8.089922,8.4178915,8.745861,9.073831,9.4018,8.636538,7.871275,7.1060123,6.3407493,5.575486,4.900025,4.224563,3.5491016,2.87364,2.1981785,2.494913,2.7916477,3.084478,3.3812122,3.6740425,4.7126136,5.7511845,6.785851,7.824422,8.862993,7.3715115,5.8761253,4.3846436,2.893162,1.4016805,1.1205635,0.8394465,0.5583295,0.28111696,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09761006,0.19522011,0.29283017,0.39044023,0.48805028,0.60127795,0.7106012,0.8238289,0.93705654,1.0502841,0.8628729,0.6754616,0.48805028,0.30063897,0.113227665,0.24207294,0.3709182,0.5036679,0.63251317,0.76135844,3.7287042,6.6921453,9.659492,12.622932,15.586374,13.153932,10.717585,8.281238,5.8487945,3.4124475,2.7291772,2.0459068,1.3665408,0.6832704,0.0,0.20693332,0.41386664,0.62079996,0.8316377,1.038571,1.1986516,1.3626363,1.5266213,1.6867018,1.8506867,2.194274,2.533957,2.8775444,3.2211318,3.5608149,3.1313305,2.7018464,2.2723622,1.8428779,1.4133936,1.6632754,1.9170616,2.1708477,2.4207294,2.6745155,3.3734035,4.0761957,4.775084,5.473972,6.1767645,6.3993154,6.6257706,6.8483214,7.0747766,7.3012323,6.6374836,5.9737353,5.3138914,4.650143,3.9863946,4.087909,4.1894236,4.2870336,4.388548,4.4861584,3.9668727,3.4436827,2.920493,2.397303,1.8741131,1.8975395,1.9209659,1.9443923,1.9639144,1.9873407,1.7647898,1.542239,1.319688,1.097137,0.8745861,0.92924774,0.98000497,1.0307622,1.0854238,1.1361811,1.2689307,1.397776,1.5266213,1.6593709,1.7882162,1.4836729,1.183034,0.8784905,0.57785153,0.27330816,0.25378615,0.23426414,0.21474212,0.19522011,0.1756981,0.1678893,0.16008049,0.15227169,0.14446288,0.13665408,14.461906,13.138313,11.810817,10.487225,9.163632,7.8361354,6.9381227,6.044015,5.1460023,4.2479897,3.349977,3.018103,2.690133,2.358259,2.0302892,1.698415,1.6242313,1.5500476,1.475864,1.4016805,1.3235924,1.1400855,0.95657855,0.76916724,0.58566034,0.39824903,0.8355421,1.2767396,1.7140326,2.1513257,2.5886188,5.5832953,8.577971,11.572648,14.567325,17.562002,20.076437,22.586967,25.101402,27.611933,30.126368,29.443098,28.759827,28.076557,27.393286,26.71392,23.516214,20.31851,17.120804,13.923099,10.725393,14.239355,17.753317,21.271183,24.785145,28.299107,27.119978,25.94085,24.761719,23.578686,22.399555,20.845604,19.29165,17.733795,16.179844,14.625891,16.261835,17.901684,19.537628,21.173573,22.813423,19.728945,16.64837,13.563893,10.48332,7.3988423,6.7702336,6.141625,5.5091114,4.8805027,4.251894,3.978586,3.7052777,3.4319696,3.1586614,2.8892577,2.8580225,2.8306916,2.803361,2.77603,2.7486992,2.1981785,1.6515622,1.1010414,0.5505207,0.0,0.737932,1.475864,2.2137961,2.951728,3.6857557,4.755562,5.8292727,6.899079,7.968885,9.0386915,7.289519,5.5364423,3.78727,2.0380979,0.28892577,0.3357786,0.38263142,0.42948425,0.47633708,0.5231899,0.9956226,1.4680552,1.9443923,2.416825,2.8892577,4.0488653,5.2084727,6.36808,7.5276875,8.687295,9.448653,10.206107,10.967466,11.728825,12.486279,12.595602,12.708829,12.818152,12.927476,13.036799,11.354002,9.671205,7.988407,6.3056097,4.6267166,4.7907014,4.9546866,5.1186714,5.2865605,5.4505453,5.5013027,5.5559645,5.606722,5.661383,5.7121406,5.630148,5.548156,5.466163,5.3841705,5.298274,5.192855,5.083532,4.9781127,4.8687897,4.7633705,5.794133,6.8209906,7.8517528,8.882515,9.913278,9.858616,9.803954,9.749292,9.690726,9.636065,8.999647,8.36323,7.726812,7.08649,6.4500723,5.606722,4.7633705,3.9239242,3.0805733,2.2372224,2.4090161,2.5808098,2.7565079,2.9283018,3.1000953,2.5261483,1.9482968,1.3743496,0.80040246,0.22645533,0.19912452,0.1756981,0.14836729,0.12494087,0.10151446,0.1639849,0.23035973,0.29673457,0.359205,0.42557985,0.3670138,0.30844778,0.25378615,0.19522011,0.13665408,0.13274968,0.12884527,0.12103647,0.11713207,0.113227665,0.093705654,0.078088045,0.058566034,0.042948425,0.023426414,0.3279698,0.62860876,0.93315214,1.2337911,1.5383345,1.2806439,1.0268579,0.77307165,0.5192855,0.26159495,0.21083772,0.15617609,0.10541886,0.05075723,0.0,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,0.5388075,0.44900626,0.3631094,0.27330816,0.18741131,0.23816854,0.28892577,0.3357786,0.38653582,0.43729305,0.8980125,1.358732,1.8194515,2.2762666,2.736986,3.408543,4.084005,4.755562,5.4271193,6.098676,5.805846,5.5169206,5.22409,4.93126,4.6384296,5.3217,6.008875,6.6921453,7.37932,8.062591,6.6687193,5.278752,3.8848803,2.4910088,1.1010414,1.3821584,1.6632754,1.9482968,2.2294137,2.5105307,3.513962,4.5173936,5.520825,6.524256,7.523783,6.957645,6.3915067,5.8214636,5.2553253,4.689187,4.6657605,4.646239,4.6267166,4.607195,4.5876727,4.806319,5.02887,5.2475166,5.466163,5.688714,5.6145306,5.5442514,5.4700675,5.395884,5.3256044,5.364649,5.4036927,5.446641,5.4856853,5.5247293,5.9151692,6.3056097,6.6960497,7.08649,7.473026,7.9727893,8.468649,8.968412,9.464272,9.964035,7.9766936,5.9932575,4.0059166,2.0224805,0.039044023,1.5734742,3.1118085,4.650143,6.1884775,7.726812,6.5281606,5.3295093,4.1308575,2.9361105,1.737459,1.8780174,2.018576,2.1591344,2.2957885,2.436347,4.31046,6.180669,8.054782,9.928895,11.799104,12.111456,12.419904,12.728352,13.040704,13.349152,15.613705,17.874353,20.138906,22.399555,24.664108,26.479656,28.299107,30.114655,31.934107,33.749653,33.105427,32.4612,31.816975,31.168842,30.524616,29.033134,27.545557,26.054077,24.5665,23.075018,24.328331,25.581644,26.831053,28.084366,29.337679,27.455757,25.57774,23.695818,21.8178,19.935879,20.423927,20.911978,21.400028,21.888079,22.37613,19.803127,17.230127,14.657126,12.084125,9.511124,13.040704,16.574188,20.103767,23.633347,27.162926,24.031595,20.90417,17.772839,14.641508,11.514082,10.944039,10.377901,9.811763,9.24172,8.675582,7.9805984,7.2856145,6.590631,5.8956475,5.2006636,4.423688,3.6506162,2.87364,2.1005683,1.3235924,5.4115014,9.499411,13.58732,17.675228,21.763138,17.519053,13.2788725,9.034787,4.7907014,0.5505207,0.58175594,0.60908675,0.64032197,0.6715572,0.698888,0.76916724,0.8394465,0.9097257,0.98000497,1.0502841,0.92143893,0.78868926,0.659844,0.5309987,0.39824903,1.3431144,2.2840753,3.2289407,4.169902,5.1108627,4.6110992,4.1074314,3.6037633,3.1039999,2.6003318,2.7526035,2.9048753,3.057147,3.2094188,3.3616903,3.135235,2.9087796,2.67842,2.4519646,2.2255092,3.513962,4.806319,6.094772,7.3832245,8.675582,7.1216297,5.571582,4.01763,2.463678,0.9136301,0.7340276,0.5583295,0.37872702,0.20302892,0.023426414,0.59346914,1.1596074,1.7257458,2.2957885,2.8619268,3.2484627,3.631094,4.01763,4.4041657,4.786797,5.2006636,5.618435,6.0323014,6.446168,6.8639393,7.558923,8.257811,8.956698,9.651682,10.350571,9.753197,9.155824,8.55845,7.9610763,7.363703,6.4500723,5.5364423,4.6267166,3.7130866,2.7994564,3.2914112,3.7833657,4.279225,4.7711797,5.263134,6.036206,6.813182,7.5862536,8.36323,9.136301,7.7307167,6.321227,4.9156423,3.506153,2.1005683,1.678893,1.261122,0.8394465,0.42167544,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06637484,0.12884527,0.19522011,0.26159495,0.3240654,0.39824903,0.47633708,0.5505207,0.62470436,0.698888,0.58566034,0.47633708,0.3631094,0.24988174,0.13665408,0.26940376,0.40215343,0.5349031,0.6676528,0.80040246,4.271416,7.746334,11.217348,14.688361,18.163279,15.434102,12.708829,9.979652,7.2543793,4.5252023,3.619381,2.7135596,1.8116426,0.9058213,0.0,0.30454338,0.60908675,0.9136301,1.2181735,1.5266213,1.5890918,1.6515622,1.7140326,1.7765031,1.8389735,2.4090161,2.979059,3.5491016,4.1191444,4.689187,4.0801005,3.4710135,2.8658314,2.2567444,1.6515622,1.9209659,2.194274,2.4675822,2.7408905,3.0141985,3.5764325,4.138666,4.7009,5.263134,5.825368,6.4891167,7.1489606,7.812709,8.476458,9.136301,8.101635,7.0630636,6.0244927,4.985922,3.951255,4.0996222,4.251894,4.4002614,4.548629,4.7009,4.2597027,3.8185053,3.3812122,2.9400148,2.4988174,2.4285383,2.3543546,2.2840753,2.2098918,2.135708,1.8975395,1.6593709,1.4172981,1.1791295,0.93705654,1.0229534,1.1088502,1.1908426,1.2767396,1.3626363,1.5969005,1.8272603,2.0615244,2.2918842,2.5261483,2.077142,1.6281357,1.183034,0.7340276,0.28892577,0.25769055,0.22645533,0.19912452,0.1678893,0.13665408,0.13274968,0.12884527,0.12103647,0.11713207,0.113227665,8.699008,8.335898,7.9766936,7.6135845,7.250475,6.8873653,6.1572423,5.4271193,4.6969957,3.9668727,3.2367494,2.8345962,2.4324427,2.0302892,1.6281357,1.2259823,1.1986516,1.175225,1.1517987,1.1244678,1.1010414,0.93315214,0.76526284,0.59737355,0.42948425,0.26159495,0.80040246,1.33921,1.8741131,2.4129205,2.951728,7.0357327,11.119738,15.203742,19.29165,23.375656,26.663162,29.95067,33.23818,36.525684,39.81319,38.391987,36.96688,35.545677,34.124477,32.699368,28.31863,23.941795,19.561056,15.180316,10.799577,13.470188,16.140799,18.81141,21.478117,24.148727,22.485453,20.818274,19.154997,17.491722,15.824542,14.223738,12.619028,11.018223,9.413514,7.812709,9.839094,11.861574,13.887959,15.914344,17.936825,15.879204,13.817679,11.756155,9.698535,7.6370106,6.9459314,6.2587566,5.5676775,4.8765984,4.1894236,3.6701381,3.1508527,2.6354716,2.1161861,1.6008049,1.9170616,2.233318,2.5534792,2.8697357,3.1859922,2.5495746,1.9131571,1.2767396,0.63641757,0.0,0.76135844,1.5266213,2.2879796,3.049338,3.8106966,5.4583545,7.1060123,8.75367,10.401327,12.0489855,9.675109,7.3012323,4.9234514,2.5495746,0.1756981,0.21864653,0.26159495,0.30063897,0.3435874,0.38653582,0.60518235,0.8238289,1.038571,1.2572175,1.475864,3.2679846,5.0601053,6.852226,8.644346,10.436467,11.229061,12.021654,12.814248,13.606842,14.399435,14.180789,13.958238,13.739592,13.520945,13.298394,11.814721,10.331048,8.843472,7.3597984,5.8761253,6.1064854,6.3407493,6.571109,6.805373,7.0357327,6.321227,5.602817,4.884407,4.165997,3.4514916,3.513962,3.5803368,3.6467118,3.7091823,3.775557,3.7013733,3.631094,3.5569105,3.4866312,3.4124475,3.7404175,4.068387,4.396357,4.7243266,5.0483923,5.134289,5.2201858,5.3060827,5.388075,5.473972,5.8878384,6.3017054,6.7116675,7.125534,7.5394006,6.4969254,5.4583545,4.415879,3.377308,2.338737,2.4285383,2.522244,2.6159496,2.7057507,2.7994564,2.260649,1.7257458,1.1869383,0.6481308,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.10932326,0.1639849,0.22255093,0.28111696,0.3357786,0.28892577,0.24207294,0.19522011,0.14836729,0.10151446,0.10932326,0.12103647,0.12884527,0.14055848,0.14836729,0.12103647,0.093705654,0.06637484,0.039044023,0.011713207,0.42167544,0.8277333,1.2337911,1.6437533,2.0498111,1.698415,1.3431144,0.9917182,0.64032197,0.28892577,0.23035973,0.1717937,0.113227665,0.058566034,0.0,0.1639849,0.3240654,0.48805028,0.6481308,0.81211567,0.698888,0.58566034,0.47633708,0.3631094,0.24988174,0.31235218,0.37482262,0.43729305,0.4997635,0.5622339,0.94096094,1.3235924,1.7023194,2.0810463,2.463678,3.5803368,4.6969957,5.813655,6.9342184,8.050878,6.9615493,5.8683167,4.7789884,3.68966,2.6003318,3.240654,3.8848803,4.5291066,5.169429,5.813655,4.759466,3.7091823,2.6549935,1.6008049,0.5505207,0.76135844,0.96829176,1.1791295,1.3899672,1.6008049,2.8697357,4.138666,5.4115014,6.6804323,7.9493628,7.60968,7.269997,6.930314,6.590631,6.250948,6.114294,5.9815445,5.84489,5.708236,5.575486,5.1460023,4.7204223,4.290938,3.8653584,3.435874,3.795079,4.154284,4.5095844,4.8687897,5.22409,5.407597,5.591104,5.7707067,5.9542136,6.13772,6.008875,5.8761253,5.74728,5.618435,5.4856853,6.153338,6.8209906,7.4886436,8.156297,8.823949,7.0708723,5.3138914,3.5608149,1.8038338,0.05075723,1.7140326,3.3734035,5.036679,6.699954,8.36323,7.0708723,5.7785153,4.4861584,3.193801,1.901444,2.1318035,2.366068,2.5964274,2.8306916,3.0610514,3.8067923,4.548629,5.290465,6.0323014,6.774138,8.503788,10.2334385,11.966993,13.696643,15.426293,15.914344,16.398489,16.88654,17.37459,17.86264,20.263847,22.668959,25.070168,27.471375,29.876486,31.000954,32.129326,33.257698,34.38607,35.514442,33.167896,30.821352,28.47871,26.132164,23.785618,25.32005,26.850574,28.385004,29.919434,31.44996,29.372818,27.295675,25.218534,23.141392,21.06425,21.00178,20.93931,20.876839,20.81437,20.751898,17.99539,15.238882,12.486279,9.729771,6.9732623,9.76491,12.556558,15.344301,18.135948,20.92369,19.810938,18.694279,17.581524,16.464865,15.348206,13.224211,11.096312,8.968412,6.8405128,4.7126136,4.3026514,3.892689,3.4827268,3.0727646,2.6628022,2.260649,1.8623998,1.4641509,1.0619974,0.6637484,4.6267166,8.58578,12.548749,16.511717,20.474686,16.43363,12.396477,8.355421,4.3143644,0.27330816,0.339683,0.40605783,0.46852827,0.5349031,0.60127795,0.58566034,0.5700427,0.5544251,0.5388075,0.5231899,0.46071947,0.39434463,0.3318742,0.26549935,0.19912452,1.2142692,2.2294137,3.2445583,4.2597027,5.2748475,4.493967,3.7091823,2.9283018,2.1435168,1.3626363,1.4329157,1.5031948,1.5734742,1.6437533,1.7140326,1.9287747,2.1474214,2.366068,2.5808098,2.7994564,4.4314966,6.0635366,7.699481,9.331521,10.963562,8.917655,6.871748,4.825841,2.7838387,0.737932,0.59346914,0.44900626,0.30063897,0.15617609,0.011713207,0.3279698,0.6442264,0.95657855,1.2728351,1.5890918,2.0810463,2.5730011,3.0649557,3.5569105,4.0488653,4.4314966,4.814128,5.196759,5.579391,5.9620223,7.0318284,8.097731,9.163632,10.2334385,11.29934,10.869856,10.4403715,10.010887,9.581403,9.151918,8.00012,6.8483214,5.700427,4.548629,3.4007344,4.0918136,4.7789884,5.4700675,6.1611466,6.8483214,7.363703,7.8751793,8.386656,8.898132,9.413514,8.089922,6.7663293,5.446641,4.123049,2.7994564,2.241127,1.678893,1.1205635,0.5583295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.06637484,0.09761006,0.12884527,0.1639849,0.19912452,0.23816854,0.27330816,0.31235218,0.3513962,0.31235218,0.27330816,0.23816854,0.19912452,0.1639849,0.29673457,0.43338865,0.5661383,0.7027924,0.8394465,4.8180323,8.796618,12.779109,16.757694,20.73628,17.718178,14.69617,11.678067,8.65606,5.6379566,4.5095844,3.3812122,2.2567444,1.1283722,0.0,0.40215343,0.80430686,1.2064602,1.6086137,2.0107672,1.9756275,1.9365835,1.901444,1.8623998,1.8233559,2.6237583,3.4202564,4.2167544,5.0132523,5.813655,5.02887,4.2440853,3.4593005,2.6706111,1.8858263,2.1786566,2.4714866,2.7643168,3.057147,3.349977,3.775557,4.2011366,4.6267166,5.0483923,5.473972,6.575013,7.676055,8.773191,9.874233,10.975275,9.561881,8.148487,6.7389984,5.3256044,3.912211,4.1113358,4.3143644,4.513489,4.7126136,4.911738,4.5564375,4.1972322,3.8419318,3.4827268,3.1235218,2.9556324,2.7916477,2.6237583,2.455869,2.2879796,2.0302892,1.7725986,1.5149081,1.2572175,0.999527,1.116659,1.2337911,1.3509232,1.4680552,1.5890918,1.9209659,2.2567444,2.592523,2.9283018,3.2640803,2.6706111,2.077142,1.4836729,0.8941081,0.30063897,0.26159495,0.21864653,0.1796025,0.14055848,0.10151446,0.09761006,0.093705654,0.093705654,0.08980125,0.08589685,2.9361105,3.5373883,4.138666,4.73604,5.337318,5.938596,5.376362,4.814128,4.251894,3.6857557,3.1235218,2.6510892,2.174752,1.698415,1.2259823,0.74964523,0.77307165,0.80040246,0.8238289,0.8511597,0.8745861,0.7262188,0.57394713,0.42557985,0.27330816,0.12494087,0.76135844,1.4016805,2.0380979,2.6745155,3.310933,8.488171,13.661504,18.838741,24.012074,29.189312,33.24989,37.310467,41.37495,45.439434,49.50001,47.33697,45.173935,43.010895,40.85176,38.68872,33.12495,27.561176,22.001307,16.437534,10.87376,12.70102,14.524376,16.351637,18.174992,19.998348,17.850927,15.699601,13.548276,11.400854,9.249529,7.601871,5.950309,4.298747,2.6510892,0.999527,3.4124475,5.825368,8.238289,10.651209,13.06413,12.025558,10.986988,9.948417,8.913751,7.8751793,7.125534,6.375889,5.6262436,4.8765984,4.123049,3.3616903,2.6003318,1.8389735,1.0737107,0.31235218,0.97610056,1.6359446,2.2996929,2.9634414,3.6232853,2.900971,2.174752,1.4485333,0.7262188,0.0,0.78868926,1.5734742,2.3621633,3.1508527,3.9356375,6.1611466,8.386656,10.612165,12.837675,15.063184,12.0606985,9.062118,6.0635366,3.0610514,0.062470436,0.10151446,0.13665408,0.1756981,0.21083772,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,2.4871042,4.911738,7.336372,9.761005,12.185639,13.013372,13.837202,14.661031,15.488764,16.312593,15.762072,15.211552,14.661031,14.114414,13.563893,12.27544,10.986988,9.698535,8.413987,7.125534,7.426173,7.726812,8.023546,8.324185,8.624825,7.137247,5.64967,4.1620927,2.6745155,1.1869383,1.4016805,1.6125181,1.8233559,2.0380979,2.2489357,2.2137961,2.174752,2.135708,2.1005683,2.0615244,1.6867018,1.3118792,0.93705654,0.5622339,0.18741131,0.41386664,0.63641757,0.8628729,1.0893283,1.3118792,2.77603,4.2362766,5.700427,7.1606736,8.624825,7.387129,6.1494336,4.911738,3.6740425,2.436347,2.4480603,2.463678,2.475391,2.4871042,2.4988174,1.999054,1.4992905,0.999527,0.4997635,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.5114767,1.0268579,1.5383345,2.0498111,2.5612879,2.1122816,1.6632754,1.2142692,0.76135844,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.19912452,0.39824903,0.60127795,0.80040246,0.999527,0.8628729,0.7262188,0.58566034,0.44900626,0.31235218,0.38653582,0.46071947,0.5388075,0.61299115,0.6871748,0.9878138,1.2884527,1.5890918,1.8858263,2.1864653,3.7482262,5.3138914,6.8756523,8.437413,9.999174,8.113348,6.223617,4.337791,2.4480603,0.5622339,1.1635119,1.7608855,2.3621633,2.9634414,3.5608149,2.8502135,2.135708,1.4251068,0.7106012,0.0,0.13665408,0.27330816,0.41386664,0.5505207,0.6871748,2.2255092,3.7638438,5.298274,6.8366084,8.374943,8.261715,8.148487,8.039165,7.9259367,7.812709,7.562827,7.3129454,7.0630636,6.813182,6.5633,5.4856853,4.4119744,3.338264,2.260649,1.1869383,1.9756275,2.7643168,3.5491016,4.337791,5.12648,5.4505453,5.774611,6.098676,6.426646,6.7507114,6.098676,5.4505453,4.7985106,4.1503797,3.4983444,4.337791,5.173333,6.012779,6.8483214,7.687768,6.1611466,4.6384296,3.1118085,1.5890918,0.062470436,1.8506867,3.638903,5.423215,7.211431,8.999647,7.6135845,6.223617,4.8375545,3.4514916,2.0615244,2.3855898,2.7135596,3.0376248,3.3616903,3.6857557,3.2992198,2.912684,2.5261483,2.135708,1.7491722,4.900025,8.050878,11.20173,14.348679,17.49953,16.211079,14.92653,13.638077,12.349625,11.061172,14.051944,17.03881,20.025679,23.012547,25.999414,28.900385,31.801357,34.69842,37.599392,40.500366,37.298756,34.101048,30.899439,27.701735,24.500124,26.311768,28.12341,29.938957,31.750599,33.56224,31.285975,29.013613,26.737347,24.46108,22.188719,21.575727,20.962736,20.349745,19.736753,19.123762,16.187653,13.251541,10.311526,7.375416,4.4393053,6.4891167,8.538928,10.588739,12.63855,14.688361,15.586374,16.48829,17.386303,18.28822,19.186234,15.500477,11.810817,8.125061,4.4393053,0.74964523,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,3.8380275,7.676055,11.514082,15.348206,19.186234,15.348206,11.514082,7.676055,3.8380275,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.0,0.0,0.0,0.0,0.0,1.0893283,2.174752,3.2640803,4.349504,5.4388323,4.376835,3.310933,2.2489357,1.1869383,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.7262188,1.3860629,2.0498111,2.7135596,3.3734035,5.349031,7.3246584,9.300286,11.275913,13.251541,10.71368,8.175818,5.6379566,3.1000953,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.9136301,1.5110037,2.1122816,2.7135596,3.310933,3.6623292,4.0137253,4.3612175,4.7126136,5.0640097,6.5008297,7.9376497,9.37447,10.81129,12.24811,11.986515,11.72492,11.4633255,11.20173,10.936231,9.550168,8.164105,6.774138,5.388075,3.998108,4.8883114,5.774611,6.66091,7.551114,8.437413,8.687295,8.937177,9.187058,9.43694,9.686822,8.449126,7.211431,5.9737353,4.73604,3.4983444,2.7994564,2.1005683,1.4016805,0.698888,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.3240654,0.46071947,0.60127795,0.737932,0.8745861,5.364649,9.850807,14.336966,18.823124,23.313187,19.998348,16.687416,13.376482,10.061645,6.7507114,5.3997884,4.0488653,2.7018464,1.3509232,0.0,0.4997635,0.999527,1.4992905,1.999054,2.4988174,2.3621633,2.2255092,2.0888553,1.9482968,1.8116426,2.8385005,3.8614538,4.8883114,5.911265,6.9381227,5.9737353,5.0132523,4.0488653,3.0883822,2.1239948,2.436347,2.7486992,3.0610514,3.3734035,3.6857557,3.9746814,4.263607,4.548629,4.8375545,5.12648,6.66091,8.1992445,9.737579,11.275913,12.814248,11.0260315,9.237816,7.4495993,5.661383,3.873167,4.126953,4.376835,4.6267166,4.8765984,5.12648,4.8492675,4.575959,4.298747,4.025439,3.7482262,3.4866312,3.2250361,2.9634414,2.7018464,2.436347,2.1630387,1.8858263,1.6125181,1.33921,1.0619974,1.2142692,1.3626363,1.5110037,1.6632754,1.8116426,2.2489357,2.6862288,3.1235218,3.5608149,3.998108,3.2640803,2.5261483,1.7882162,1.0502841,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,4.911738,5.036679,5.1616197,5.2865605,5.4115014,5.5364423,5.1108627,4.689187,4.263607,3.8380275,3.4124475,2.854118,2.2918842,1.7335546,1.1713207,0.61299115,0.97219616,1.3314011,1.6906061,2.0537157,2.4129205,1.9873407,1.5617609,1.1361811,0.7106012,0.28892577,1.1283722,1.9717231,2.815074,3.6584249,4.5017757,11.678067,18.854359,26.034554,33.210846,40.38714,43.799583,47.212032,50.62448,54.036926,57.449375,52.51421,47.57514,42.636074,37.70091,32.76184,27.96333,23.168722,18.370213,13.571702,8.773191,10.241247,11.705398,13.169549,14.633699,16.101755,14.532186,12.96652,11.39695,9.8312845,8.261715,7.137247,6.012779,4.8883114,3.7638438,2.639376,4.50568,6.3719845,8.238289,10.108498,11.974802,11.393045,10.81129,10.22563,9.643873,9.062118,8.492075,7.9220324,7.3519893,6.7819467,6.211904,5.263134,4.318269,3.3694992,2.4207294,1.475864,1.8194515,2.1591344,2.5027218,2.8463092,3.1859922,2.77603,2.3621633,1.9482968,1.5383345,1.1244678,1.5305257,1.9365835,2.338737,2.7447948,3.1508527,4.93126,6.7116675,8.488171,10.268578,12.0489855,9.651682,7.250475,4.8492675,2.4480603,0.05075723,0.14836729,0.24597734,0.3435874,0.44119745,0.5388075,0.5349031,0.5309987,0.5309987,0.5270943,0.5231899,2.416825,4.3065557,6.196286,8.086017,9.975748,10.67854,11.381332,12.084125,12.783013,13.4858055,13.58732,13.688834,13.786445,13.887959,13.985569,12.73616,11.482847,10.229534,8.976221,7.726812,7.6955767,7.6643414,7.633106,7.605776,7.57454,6.6531014,5.7316628,4.806319,3.8848803,2.9634414,3.0298162,3.096191,3.1664703,3.232845,3.2992198,3.0376248,2.77603,2.514435,2.2489357,1.9873407,1.893635,1.8038338,1.7101282,1.6164225,1.5266213,1.639849,1.7530766,1.8702087,1.9834363,2.1005683,3.4397783,4.7789884,6.1181984,7.461313,8.800523,8.445222,8.089922,7.734621,7.37932,7.0240197,6.1181984,5.2162814,4.31046,3.4046388,2.4988174,1.999054,1.4992905,0.999527,0.4997635,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.1717937,0.14055848,0.10932326,0.078088045,0.05075723,0.07027924,0.08980125,0.10932326,0.12884527,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.41777104,0.8355421,1.2533131,1.6710842,2.0888553,1.7843118,1.475864,1.1713207,0.8667773,0.5622339,0.48805028,0.41386664,0.3357786,0.26159495,0.18741131,0.5114767,0.8316377,1.1557031,1.475864,1.7999294,1.4914817,1.1791295,0.8706817,0.5583295,0.24988174,0.31235218,0.37482262,0.43729305,0.4997635,0.5622339,0.9956226,1.4290112,1.8584955,2.2918842,2.7252727,3.7794614,4.83365,5.891743,6.9459314,8.00012,6.5437784,5.0913405,3.6349986,2.1786566,0.7262188,1.1557031,1.5851873,2.0146716,2.4441557,2.87364,2.4012074,1.9287747,1.456342,0.98390937,0.5114767,0.5583295,0.60127795,0.6481308,0.6910792,0.737932,2.018576,3.2992198,4.575959,5.8566036,7.137247,7.1294384,7.1216297,7.113821,7.1060123,7.098203,6.7780423,6.453977,6.133816,5.8097506,5.4856853,4.8570766,4.2284675,3.5959544,2.9673457,2.338737,2.8619268,3.3812122,3.9044023,4.4275923,4.950782,5.185046,5.4193106,5.6535745,5.891743,6.126007,5.473972,4.8219366,4.165997,3.513962,2.8619268,3.521771,4.181615,4.841459,5.5013027,6.1611466,4.950782,3.736513,2.5261483,1.3118792,0.10151446,1.5461433,2.9907722,4.435401,5.8800297,7.3246584,6.375889,5.423215,4.474445,3.5256753,2.5769055,2.736986,2.900971,3.0610514,3.2250361,3.3890212,3.049338,2.7057507,2.366068,2.0263848,1.6867018,4.1777105,6.6687193,9.155824,11.6468315,14.13784,13.110983,12.08803,11.061172,10.0382185,9.01136,12.552653,16.093946,19.631334,23.172626,26.71392,28.80668,30.895535,32.988297,35.081055,37.173813,34.11667,31.055616,27.994564,24.933514,21.876366,22.946173,24.015978,25.085785,26.15559,27.225397,25.362997,23.504501,21.646006,19.783606,17.92511,17.468296,17.015385,16.55857,16.10566,15.648844,13.228115,10.81129,8.39056,5.969831,3.5491016,5.2084727,6.871748,8.531119,10.19049,11.849861,12.642454,13.435048,14.227642,15.020235,15.812829,13.435048,11.057267,8.679486,6.3017054,3.9239242,3.3031244,2.6862288,2.0654287,1.4446288,0.8238289,0.74574083,0.6715572,0.59346914,0.5153811,0.43729305,3.4202564,6.4032197,9.386183,12.369146,15.348206,12.306676,9.261242,6.2158084,3.1703746,0.12494087,0.359205,0.58956474,0.8238289,1.0541886,1.2884527,1.1205635,0.95267415,0.78478485,0.61689556,0.44900626,0.4958591,0.5466163,0.59346914,0.64032197,0.6871748,1.8389735,2.9868677,4.138666,5.2865605,6.4383593,5.4115014,4.380739,3.3538816,2.3270237,1.3001659,1.5110037,1.7218413,1.9287747,2.1396124,2.35045,2.6081407,2.8658314,3.1235218,3.3812122,3.638903,5.3295093,7.016211,8.706817,10.397423,12.08803,9.780528,7.47693,5.173333,2.8658314,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.30063897,0.60518235,0.9058213,1.2103647,1.5110037,2.2020829,2.893162,3.5842414,4.271416,4.9624953,5.267039,5.571582,5.8761253,6.180669,6.4891167,7.7814736,9.073831,10.366188,11.6585455,12.950902,12.341816,11.736633,11.127546,10.518459,9.913278,9.128492,8.347612,7.5667315,6.7819467,6.001066,6.590631,7.1841,7.7775693,8.371038,8.960603,9.198771,9.433036,9.6673,9.901564,10.135828,8.671678,7.2036223,5.735567,4.267512,2.7994564,2.241127,1.678893,1.1205635,0.5583295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.26159495,0.3709182,0.48024148,0.58956474,0.698888,4.298747,7.8947015,11.490656,15.090515,18.68647,16.863113,15.035853,13.212498,11.389141,9.561881,7.648724,5.7394714,3.8263142,1.9131571,0.0,0.4997635,0.999527,1.4992905,1.999054,2.4988174,2.8306916,3.1586614,3.4905357,3.8185053,4.1503797,4.73604,5.3217,5.903456,6.4891167,7.0747766,6.2587566,5.4388323,4.6228123,3.8067923,2.9868677,3.435874,3.8809757,4.3299823,4.7789884,5.22409,5.298274,5.368553,5.4427366,5.5169206,5.5871997,7.000593,8.413987,9.823476,11.23687,12.650263,11.084598,9.518932,7.9532676,6.3915067,4.825841,5.0054436,5.185046,5.364649,5.5442514,5.7238536,5.3412223,4.9546866,4.5681505,4.185519,3.7989833,3.7091823,3.619381,3.5295796,3.4397783,3.349977,2.9361105,2.5261483,2.1122816,1.698415,1.2884527,1.4094892,1.53443,1.6554666,1.7765031,1.901444,2.25284,2.6042364,2.9556324,3.310933,3.6623292,3.2289407,2.7916477,2.358259,1.9209659,1.4875772,1.2025559,0.91753453,0.63251317,0.3474918,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,6.8873653,6.5359693,6.1884775,5.8370814,5.4856853,5.138193,4.8492675,4.564246,4.2753205,3.9863946,3.7013733,3.0532427,2.4090161,1.7647898,1.1205635,0.47633708,1.1713207,1.8663043,2.5612879,3.2562714,3.951255,3.2484627,2.5495746,1.8506867,1.1517987,0.44900626,1.4992905,2.5456703,3.59205,4.6384296,5.688714,14.867964,24.047213,33.226463,42.40962,51.588867,54.34928,57.113598,59.87401,62.638325,65.398735,57.687542,49.97635,42.26125,34.550056,26.838861,22.805614,18.772366,14.739119,10.705871,6.676528,7.7814736,8.886419,9.991365,11.096312,12.201257,11.213444,10.229534,9.245625,8.261715,7.2739015,6.676528,6.0752497,5.473972,4.8765984,4.2753205,5.5989127,6.918601,8.242193,9.565785,10.889378,10.760532,10.631687,10.506746,10.377901,10.249056,9.858616,9.468176,9.081639,8.691199,8.300759,7.168483,6.036206,4.903929,3.7716527,2.639376,2.6588979,2.6823244,2.7057507,2.7291772,2.7486992,2.6510892,2.5495746,2.4480603,2.35045,2.2489357,2.2723622,2.2957885,2.3192148,2.338737,2.3621633,3.697469,5.0327744,6.36808,7.703386,9.0386915,7.238762,5.4388323,3.638903,1.8389735,0.039044023,0.19522011,0.3513962,0.5114767,0.6676528,0.8238289,0.8589685,0.8902037,0.92143893,0.95657855,0.9878138,2.3426414,3.697469,5.0522966,6.407124,7.7619514,8.343708,8.921559,9.503315,10.081166,10.662923,11.412568,12.162213,12.911859,13.661504,14.411149,13.196879,11.978706,10.760532,9.542359,8.324185,7.9649806,7.605776,7.2465706,6.883461,6.524256,6.168956,5.8097506,5.4505453,5.095245,4.73604,4.661856,4.5837684,4.50568,4.4275923,4.349504,3.8614538,3.3734035,2.8892577,2.4012074,1.9131571,2.1005683,2.2918842,2.4831998,2.6706111,2.8619268,2.8658314,2.87364,2.8775444,2.8814487,2.8892577,4.1035266,5.3217,6.5398736,7.758047,8.976221,9.503315,10.03041,10.557504,11.084598,11.611692,9.788337,7.968885,6.1455293,4.322173,2.4988174,1.999054,1.4992905,0.999527,0.4997635,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.12884527,0.10541886,0.08199245,0.058566034,0.039044023,0.05075723,0.06637484,0.08199245,0.09761006,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.3240654,0.6442264,0.96829176,1.2884527,1.6125181,1.4524376,1.2923572,1.1322767,0.97219616,0.81211567,0.7262188,0.63641757,0.5505207,0.46071947,0.37482262,0.8199245,1.2650263,1.7101282,2.15523,2.6003318,2.1161861,1.6359446,1.1517987,0.6715572,0.18741131,0.23816854,0.28892577,0.3357786,0.38653582,0.43729305,1.0034313,1.5656652,2.1318035,2.697942,3.2640803,3.8106966,4.357313,4.903929,5.4505453,6.001066,4.9781127,3.9551594,2.9322062,1.9092526,0.8862993,1.1478943,1.4055848,1.6671798,1.9287747,2.1864653,1.9561055,1.7218413,1.4914817,1.2572175,1.0268579,0.97610056,0.92924774,0.8823949,0.8355421,0.78868926,1.8116426,2.8306916,3.853645,4.8765984,5.899552,5.997162,6.094772,6.192382,6.289992,6.387602,5.9932575,5.5989127,5.2006636,4.806319,4.4119744,4.2284675,4.041056,3.8575494,3.6740425,3.4866312,3.7443218,4.0020123,4.2597027,4.5173936,4.775084,4.919547,5.0640097,5.2084727,5.35684,5.5013027,4.845363,4.1894236,3.533484,2.8814487,2.2255092,2.7057507,3.1898966,3.6740425,4.154284,4.6384296,3.736513,2.8385005,1.9365835,1.038571,0.13665408,1.2415999,2.3426414,3.4436827,4.548629,5.64967,5.138193,4.6267166,4.1113358,3.5998588,3.0883822,3.0883822,3.0883822,3.0883822,3.0883822,3.0883822,2.795552,2.5027218,2.2098918,1.9170616,1.6242313,3.455396,5.2865605,7.113821,8.944985,10.77615,10.010887,9.249529,8.488171,7.726812,6.9615493,11.053363,15.14908,19.240894,23.332708,27.424522,28.70907,29.993618,31.278166,32.56662,33.851166,30.930676,28.010181,25.08969,22.169195,19.248703,19.576674,19.904642,20.232613,20.560583,20.888552,19.443924,17.999294,16.55076,15.1061325,13.661504,13.364769,13.068034,12.771299,12.470661,12.173926,10.272482,8.371038,6.46569,4.564246,2.6628022,3.9317331,5.2006636,6.473499,7.7424297,9.01136,9.698535,10.381805,11.06898,11.752251,12.439425,11.369619,10.303718,9.2339115,8.16801,7.098203,5.985449,4.8687897,3.7560349,2.639376,1.5266213,1.3938715,1.2650263,1.1361811,1.0034313,0.8745861,3.0024853,5.1303844,7.2582836,9.386183,11.514082,9.261242,7.008402,4.755562,2.5027218,0.24988174,0.61689556,0.98000497,1.3431144,1.7101282,2.0732377,1.8389735,1.6047094,1.3704453,1.1361811,0.9019169,0.9956226,1.0893283,1.1869383,1.2806439,1.3743496,2.5886188,3.7989833,5.0132523,6.223617,7.437886,6.446168,5.45445,4.4588275,3.4671092,2.475391,2.9087796,3.338264,3.7716527,4.2050414,4.6384296,4.4900627,4.3416953,4.193328,4.0488653,3.900498,5.3060827,6.7116675,8.113348,9.518932,10.924518,8.85128,6.7819467,4.7087092,2.6354716,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.5427119,1.0854238,1.6281357,2.1708477,2.7135596,3.49444,4.271416,5.0522966,5.833177,6.6140575,6.871748,7.1333427,7.3910336,7.6526284,7.914223,9.058213,10.206107,11.354002,12.501896,13.64979,12.697116,11.744442,10.791768,9.839094,8.886419,8.710721,8.531119,8.355421,8.175818,8.00012,8.296855,8.59359,8.894228,9.190963,9.487698,9.706344,9.928895,10.147541,10.366188,10.588739,8.890324,7.191909,5.493494,3.7989833,2.1005683,1.678893,1.261122,0.8394465,0.42167544,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.19522011,0.27721256,0.359205,0.44119745,0.5231899,3.232845,5.938596,8.648251,11.354002,14.063657,13.723974,13.388195,13.048512,12.712734,12.376955,9.901564,7.426173,4.950782,2.475391,0.0,0.4997635,0.999527,1.4992905,1.999054,2.4988174,3.2992198,4.095718,4.892216,5.688714,6.4891167,6.6335793,6.7780423,6.9225054,7.066968,7.211431,6.5398736,5.8683167,5.196759,4.521298,3.8497405,4.4314966,5.0132523,5.5989127,6.180669,6.7624245,6.621866,6.477403,6.336845,6.192382,6.0518236,7.336372,8.624825,9.913278,11.20173,12.486279,11.143164,9.803954,8.460839,7.1177254,5.774611,5.883934,5.9932575,6.1064854,6.2158084,6.3251314,5.8292727,5.3334136,4.841459,4.3455997,3.8497405,3.9317331,4.0137253,4.095718,4.181615,4.263607,3.7130866,3.1625657,2.612045,2.0615244,1.5110037,1.6086137,1.7023194,1.796025,1.893635,1.9873407,2.2567444,2.522244,2.7916477,3.057147,3.3265507,3.193801,3.0610514,2.9283018,2.795552,2.6628022,2.1435168,1.6242313,1.1010414,0.58175594,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,8.862993,8.039165,7.211431,6.387602,5.563773,4.73604,4.5876727,4.4393053,4.2870336,4.138666,3.9863946,3.2562714,2.5261483,1.796025,1.0659018,0.3357786,1.3665408,2.397303,3.4280653,4.4588275,5.4856853,4.513489,3.5373883,2.5612879,1.5890918,0.61299115,1.8663043,3.1157131,4.369026,5.6223392,6.8756523,18.057861,29.240068,40.422276,51.604485,62.786694,64.89897,67.01125,69.123535,71.23582,73.3481,62.860878,52.373653,41.88643,31.399202,20.911978,17.643993,14.376009,11.108025,7.843944,4.575959,5.3217,6.0635366,6.8092775,7.5550184,8.300759,7.898606,7.4964523,7.094299,6.688241,6.2860875,6.211904,6.13772,6.0635366,5.989353,5.911265,6.688241,7.4691215,8.246098,9.023073,9.80005,10.128019,10.455989,10.783959,11.111929,11.435994,11.229061,11.018223,10.807385,10.596548,10.38571,9.069926,7.7541428,6.434455,5.1186714,3.7989833,3.5022488,3.2055142,2.9087796,2.6081407,2.3114061,2.5261483,2.736986,2.951728,3.1625657,3.3734035,3.0141985,2.6549935,2.2957885,1.9365835,1.5734742,2.463678,3.3538816,4.2440853,5.134289,6.0244927,4.825841,3.6232853,2.4246337,1.2259823,0.023426414,0.24207294,0.46071947,0.679366,0.8941081,1.1127546,1.1791295,1.2494087,1.3157835,1.3821584,1.4485333,2.2684577,3.0883822,3.9083066,4.728231,5.548156,6.008875,6.46569,6.9225054,7.37932,7.8361354,9.237816,10.6355915,12.037272,13.438952,14.836729,13.653695,12.470661,11.291532,10.108498,8.925464,8.234385,7.5433054,6.8561306,6.165051,5.473972,5.6809053,5.891743,6.098676,6.3056097,6.5125427,6.289992,6.067441,5.84489,5.6223392,5.3997884,4.689187,3.9746814,3.2640803,2.5495746,1.8389735,2.3114061,2.7838387,3.2562714,3.7287042,4.2011366,4.095718,3.9902992,3.8848803,3.7794614,3.6740425,4.7711797,5.8644123,6.9615493,8.054782,9.151918,10.561408,11.970898,13.380386,14.789876,16.199366,13.458474,10.721489,7.9805984,5.239708,2.4988174,1.999054,1.4992905,0.999527,0.4997635,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.08589685,0.07027924,0.05466163,0.039044023,0.023426414,0.03513962,0.046852827,0.05466163,0.06637484,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.22645533,0.45681506,0.6832704,0.9097257,1.1361811,1.1205635,1.1088502,1.0932326,1.077615,1.0619974,0.96438736,0.8628729,0.76135844,0.6637484,0.5622339,1.1283722,1.698415,2.2645533,2.8306916,3.4007344,2.7447948,2.0888553,1.43682,0.78088045,0.12494087,0.1639849,0.19912452,0.23816854,0.27330816,0.31235218,1.0112402,1.7062237,2.4051118,3.1039999,3.7989833,3.8419318,3.8809757,3.9200199,3.959064,3.998108,3.408543,2.8189783,2.2294137,1.639849,1.0502841,1.1400855,1.2298868,1.319688,1.4094892,1.4992905,1.5070993,1.5149081,1.5227169,1.5305257,1.5383345,1.397776,1.2572175,1.116659,0.97610056,0.8394465,1.6008049,2.366068,3.1313305,3.8965936,4.661856,4.8648853,5.067914,5.270943,5.473972,5.6730967,5.2084727,4.7399445,4.271416,3.8067923,3.338264,3.5959544,3.8575494,4.1191444,4.376835,4.6384296,4.630621,4.6228123,4.6150036,4.607195,4.5993857,4.6540475,4.7087092,4.7633705,4.8219366,4.8765984,4.2167544,3.5608149,2.900971,2.2450314,1.5890918,1.893635,2.1981785,2.5027218,2.8072653,3.1118085,2.5261483,1.9365835,1.3509232,0.76135844,0.1756981,0.93315214,1.6945106,2.455869,3.213323,3.9746814,3.900498,3.8263142,3.7482262,3.6740425,3.5998588,3.435874,3.2757936,3.1118085,2.951728,2.787743,2.541766,2.2957885,2.0537157,1.8077383,1.5617609,2.7330816,3.9044023,5.0718184,6.2431393,7.4144597,6.910792,6.4110284,5.911265,5.4115014,4.911738,9.557977,14.204215,18.84655,23.492788,28.139027,28.615364,29.091702,29.571943,30.048279,30.524616,27.744682,24.964748,22.184814,19.404879,16.624945,16.211079,15.793307,15.37944,14.965574,14.551707,13.520945,12.490183,11.45942,10.4286585,9.4018,9.261242,9.120684,8.980125,8.839567,8.699008,7.3168497,5.930787,4.5447245,3.1586614,1.7765031,2.6549935,3.533484,4.415879,5.2943697,6.1767645,6.7507114,7.328563,7.9064145,8.484266,9.062118,9.304191,9.546264,9.788337,10.034314,10.276386,8.663869,7.055255,5.446641,3.8341231,2.2255092,2.0420024,1.8584955,1.678893,1.4953861,1.3118792,2.5847144,3.8575494,5.1303844,6.4032197,7.676055,6.2158084,4.755562,3.2953155,1.8350691,0.37482262,0.8706817,1.3704453,1.8663043,2.366068,2.8619268,2.5612879,2.2567444,1.9561055,1.6515622,1.3509232,1.4914817,1.6359446,1.7765031,1.9209659,2.0615244,3.338264,4.6110992,5.8878384,7.1606736,8.437413,7.480835,6.524256,5.563773,4.607195,3.6506162,4.3065557,4.958591,5.6145306,6.27047,6.9264097,6.3719845,5.8214636,5.267039,4.716518,4.1620927,5.282656,6.4032197,7.523783,8.644346,9.761005,7.9220324,6.083059,4.2440853,2.4012074,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.78088045,1.5656652,2.3465457,3.1313305,3.912211,4.7828927,5.6535745,6.524256,7.3910336,8.261715,8.476458,8.691199,8.905942,9.120684,9.339331,10.338858,11.342289,12.34572,13.349152,14.348679,13.052417,11.756155,10.455989,9.159728,7.8634663,8.289046,8.718531,9.14411,9.573594,9.999174,10.003078,10.003078,10.006983,10.010887,10.010887,10.217821,10.42085,10.627783,10.8308115,11.037745,9.108971,7.1841,5.2553253,3.3265507,1.4016805,1.1205635,0.8394465,0.5583295,0.28111696,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.12884527,0.1835069,0.23816854,0.29673457,0.3513962,2.1669433,3.9863946,5.801942,7.621393,9.43694,10.588739,11.736633,12.888432,14.036326,15.188125,12.150499,9.112875,6.0752497,3.0376248,0.0,0.4997635,0.999527,1.4992905,1.999054,2.4988174,3.7638438,5.02887,6.2938967,7.558923,8.823949,8.531119,8.234385,7.941554,7.6448197,7.348085,6.8209906,6.2938967,5.7668023,5.239708,4.7126136,5.4310236,6.1455293,6.8639393,7.5823493,8.300759,7.941554,7.5862536,7.2270484,6.871748,6.5125427,7.676055,8.839567,9.999174,11.162686,12.326198,11.205634,10.085071,8.964508,7.843944,6.7233806,6.7663293,6.805373,6.844417,6.883461,6.9264097,6.321227,5.716045,5.1108627,4.50568,3.900498,4.154284,4.4119744,4.6657605,4.919547,5.173333,4.4861584,3.7989833,3.1118085,2.4246337,1.737459,1.8038338,1.8741131,1.9404879,2.0068626,2.0732377,2.2567444,2.4402514,2.6237583,2.803361,2.9868677,3.1586614,3.3265507,3.4983444,3.6662338,3.8380275,3.0805733,2.3270237,1.5734742,0.8160201,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,10.838621,9.538455,8.238289,6.9381227,5.6379566,4.337791,4.3260775,4.3143644,4.298747,4.2870336,4.2753205,3.4593005,2.6432803,1.8311646,1.0151446,0.19912452,1.5656652,2.9283018,4.2948427,5.661383,7.0240197,5.774611,4.5252023,3.2757936,2.0263848,0.77307165,2.233318,3.68966,5.1460023,6.606249,8.062591,21.247757,34.432922,47.61809,60.803257,73.98843,75.44867,76.91282,78.37697,79.83722,81.30137,68.03812,54.77486,41.511604,28.24835,14.989,12.486279,9.983557,7.480835,4.9781127,2.475391,2.8580225,3.2445583,3.631094,4.0137253,4.4002614,4.579864,4.759466,4.939069,5.1186714,5.298274,5.7511845,6.2001905,6.649197,7.098203,7.551114,7.7814736,8.015738,8.246098,8.480362,8.710721,9.495506,10.276386,11.061172,11.842052,12.626837,12.595602,12.564366,12.533132,12.5058,12.4745655,10.971371,9.468176,7.968885,6.46569,4.9624953,4.3455997,3.7287042,3.1118085,2.4910088,1.8741131,2.4012074,2.9243972,3.4514916,3.9746814,4.5017757,3.7560349,3.0141985,2.2723622,1.5305257,0.78868926,1.2337911,1.678893,2.1239948,2.5690966,3.0141985,2.4129205,1.8116426,1.2142692,0.61299115,0.011713207,0.28892577,0.5661383,0.8433509,1.1205635,1.4016805,1.5031948,1.6047094,1.7062237,1.8116426,1.9131571,2.1981785,2.4831998,2.7682211,3.0532427,3.338264,3.6740425,4.0059166,4.3416953,4.677474,5.0132523,7.0630636,9.112875,11.162686,13.212498,15.262308,14.114414,12.96652,11.818625,10.670732,9.526741,8.503788,7.4847393,6.46569,5.446641,4.423688,5.196759,5.969831,6.7429028,7.5159745,8.289046,7.918128,7.551114,7.1841,6.817086,6.4500723,5.5130157,4.575959,3.638903,2.7018464,1.7608855,2.5183394,3.2718892,4.029343,4.7828927,5.5364423,5.3217,5.1069584,4.892216,4.677474,4.462732,5.434928,6.407124,7.37932,8.351517,9.323712,11.615597,13.911386,16.20327,18.495153,20.787037,17.128613,13.4740925,9.815667,6.1572423,2.4988174,1.999054,1.4992905,0.999527,0.4997635,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.042948425,0.03513962,0.027330816,0.019522011,0.011713207,0.015617609,0.023426414,0.027330816,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.13274968,0.26549935,0.39824903,0.5309987,0.6637484,0.79259366,0.92143893,1.0541886,1.183034,1.3118792,1.1986516,1.0893283,0.97610056,0.8628729,0.74964523,1.4407244,2.1318035,2.8189783,3.5100577,4.2011366,3.3734035,2.5456703,1.717937,0.8902037,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,1.0190489,1.8467822,2.67842,3.506153,4.337791,3.8692627,3.4007344,2.9361105,2.4675822,1.999054,1.8428779,1.6867018,1.5266213,1.3704453,1.2142692,1.1322767,1.0541886,0.97219616,0.8941081,0.81211567,1.0580931,1.3079748,1.5539521,1.8038338,2.0498111,1.8194515,1.5851873,1.3509232,1.1205635,0.8862993,1.3938715,1.901444,2.4090161,2.9165885,3.4241607,3.7326086,4.041056,4.3455997,4.6540475,4.9624953,4.423688,3.8809757,3.3421683,2.803361,2.260649,2.9673457,3.6740425,4.376835,5.083532,5.786324,5.5169206,5.2436123,4.970304,4.6969957,4.423688,4.388548,4.3534083,4.318269,4.283129,4.251894,3.5881457,2.9283018,2.2684577,1.6086137,0.94876975,1.077615,1.2064602,1.3314011,1.4602464,1.5890918,1.3118792,1.038571,0.76135844,0.48805028,0.21083772,0.62860876,1.0463798,1.4641509,1.8819219,2.2996929,2.6628022,3.0259118,3.3890212,3.7482262,4.1113358,3.78727,3.4632049,3.1391394,2.8111696,2.4871042,2.2918842,2.0927596,1.893635,1.698415,1.4992905,2.0107672,2.5183394,3.0298162,3.541293,4.0488653,3.8106966,3.5764325,3.338264,3.1000953,2.8619268,8.058686,13.2554455,18.45611,23.652868,28.849628,28.521658,28.189785,27.861814,27.52994,27.198067,24.558691,21.919313,19.279938,16.640562,14.001186,12.841579,11.685876,10.526268,9.370565,8.210958,7.5979667,6.9810715,6.36808,5.7511845,5.138193,5.153811,5.173333,5.1889505,5.2084727,5.22409,4.357313,3.4905357,2.6237583,1.7530766,0.8862993,1.3782539,1.8663043,2.358259,2.8463092,3.338264,3.8067923,4.279225,4.747753,5.2162814,5.688714,7.238762,8.792714,10.346666,11.896713,13.450665,11.346193,9.24172,7.1333427,5.02887,2.9243972,2.690133,2.455869,2.2216048,1.9834363,1.7491722,2.1669433,2.5847144,3.0024853,3.4202564,3.8380275,3.1703746,2.5027218,1.8350691,1.1674163,0.4997635,1.1283722,1.7608855,2.3894942,3.018103,3.6506162,3.279698,2.9087796,2.541766,2.1708477,1.7999294,1.9912452,2.1786566,2.3699722,2.5612879,2.7486992,4.087909,5.423215,6.7624245,8.101635,9.43694,8.515501,7.5940623,6.6687193,5.74728,4.825841,5.704332,6.578918,7.4574084,8.335898,9.21439,8.253906,7.297328,6.3407493,5.3841705,4.423688,5.2592297,6.094772,6.930314,7.7658563,8.601398,6.9927845,5.3841705,3.775557,2.1708477,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,1.0229534,2.0459068,3.06886,4.0918136,5.1108627,6.0713453,7.0318284,7.9923115,8.952794,9.913278,10.081166,10.25296,10.42085,10.592644,10.764437,11.619501,12.47847,13.333533,14.192502,15.051471,13.407718,11.763964,10.124115,8.480362,6.8366084,7.871275,8.902037,9.936704,10.967466,11.998228,11.709302,11.416472,11.123642,10.8308115,10.537982,10.729298,10.916709,11.108025,11.29934,11.486752,9.331521,7.172387,5.0132523,2.8580225,0.698888,0.5583295,0.42167544,0.28111696,0.14055848,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.06637484,0.093705654,0.12103647,0.14836729,0.1756981,1.1010414,2.0302892,2.9556324,3.8848803,4.814128,7.4495993,10.088976,12.724447,15.363823,17.999294,14.399435,10.799577,7.1997175,3.5998588,0.0,0.4997635,0.999527,1.4992905,1.999054,2.4988174,4.2323723,5.9659266,7.699481,9.4291315,11.162686,10.4286585,9.690726,8.956698,8.2226715,7.4886436,7.1060123,6.7233806,6.3407493,5.958118,5.575486,6.426646,7.28171,8.13287,8.98403,9.839094,9.265146,8.691199,8.121157,7.5472097,6.9732623,8.011833,9.050405,10.088976,11.123642,12.162213,11.2642,10.366188,9.468176,8.574067,7.676055,7.6448197,7.6135845,7.5862536,7.5550184,7.523783,6.8092775,6.094772,5.380266,4.6657605,3.951255,4.376835,4.806319,5.2318993,5.661383,6.086963,5.263134,4.4393053,3.611572,2.787743,1.9639144,2.0029583,2.0420024,2.0810463,2.1239948,2.1630387,2.260649,2.358259,2.455869,2.5534792,2.6510892,3.1235218,3.5959544,4.068387,4.5408196,5.0132523,4.0215344,3.0337205,2.0420024,1.0541886,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,12.814248,11.037745,9.261242,7.4886436,5.7121406,3.9356375,4.0605783,4.1894236,4.3143644,4.4393053,4.564246,3.6623292,2.7643168,1.8623998,0.96438736,0.062470436,1.7608855,3.4632049,5.1616197,6.8639393,8.562354,7.0357327,5.5130157,3.9863946,2.463678,0.93705654,2.6003318,4.263607,5.9268827,7.5862536,9.249529,24.437654,39.62578,54.813904,70.00203,85.18625,85.99837,86.814384,87.6265,88.438614,89.25073,73.21145,57.176067,41.136784,25.101402,9.062118,7.3246584,5.5871997,3.8497405,2.1122816,0.37482262,0.39824903,0.42557985,0.44900626,0.47633708,0.4997635,1.261122,2.0263848,2.787743,3.5491016,4.3143644,5.2865605,6.262661,7.238762,8.210958,9.187058,8.874706,8.562354,8.250002,7.9376497,7.6252975,8.862993,10.100689,11.338385,12.576079,13.813775,13.962143,14.114414,14.262781,14.411149,14.56342,12.8767185,11.186112,9.499411,7.812709,6.126007,5.1889505,4.251894,3.310933,2.3738766,1.43682,2.2762666,3.1118085,3.951255,4.786797,5.6262436,4.5017757,3.3734035,2.2489357,1.1244678,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3357786,0.6754616,1.0112402,1.3509232,1.6867018,1.8233559,1.9639144,2.1005683,2.2372224,2.3738766,2.1239948,1.8741131,1.6242313,1.3743496,1.1244678,1.33921,1.5500476,1.7608855,1.9756275,2.1864653,4.8883114,7.5862536,10.2881,12.986042,15.687888,14.575133,13.462379,12.349625,11.23687,10.124115,8.773191,7.426173,6.0752497,4.7243266,3.3734035,4.7126136,6.0518236,7.387129,8.726339,10.061645,9.550168,9.0386915,8.52331,8.011833,7.5003567,6.336845,5.173333,4.0137253,2.8502135,1.6867018,2.7252727,3.7638438,4.7985106,5.8370814,6.8756523,6.551587,6.223617,5.899552,5.575486,5.251421,6.098676,6.949836,7.800996,8.648251,9.499411,12.67369,15.847969,19.026152,22.200432,25.37471,20.79875,16.226696,11.650736,7.0747766,2.4988174,1.999054,1.4992905,0.999527,0.4997635,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.46071947,0.737932,1.0112402,1.2884527,1.5617609,1.43682,1.3118792,1.1869383,1.0619974,0.93705654,1.7491722,2.5612879,3.3734035,4.1894236,5.001539,3.998108,2.998581,1.999054,0.999527,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,1.0268579,1.9873407,2.951728,3.912211,4.8765984,3.900498,2.9243972,1.9482968,0.97610056,0.0,0.27330816,0.5505207,0.8238289,1.1010414,1.3743496,1.1244678,0.8745861,0.62470436,0.37482262,0.12494087,0.61299115,1.1010414,1.5890918,2.0732377,2.5612879,2.2372224,1.9131571,1.5890918,1.261122,0.93705654,1.1869383,1.43682,1.6867018,1.9365835,2.1864653,2.6003318,3.0141985,3.4241607,3.8380275,4.251894,3.638903,3.0259118,2.4129205,1.7999294,1.1869383,2.338737,3.4866312,4.6384296,5.786324,6.9381227,6.3993154,5.8644123,5.3256044,4.786797,4.251894,4.126953,3.998108,3.873167,3.7482262,3.6232853,2.9634414,2.2996929,1.6359446,0.97610056,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.10151446,0.13665408,0.1756981,0.21083772,0.24988174,0.3240654,0.39824903,0.47633708,0.5505207,0.62470436,1.4251068,2.2255092,3.0259118,3.8263142,4.6267166,4.138666,3.6506162,3.1625657,2.6745155,2.1864653,2.0380979,1.8858263,1.737459,1.5890918,1.43682,1.2884527,1.1361811,0.9878138,0.8394465,0.6871748,0.7106012,0.737932,0.76135844,0.78868926,0.81211567,6.5633,12.31058,18.061766,23.81295,29.564135,28.42405,27.287867,26.151686,25.0116,23.87542,21.376602,18.87388,16.375063,13.8762455,11.373524,9.475985,7.57454,5.6730967,3.775557,1.8741131,1.6749885,1.475864,1.2767396,1.0737107,0.8745861,1.0502841,1.2259823,1.4016805,1.5734742,1.7491722,1.4016805,1.0502841,0.698888,0.3513962,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.8628729,1.2259823,1.5890918,1.9482968,2.3114061,5.173333,8.039165,10.901091,13.763018,16.624945,14.024612,11.424281,8.823949,6.223617,3.6232853,3.338264,3.049338,2.7643168,2.475391,2.1864653,1.7491722,1.3118792,0.8745861,0.43729305,0.0,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,1.3860629,2.1513257,2.912684,3.6740425,4.4393053,3.998108,3.5608149,3.1235218,2.6862288,2.2489357,2.4871042,2.7252727,2.9634414,3.2016098,3.435874,4.8375545,6.239235,7.6370106,9.0386915,10.436467,9.550168,8.663869,7.773665,6.8873653,6.001066,7.098203,8.1992445,9.300286,10.401327,11.498465,10.135828,8.773191,7.4105554,6.0518236,4.689187,5.2358036,5.786324,6.336845,6.8873653,7.437886,6.0635366,4.689187,3.310933,1.9365835,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,1.261122,2.5261483,3.78727,5.0483923,6.3134184,7.363703,8.413987,9.464272,10.510651,11.560935,11.685876,11.810817,11.935758,12.0606985,12.185639,12.900145,13.610746,14.325252,15.035853,15.750359,13.763018,11.775677,9.788337,7.800996,5.813655,7.4495993,9.085544,10.725393,12.361338,14.001186,13.411622,12.825961,12.236397,11.650736,11.061172,11.23687,11.412568,11.588266,11.763964,11.935758,9.550168,7.1606736,4.775084,2.3855898,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,4.3143644,8.437413,12.564366,16.687416,20.81437,16.64837,12.486279,8.324185,4.1620927,0.0,0.4997635,0.999527,1.4992905,1.999054,2.4988174,4.7009,6.899079,9.101162,11.29934,13.501423,12.326198,11.150972,9.975748,8.800523,7.6252975,7.387129,7.1489606,6.910792,6.676528,6.4383593,7.426173,8.413987,9.4018,10.38571,11.373524,10.588739,9.80005,9.01136,8.226576,7.437886,8.351517,9.261242,10.174872,11.088503,11.998228,11.326671,10.651209,9.975748,9.300286,8.624825,8.52331,8.4257,8.324185,8.226576,8.125061,7.3012323,6.473499,5.64967,4.825841,3.998108,4.5993857,5.2006636,5.801942,6.3993154,7.000593,6.036206,5.0757227,4.1113358,3.1508527,2.1864653,2.1981785,2.2137961,2.2255092,2.2372224,2.2489357,2.260649,2.2762666,2.2879796,2.2996929,2.3114061,3.0883822,3.8614538,4.6384296,5.4115014,6.1884775,4.9624953,3.736513,2.5105307,1.2884527,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,10.986988,9.460366,7.9337454,6.4032197,4.8765984,3.349977,3.408543,3.4710135,3.5295796,3.5881457,3.6506162,3.377308,3.1039999,2.8306916,2.5612879,2.2879796,3.2484627,4.2089458,5.169429,6.126007,7.08649,5.872221,4.657952,3.4436827,2.2294137,1.0112402,3.2757936,5.5364423,7.800996,10.061645,12.326198,24.78124,37.24019,49.699135,62.15418,74.61313,74.605316,74.59751,74.5897,74.581894,74.57408,61.334255,48.094425,34.8546,21.61477,8.374943,7.191909,6.0049706,4.8219366,3.6349986,2.4519646,2.7486992,3.0454338,3.3421683,3.638903,3.9356375,4.2011366,4.466636,4.732136,4.997635,5.263134,5.7902284,6.3173227,6.844417,7.3715115,7.898606,7.7307167,7.5667315,7.3988423,7.230953,7.0630636,7.9532676,8.847376,9.741484,10.631687,11.525795,11.752251,11.978706,12.209065,12.435521,12.661977,11.701493,10.741011,9.780528,8.823949,7.8634663,6.551587,5.2436123,3.9317331,2.6237583,1.3118792,2.0224805,2.7330816,3.4436827,4.154284,4.860981,4.142571,3.4241607,2.7018464,1.9834363,1.261122,1.038571,0.81211567,0.58566034,0.3631094,0.13665408,0.30454338,0.47243267,0.64032197,0.80821127,0.97610056,1.1283722,1.2845483,1.4407244,1.5969005,1.7491722,2.2137961,2.67842,3.1469483,3.611572,4.0761957,4.3338866,4.5954814,4.853172,5.114767,5.376362,5.192855,5.009348,4.825841,4.646239,4.462732,6.329036,8.1992445,10.065549,11.931853,13.798158,12.771299,11.744442,10.717585,9.690726,8.663869,7.480835,6.297801,5.114767,3.9317331,2.7486992,3.8185053,4.884407,5.9542136,7.0201154,8.086017,7.676055,7.266093,6.8561306,6.446168,6.036206,5.1030536,4.165997,3.232845,2.2957885,1.3626363,2.241127,3.1235218,4.0020123,4.884407,5.7628975,5.45445,5.1460023,4.841459,4.533011,4.224563,4.903929,5.5832953,6.266566,6.9459314,7.6252975,10.666827,13.708356,16.75379,19.795319,22.83685,18.95197,15.067088,11.182208,7.297328,3.4124475,2.822883,2.233318,1.6437533,1.0541886,0.46071947,0.42948425,0.39824903,0.3631094,0.3318742,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.031235218,0.06637484,0.09761006,0.12884527,0.1639849,0.37872702,0.59737355,0.8160201,1.0307622,1.2494087,1.1517987,1.0502841,0.94876975,0.8511597,0.74964523,1.4016805,2.0498111,2.7018464,3.349977,3.998108,3.2016098,2.4012074,1.6008049,0.80040246,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.8199245,1.5890918,2.358259,3.1313305,3.900498,3.1235218,2.35045,1.5734742,0.80040246,0.023426414,0.23816854,0.45681506,0.6715572,0.8862993,1.1010414,0.9019169,0.698888,0.4997635,0.30063897,0.10151446,0.4958591,0.8902037,1.2845483,1.678893,2.0732377,1.9209659,1.7686942,1.6164225,1.4641509,1.3118792,1.4016805,1.4914817,1.5812829,1.6710842,1.7608855,2.1396124,2.5183394,2.893162,3.2718892,3.6506162,3.1313305,2.6159496,2.096664,1.5812829,1.0619974,1.9717231,2.8775444,3.7833657,4.6930914,5.5989127,5.165524,4.728231,4.2948427,3.8614538,3.4241607,3.3460727,3.2640803,3.1859922,3.1039999,3.0259118,2.7213683,2.4207294,2.1161861,1.815547,1.5110037,1.2259823,0.94096094,0.6559396,0.3709182,0.08589685,0.15227169,0.21864653,0.28111696,0.3474918,0.41386664,0.4958591,0.57785153,0.659844,0.7418364,0.8238289,1.5578566,2.2918842,3.0220075,3.7560349,4.4861584,4.173806,3.8614538,3.5491016,3.2367494,2.9243972,2.7291772,2.533957,2.338737,2.1435168,1.9482968,1.678893,1.4094892,1.1400855,0.8706817,0.60127795,0.71841,0.8355421,0.95267415,1.0698062,1.1869383,5.9737353,10.760532,15.551234,20.338032,25.124828,24.148727,23.168722,22.192623,21.216522,20.236517,18.081287,15.926057,13.770826,11.615597,9.464272,7.871275,6.278279,4.6852827,3.0922866,1.4992905,1.33921,1.1791295,1.0190489,0.8589685,0.698888,0.8433509,0.9917182,1.1361811,1.2806439,1.4251068,1.43682,1.4446288,1.456342,1.4641509,1.475864,1.3157835,1.1596074,1.0034313,0.8433509,0.6871748,1.5461433,2.4012074,3.260176,4.1191444,4.9742084,6.699954,8.4257,10.151445,11.873287,13.599033,12.271536,10.944039,9.616543,8.289046,6.9615493,7.098203,7.238762,7.375416,7.5120697,7.648724,6.9264097,6.2001905,5.473972,4.7516575,4.025439,3.8185053,3.6154766,3.408543,3.2055142,2.998581,4.123049,5.2436123,6.36808,7.4886436,8.6131115,7.715099,6.817086,5.919074,5.0210614,4.126953,4.318269,4.5095844,4.7009,4.8961205,5.087436,6.1572423,7.2270484,8.296855,9.366661,10.436467,9.788337,9.14411,8.495979,7.8478484,7.1997175,8.027451,8.855185,9.682918,10.510651,11.338385,10.0147915,8.691199,7.3715115,6.0479193,4.7243266,5.0718184,5.4193106,5.7668023,6.114294,6.461786,5.349031,4.2323723,3.1157131,2.0029583,0.8862993,0.8238289,0.75745404,0.6910792,0.62860876,0.5622339,1.6867018,2.8072653,3.9317331,5.0522966,6.1767645,7.211431,8.250002,9.288573,10.323239,11.361811,11.174399,10.986988,10.799577,10.612165,10.424754,11.326671,12.224684,13.1266,14.024612,14.92653,13.302299,11.681972,10.05774,8.433509,6.813182,7.996216,9.183154,10.366188,11.553126,12.73616,12.677594,12.619028,12.556558,12.497992,12.439425,11.869383,11.29934,10.729298,10.159255,9.589212,7.6682463,5.7511845,3.8341231,1.9170616,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,3.4983444,6.8483214,10.198298,13.548276,16.898252,13.520945,10.139732,6.75852,3.3812122,0.0,0.43729305,0.8745861,1.3118792,1.7491722,2.1864653,4.4002614,6.6140575,8.823949,11.037745,13.251541,11.873287,10.495033,9.116779,7.7385254,6.364176,6.844417,7.320754,7.800996,8.281238,8.761478,9.714153,10.662923,11.611692,12.564366,13.513136,12.888432,12.267632,11.6468315,11.022127,10.401327,10.967466,11.533605,12.103647,12.6697855,13.235924,12.743969,12.24811,11.752251,11.256392,10.764437,10.6590185,10.557504,10.455989,10.354475,10.249056,9.226103,8.203149,7.1841,6.1611466,5.138193,5.6262436,6.1181984,6.606249,7.098203,7.5862536,6.4695945,5.3529353,4.2362766,3.1157131,1.999054,2.0498111,2.1005683,2.1513257,2.1981785,2.2489357,2.25284,2.2567444,2.2567444,2.260649,2.260649,3.2016098,4.138666,5.0757227,6.012779,6.949836,5.6145306,4.279225,2.9439192,1.6086137,0.27330816,0.23426414,0.19131571,0.14836729,0.10541886,0.062470436,9.163632,7.882988,6.602344,5.3217,4.041056,2.7643168,2.7565079,2.7526035,2.7486992,2.7408905,2.736986,3.0922866,3.4475873,3.802888,4.1581883,4.513489,4.732136,4.950782,5.173333,5.3919797,5.610626,4.7087092,3.802888,2.8970666,1.9912452,1.0893283,3.951255,6.813182,9.675109,12.537036,15.398962,25.128733,34.8546,44.58437,54.310234,64.0361,63.208366,62.380634,61.556805,60.729073,59.90134,49.45706,39.016693,28.572416,18.12814,7.687768,7.055255,6.422742,5.7902284,5.1577153,4.5252023,5.095245,5.6652875,6.2353306,6.805373,7.375416,7.141152,6.910792,6.676528,6.446168,6.211904,6.2938967,6.3719845,6.453977,6.532065,6.6140575,6.590631,6.5672045,6.5437784,6.524256,6.5008297,7.0474463,7.5940623,8.140678,8.691199,9.237816,9.542359,9.846903,10.151445,10.455989,10.764437,10.530173,10.295909,10.065549,9.8312845,9.600925,7.918128,6.2353306,4.552533,2.8697357,1.1869383,1.7686942,2.3543546,2.9361105,3.5178664,4.0996222,3.7833657,3.4710135,3.154757,2.8385005,2.5261483,2.0732377,1.6242313,1.175225,0.7262188,0.27330816,0.60908675,0.94486535,1.2806439,1.6164225,1.9482968,1.9209659,1.893635,1.8663043,1.8389735,1.8116426,2.6042364,3.39683,4.1894236,4.9820175,5.774611,6.5437784,7.3168497,8.086017,8.855185,9.6243515,9.0465,8.468649,7.890797,7.3168497,6.7389984,7.773665,8.8083315,9.8429985,10.877665,11.912332,10.971371,10.0265045,9.085544,8.140678,7.1997175,6.184573,5.169429,4.154284,3.1391394,2.1239948,2.9243972,3.7208953,4.5173936,5.3138914,6.114294,5.805846,5.4973984,5.1889505,4.884407,4.575959,3.8692627,3.1586614,2.4519646,1.7452679,1.038571,1.7608855,2.4831998,3.2055142,3.9278288,4.650143,4.3612175,4.068387,3.7794614,3.4905357,3.2016098,3.7091823,4.220659,4.728231,5.239708,5.7511845,8.659965,11.568744,14.481428,17.390207,20.298986,17.105186,13.911386,10.71368,7.519879,4.3260775,3.6467118,2.9634414,2.2840753,1.6047094,0.92534333,0.8589685,0.79649806,0.7301232,0.6637484,0.60127795,0.48024148,0.359205,0.23816854,0.12103647,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.29673457,0.45681506,0.61689556,0.77697605,0.93705654,0.8628729,0.78868926,0.7106012,0.63641757,0.5622339,1.0502841,1.5383345,2.0263848,2.514435,2.998581,2.4012074,1.7999294,1.1986516,0.60127795,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.61689556,1.1908426,1.7686942,2.3465457,2.9243972,2.35045,1.7765031,1.1986516,0.62470436,0.05075723,0.20693332,0.359205,0.5153811,0.6715572,0.8238289,0.6754616,0.5231899,0.37482262,0.22645533,0.07418364,0.37872702,0.679366,0.98390937,1.2845483,1.5890918,1.6086137,1.6281357,1.6476578,1.6671798,1.6867018,1.6164225,1.5461433,1.475864,1.4055848,1.33921,1.678893,2.0224805,2.366068,2.7057507,3.049338,2.6276627,2.2059872,1.7843118,1.358732,0.93705654,1.6008049,2.2684577,2.9322062,3.5959544,4.263607,3.9317331,3.5959544,3.2640803,2.9322062,2.6003318,2.5651922,2.5300527,2.494913,2.4597735,2.4246337,2.4831998,2.541766,2.5964274,2.6549935,2.7135596,2.194274,1.6710842,1.1517987,0.63251317,0.113227665,0.20693332,0.29673457,0.39044023,0.48414588,0.57394713,0.6637484,0.75354964,0.8433509,0.93315214,1.0268579,1.6906061,2.3543546,3.018103,3.6857557,4.349504,4.21285,4.0761957,3.9356375,3.7989833,3.6623292,3.4241607,3.182088,2.9439192,2.7018464,2.463678,2.0732377,1.6827974,1.2923572,0.9019169,0.5114767,0.7223144,0.93315214,1.1439898,1.3509232,1.5617609,5.388075,9.2104845,13.036799,16.863113,20.685524,19.869503,19.053482,18.233559,17.417538,16.601519,14.789876,12.978233,11.170495,9.358852,7.551114,6.266566,4.9781127,3.6935644,2.4090161,1.1244678,1.0034313,0.8862993,0.76526284,0.6442264,0.5231899,0.64032197,0.75354964,0.8706817,0.98390937,1.1010414,1.4719596,1.8389735,2.2098918,2.5808098,2.951728,2.533957,2.1200905,1.7062237,1.2884527,0.8745861,2.2294137,3.5803368,4.93126,6.2860875,7.6370106,8.226576,8.812236,9.4018,9.987461,10.573121,10.518459,10.4637985,10.409137,10.354475,10.299813,10.862047,11.424281,11.986515,12.548749,13.110983,12.099743,11.088503,10.073358,9.062118,8.050878,7.5159745,6.9810715,6.446168,5.911265,5.376362,6.8561306,8.339804,9.823476,11.303245,12.786918,11.428185,10.073358,8.714626,7.355894,6.001066,6.1494336,6.2938967,6.4422636,6.590631,6.7389984,7.47693,8.218767,8.956698,9.698535,10.436467,10.03041,9.6243515,9.21439,8.8083315,8.398369,8.956698,9.511124,10.065549,10.619974,11.174399,9.893755,8.609207,7.328563,6.044015,4.7633705,4.9078336,5.0522966,5.196759,5.3412223,5.4856853,4.630621,3.7794614,2.9243972,2.069333,1.2142692,1.1947471,1.1791295,1.1596074,1.1439898,1.1244678,2.1083772,3.0883822,4.0722914,5.056201,6.036206,7.0630636,8.086017,9.112875,10.135828,11.162686,10.662923,10.163159,9.663396,9.163632,8.663869,9.749292,10.838621,11.924045,13.013372,14.098797,12.841579,11.584361,10.327144,9.069926,7.812709,8.546737,9.276859,10.010887,10.741011,11.475039,11.943566,12.408191,12.8767185,13.345247,13.813775,12.497992,11.182208,9.866425,8.550641,7.238762,5.7902284,4.3416953,2.893162,1.4485333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,2.6862288,5.263134,7.8361354,10.413041,12.986042,10.389614,7.793187,5.196759,2.5964274,0.0,0.37482262,0.74964523,1.1244678,1.4992905,1.8741131,4.0996222,6.3251314,8.550641,10.77615,13.001659,11.420377,9.839094,8.261715,6.6804323,5.099149,6.297801,7.4964523,8.691199,9.889851,11.088503,11.998228,12.911859,13.825488,14.739119,15.648844,15.192029,14.735214,14.278399,13.821584,13.360865,13.583415,13.805966,14.028518,14.251068,14.473619,14.161267,13.845011,13.528754,13.216402,12.900145,12.794726,12.689307,12.583888,12.47847,12.376955,11.154878,9.936704,8.714626,7.4964523,6.2743745,6.6531014,7.0357327,7.4144597,7.793187,8.175818,6.902983,5.630148,4.357313,3.084478,1.8116426,1.901444,1.9873407,2.0732377,2.1630387,2.2489357,2.241127,2.233318,2.2294137,2.2216048,2.2137961,3.310933,4.4119744,5.5130157,6.6140575,7.7111945,6.266566,4.8219366,3.377308,1.9326792,0.48805028,0.40215343,0.31625658,0.23426414,0.14836729,0.062470436,7.336372,6.3056097,5.270943,4.240181,3.2094188,2.174752,2.1044729,2.0341935,1.9639144,1.893635,1.8233559,2.8072653,3.7911747,4.7711797,5.755089,6.7389984,6.2158084,5.6965227,5.1772375,4.657952,4.138666,3.541293,2.9478238,2.3543546,1.756981,1.1635119,4.6267166,8.086017,11.549222,15.012426,18.475632,25.47232,32.46901,39.4696,46.46629,53.46298,51.815323,50.167664,48.520008,46.87235,45.22469,37.579872,29.935053,22.290232,14.645412,7.000593,6.918601,6.8405128,6.75852,6.6804323,6.5984397,7.4417906,8.285142,9.128492,9.971844,10.81129,10.081166,9.351044,8.62092,7.890797,7.1606736,6.79366,6.426646,6.0596323,5.6926184,5.3256044,5.446641,5.571582,5.6926184,5.813655,5.938596,6.141625,6.3407493,6.5437784,6.746807,6.949836,7.3324676,7.715099,8.097731,8.480362,8.862993,9.358852,9.850807,10.346666,10.8425255,11.338385,9.280765,7.2270484,5.173333,3.1157131,1.0619974,1.5188124,1.9717231,2.4285383,2.8814487,3.338264,3.4280653,3.5178664,3.6076677,3.697469,3.78727,3.1118085,2.436347,1.7608855,1.0893283,0.41386664,0.9136301,1.4172981,1.9209659,2.4207294,2.9243972,2.7135596,2.5066261,2.2957885,2.084951,1.8741131,2.9946766,4.11524,5.2358036,6.356367,7.47693,8.75367,10.034314,11.314958,12.595602,13.8762455,12.90405,11.931853,10.955752,9.983557,9.01136,9.21439,9.4174185,9.620447,9.823476,10.0265045,9.167537,8.308568,7.453504,6.5945354,5.735567,4.8883114,4.041056,3.193801,2.3465457,1.4992905,2.0263848,2.5534792,3.084478,3.611572,4.138666,3.9317331,3.7287042,3.521771,3.3187418,3.1118085,2.631567,2.1513257,1.6710842,1.1908426,0.7106012,1.2767396,1.8428779,2.4090161,2.97125,3.5373883,3.2640803,2.9907722,2.7213683,2.4480603,2.174752,2.514435,2.854118,3.193801,3.533484,3.873167,6.6531014,9.4291315,12.209065,14.985096,17.761126,15.258404,12.751778,10.249056,7.7424297,5.2358036,4.466636,3.697469,2.9283018,2.1591344,1.3860629,1.2884527,1.1908426,1.0932326,0.9956226,0.9019169,0.71841,0.5388075,0.359205,0.1796025,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.21474212,0.31625658,0.42167544,0.5231899,0.62470436,0.57394713,0.5231899,0.47633708,0.42557985,0.37482262,0.698888,1.0268579,1.3509232,1.6749885,1.999054,1.6008049,1.1986516,0.80040246,0.39824903,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.40996224,0.79649806,1.1791295,1.5656652,1.9482968,1.5734742,1.1986516,0.8238289,0.44900626,0.07418364,0.1717937,0.26549935,0.359205,0.45681506,0.5505207,0.44900626,0.3513962,0.24988174,0.14836729,0.05075723,0.26159495,0.46852827,0.679366,0.8902037,1.1010414,1.2923572,1.4836729,1.678893,1.8702087,2.0615244,1.8311646,1.6008049,1.3743496,1.1439898,0.9136301,1.2181735,1.5266213,1.8350691,2.1435168,2.4480603,2.1239948,1.796025,1.4680552,1.1400855,0.81211567,1.2337911,1.6593709,2.0810463,2.5027218,2.9243972,2.6940374,2.463678,2.233318,2.0068626,1.7765031,1.7843118,1.796025,1.8038338,1.815547,1.8233559,2.241127,2.6588979,3.076669,3.49444,3.912211,3.1586614,2.4012074,1.6476578,0.8941081,0.13665408,0.25769055,0.37872702,0.4958591,0.61689556,0.737932,0.8355421,0.93315214,1.0307622,1.1283722,1.2259823,1.8233559,2.4207294,3.018103,3.6154766,4.21285,4.251894,4.2870336,4.3260775,4.3612175,4.4002614,4.11524,3.8302186,3.5451972,3.260176,2.9751544,2.463678,1.9561055,1.4446288,0.93315214,0.42557985,0.7262188,1.0307622,1.3314011,1.6359446,1.9365835,4.7985106,7.6643414,10.526268,13.388195,16.250122,15.594183,14.934339,14.278399,13.618555,12.962616,11.498465,10.034314,8.566258,7.1021075,5.6379566,4.661856,3.6818514,2.7057507,1.7257458,0.74964523,0.6715572,0.58956474,0.5114767,0.42948425,0.3513962,0.43338865,0.5192855,0.60518235,0.6910792,0.77307165,1.5031948,2.233318,2.9634414,3.6935644,4.423688,3.7521305,3.0805733,2.4090161,1.7335546,1.0619974,2.9087796,4.755562,6.606249,8.453031,10.299813,9.749292,9.198771,8.648251,8.101635,7.551114,8.769287,9.983557,11.20173,12.419904,13.638077,14.625891,15.613705,16.601519,17.589333,18.573242,17.273075,15.976814,14.676648,13.376482,12.076316,11.209538,10.346666,9.479889,8.6131115,7.7502384,9.593117,11.435994,13.2788725,15.12175,16.960724,15.145176,13.325725,11.510178,9.690726,7.8751793,7.9766936,8.078208,8.183627,8.285142,8.386656,8.796618,9.20658,9.616543,10.0265045,10.436467,10.268578,10.100689,9.936704,9.768814,9.600925,9.882042,10.163159,10.44818,10.729298,11.014318,9.768814,8.527214,7.2856145,6.044015,4.7985106,4.743849,4.6852827,4.6267166,4.5681505,4.513489,3.9161155,3.3226464,2.7291772,2.1318035,1.5383345,1.5656652,1.5969005,1.6281357,1.6593709,1.6867018,2.5300527,3.3734035,4.2167544,5.056201,5.899552,6.910792,7.9259367,8.937177,9.948417,10.963562,10.151445,9.339331,8.52331,7.7111945,6.899079,8.175818,9.448653,10.725393,11.998228,13.274967,12.380859,11.490656,10.596548,9.706344,8.812236,9.093353,9.370565,9.651682,9.932799,10.213917,11.205634,12.201257,13.196879,14.192502,15.188125,13.1266,11.06898,9.007456,6.9459314,4.8883114,3.9083066,2.9322062,1.9561055,0.97610056,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,1.8741131,3.6740425,5.473972,7.2739015,9.073831,7.2582836,5.446641,3.631094,1.815547,0.0,0.31235218,0.62470436,0.93705654,1.2494087,1.5617609,3.7989833,6.036206,8.273428,10.510651,12.751778,10.967466,9.183154,7.4027467,5.618435,3.8380275,5.7511845,7.6682463,9.581403,11.498465,13.411622,14.286208,15.160794,16.039284,16.91387,17.788456,17.495626,17.202797,16.909966,16.617136,16.324306,16.20327,16.07833,15.957292,15.836256,15.711315,15.578565,15.441911,15.309161,15.172507,15.035853,14.930434,14.821111,14.7156925,14.606369,14.50095,13.083652,11.666354,10.249056,8.831758,7.4105554,7.6838636,7.9532676,8.2226715,8.492075,8.761478,7.336372,5.9073606,4.478349,3.0532427,1.6242313,1.7491722,1.8741131,1.999054,2.1239948,2.2489357,2.233318,2.2137961,2.1981785,2.1786566,2.1630387,3.4241607,4.689187,5.950309,7.211431,8.476458,6.918601,5.364649,3.8106966,2.2567444,0.698888,0.57394713,0.44510186,0.31625658,0.19131571,0.062470436,5.5130157,4.728231,3.9434462,3.1586614,2.3738766,1.5890918,1.4524376,1.3157835,1.183034,1.0463798,0.9136301,2.522244,4.1308575,5.743376,7.3519893,8.960603,7.703386,6.4422636,5.181142,3.9239242,2.6628022,2.377781,2.0927596,1.8077383,1.5227169,1.2376955,5.298274,9.362757,13.423335,17.487818,21.548395,25.815908,30.08342,34.35093,38.618443,42.885956,40.418373,37.95079,35.483208,33.015625,30.548042,25.70268,20.853413,16.008049,11.158782,6.3134184,6.785851,7.2582836,7.7307167,8.203149,8.675582,9.788337,10.904996,12.021654,13.134409,14.251068,13.021181,11.795199,10.569217,9.339331,8.113348,7.297328,6.481308,5.6691923,4.853172,4.037152,4.3065557,4.572055,4.841459,5.1069584,5.376362,5.2318993,5.0913405,4.9468775,4.806319,4.661856,5.1225758,5.5832953,6.044015,6.5008297,6.9615493,8.183627,9.405705,10.631687,11.8537655,13.075843,10.647305,8.218767,5.794133,3.3655949,0.93705654,1.2650263,1.5929961,1.9209659,2.2489357,2.5769055,3.06886,3.5647192,4.0605783,4.5564375,5.0483923,4.1503797,3.2484627,2.35045,1.4485333,0.5505207,1.2181735,1.8897307,2.5612879,3.2289407,3.900498,3.506153,3.1157131,2.7213683,2.330928,1.9365835,3.3851168,4.83365,6.278279,7.726812,9.175345,10.963562,12.755682,14.543899,16.33602,18.124235,16.757694,15.391153,14.020708,12.654168,11.287627,10.6590185,10.0265045,9.397896,8.769287,8.136774,7.363703,6.590631,5.8214636,5.0483923,4.2753205,3.5959544,2.9165885,2.233318,1.5539521,0.8745861,1.1322767,1.3899672,1.6476578,1.9053483,2.1630387,2.0615244,1.9561055,1.8545911,1.7530766,1.6515622,1.397776,1.1439898,0.8941081,0.64032197,0.38653582,0.79649806,1.2025559,1.6086137,2.018576,2.4246337,2.1708477,1.9131571,1.6593709,1.4055848,1.1517987,1.319688,1.4914817,1.6593709,1.8311646,1.999054,4.646239,7.289519,9.936704,12.579984,15.223265,13.411622,11.596075,9.780528,7.9649806,6.1494336,5.290465,4.4314966,3.5686235,2.7096553,1.8506867,1.7218413,1.5890918,1.4602464,1.3314011,1.1986516,0.96048295,0.71841,0.48024148,0.23816854,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.13274968,0.1756981,0.22255093,0.26940376,0.31235218,0.28892577,0.26159495,0.23816854,0.21083772,0.18741131,0.3513962,0.5114767,0.6754616,0.8355421,0.999527,0.80040246,0.60127795,0.39824903,0.19912452,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.20693332,0.39824903,0.58956474,0.78088045,0.97610056,0.80040246,0.62470436,0.44900626,0.27330816,0.10151446,0.13665408,0.1717937,0.20693332,0.23816854,0.27330816,0.22645533,0.1756981,0.12494087,0.07418364,0.023426414,0.14055848,0.26159495,0.37872702,0.4958591,0.61299115,0.97610056,1.3431144,1.7062237,2.0732377,2.436347,2.0459068,1.6593709,1.2689307,0.8784905,0.48805028,0.76135844,1.0307622,1.3040704,1.5773785,1.8506867,1.6164225,1.3860629,1.1517987,0.92143893,0.6871748,0.8667773,1.0463798,1.2259823,1.4055848,1.5890918,1.4602464,1.3314011,1.2064602,1.077615,0.94876975,1.0034313,1.0580931,1.116659,1.1713207,1.2259823,2.0029583,2.7799344,3.5569105,4.3338866,5.1108627,4.123049,3.1313305,2.1435168,1.1517987,0.1639849,0.30844778,0.45681506,0.60518235,0.75354964,0.9019169,1.0034313,1.1088502,1.2142692,1.319688,1.4251068,1.9561055,2.4831998,3.0141985,3.5451972,4.0761957,4.2870336,4.5017757,4.7126136,4.9234514,5.138193,4.806319,4.478349,4.1464753,3.8185053,3.4866312,2.8580225,2.2294137,1.5969005,0.96829176,0.3357786,0.7340276,1.1283722,1.5227169,1.9170616,2.3114061,4.21285,6.114294,8.011833,9.913278,11.810817,11.314958,10.819098,10.319335,9.823476,9.323712,8.203149,7.08649,5.9659266,4.845363,3.7247996,3.0532427,2.3855898,1.7140326,1.0463798,0.37482262,0.3357786,0.29673457,0.25378615,0.21474212,0.1756981,0.23035973,0.28502136,0.339683,0.39434463,0.44900626,1.5383345,2.631567,3.7208953,4.8102236,5.899552,4.970304,4.041056,3.1118085,2.1786566,1.2494087,3.59205,5.9346914,8.277332,10.619974,12.962616,11.275913,9.589212,7.898606,6.211904,4.5252023,7.016211,9.503315,11.994324,14.4853325,16.976341,18.38583,19.799223,21.212618,22.62601,24.039404,22.450314,20.861221,19.276033,17.686943,16.101755,14.903104,13.708356,12.513609,11.318862,10.124115,12.326198,14.528281,16.734268,18.936352,21.138433,18.858263,16.581997,14.30573,12.025558,9.749292,9.807858,9.866425,9.921086,9.979652,10.0382185,10.116306,10.198298,10.276386,10.358379,10.436467,10.510651,10.58093,10.655114,10.729298,10.799577,10.81129,10.819098,10.8308115,10.838621,10.850334,9.647778,8.445222,7.2426662,6.04011,4.8375545,4.575959,4.318269,4.056674,3.7989833,3.5373883,3.2016098,2.8658314,2.533957,2.1981785,1.8623998,1.9404879,2.018576,2.096664,2.1708477,2.2489357,2.951728,3.6545205,4.357313,5.0601053,5.7628975,6.7624245,7.7619514,8.761478,9.761005,10.764437,9.636065,8.511597,7.387129,6.262661,5.138193,6.5984397,8.062591,9.526741,10.986988,12.4511385,11.924045,11.39695,10.865952,10.338858,9.811763,9.639969,9.468176,9.296382,9.120684,8.94889,10.471607,11.994324,13.51704,15.039758,16.562475,13.759113,10.951848,8.148487,5.3412223,2.5378613,2.0302892,1.5227169,1.0151446,0.5075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,1.0619974,2.0888553,3.1118085,4.138666,5.1616197,4.1308575,3.096191,2.0654287,1.0307622,0.0,0.24988174,0.4997635,0.74964523,0.999527,1.2494087,3.4983444,5.7511845,8.00012,10.249056,12.501896,10.514555,8.531119,6.5437784,4.560342,2.5769055,5.2084727,7.8400397,10.471607,13.103174,15.738646,16.574188,17.413633,18.249176,19.088623,19.924164,19.799223,19.670378,19.541533,19.416592,19.287746,18.81922,18.35069,17.886066,17.417538,16.94901,16.995863,17.03881,17.085665,17.128613,17.175465,17.066143,16.95682,16.843592,16.734268,16.624945,15.008522,13.396004,11.779582,10.167064,8.550641,8.710721,8.870802,9.030883,9.190963,9.351044,7.7658563,6.184573,4.60329,3.0220075,1.43682,1.6008049,1.7608855,1.9248703,2.0888553,2.2489357,2.2216048,2.194274,2.1669433,2.1396124,2.1122816,3.5373883,4.9624953,6.387602,7.812709,9.237816,7.570636,5.9073606,4.2440853,2.5769055,0.9136301,0.7418364,0.57394713,0.40215343,0.23426414,0.062470436,3.6857557,3.1508527,2.612045,2.0732377,1.5383345,0.999527,0.80040246,0.60127795,0.39824903,0.19912452,0.0,2.2372224,4.474445,6.7116675,8.94889,11.186112,9.187058,7.1880045,5.1889505,3.1859922,1.1869383,1.2142692,1.2376955,1.261122,1.2884527,1.3118792,5.9737353,10.6355915,15.3013525,19.96321,24.625065,26.163399,27.701735,29.236164,30.774498,32.31283,29.025326,25.73782,22.450314,19.162806,15.875299,13.825488,11.775677,9.725866,7.676055,5.6262436,6.649197,7.676055,8.699008,9.725866,10.748819,12.138786,13.524849,14.9109125,16.300879,17.686943,15.961197,14.239355,12.513609,10.787864,9.062118,7.800996,6.5359693,5.2748475,4.0137253,2.7486992,3.1625657,3.5764325,3.9863946,4.4002614,4.814128,4.3260775,3.8380275,3.349977,2.8619268,2.3738766,2.912684,3.4514916,3.9863946,4.5252023,5.0640097,7.012306,8.960603,10.912805,12.861101,14.813302,12.013845,9.21439,6.4110284,3.611572,0.81211567,1.0112402,1.2142692,1.4133936,1.6125181,1.8116426,2.7135596,3.611572,4.513489,5.4115014,6.3134184,5.1889505,4.0644827,2.9361105,1.8116426,0.6871748,1.5266213,2.3621633,3.2016098,4.037152,4.8765984,4.298747,3.7247996,3.1508527,2.5769055,1.999054,3.775557,5.548156,7.3246584,9.101162,10.87376,13.173453,15.473146,17.776743,20.076437,22.37613,20.61134,18.850454,17.085665,15.324779,13.563893,12.099743,10.639496,9.175345,7.7111945,6.250948,5.563773,4.8765984,4.1894236,3.4983444,2.8111696,2.2996929,1.7882162,1.2767396,0.76135844,0.24988174,0.23816854,0.22645533,0.21083772,0.19912452,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.31235218,0.5622339,0.81211567,1.0619974,1.3118792,1.0737107,0.8394465,0.60127795,0.3631094,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,2.639376,5.1499066,7.6643414,10.174872,12.689307,11.560935,10.436467,9.311999,8.187531,7.0630636,6.114294,5.1616197,4.21285,3.2640803,2.3114061,2.1513257,1.9873407,1.8233559,1.6632754,1.4992905,1.1986516,0.9019169,0.60127795,0.30063897,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.6637484,1.1986516,1.737459,2.2762666,2.8111696,2.260649,1.7140326,1.1635119,0.61299115,0.062470436,0.30063897,0.5388075,0.77307165,1.0112402,1.2494087,1.1127546,0.97610056,0.8394465,0.698888,0.5622339,0.4997635,0.43729305,0.37482262,0.31235218,0.24988174,0.22645533,0.19912452,0.1756981,0.14836729,0.12494087,0.22645533,0.3240654,0.42557985,0.5231899,0.62470436,1.7608855,2.900971,4.037152,5.173333,6.3134184,5.087436,3.8614538,2.639376,1.4133936,0.18741131,0.3631094,0.5388075,0.7106012,0.8862993,1.0619974,1.175225,1.2884527,1.4016805,1.5110037,1.6242313,2.0888553,2.5495746,3.0141985,3.474918,3.9356375,4.3260775,4.7126136,5.099149,5.4856853,5.8761253,5.5013027,5.12648,4.7516575,4.376835,3.998108,3.2484627,2.4988174,1.7491722,0.999527,0.24988174,0.737932,1.2259823,1.7140326,2.1981785,2.6862288,3.6232853,4.564246,5.5013027,6.4383593,7.375416,7.0357327,6.699954,6.364176,6.0244927,5.688714,4.911738,4.138666,3.3616903,2.5886188,1.8116426,1.4485333,1.0893283,0.7262188,0.3631094,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,1.5734742,3.0259118,4.474445,5.9268827,7.375416,6.1884775,5.001539,3.8106966,2.6237583,1.43682,4.2753205,7.113821,9.948417,12.786918,15.625418,12.798631,9.975748,7.1489606,4.3260775,1.4992905,5.263134,9.023073,12.786918,16.55076,20.310701,22.149673,23.988647,25.823717,27.66269,29.501663,27.623646,25.749533,23.87542,22.001307,20.12329,18.600573,17.073952,15.551234,14.024612,12.501896,15.063184,17.624472,20.18576,22.750952,25.31224,22.575254,19.838268,17.101282,14.364296,11.623405,11.639023,11.650736,11.66245,11.674163,11.685876,11.435994,11.186112,10.936231,10.686349,10.436467,10.748819,11.061172,11.373524,11.685876,11.998228,11.736633,11.475039,11.213444,10.951848,10.686349,9.526741,8.36323,7.1997175,6.036206,4.8765984,4.4119744,3.951255,3.4866312,3.0259118,2.5612879,2.4871042,2.4129205,2.338737,2.260649,2.1864653,2.3114061,2.436347,2.5612879,2.6862288,2.8111696,3.3734035,3.9356375,4.5017757,5.0640097,5.6262436,6.6140575,7.601871,8.58578,9.573594,10.561408,9.124588,7.687768,6.250948,4.814128,3.3734035,5.024966,6.676528,8.324185,9.975748,11.623405,11.4633255,11.29934,11.139259,10.975275,10.81129,10.186585,9.561881,8.937177,8.312472,7.687768,9.737579,11.787391,13.837202,15.8870125,17.936825,14.387722,10.838621,7.2856145,3.736513,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24988174,0.4997635,0.74964523,0.999527,1.2494087,0.999527,0.74964523,0.4997635,0.24988174,0.0,0.18741131,0.37482262,0.5622339,0.74964523,0.93705654,3.2016098,5.462259,7.726812,9.987461,12.24811,10.061645,7.8751793,5.688714,3.4983444,1.3118792,4.661856,8.011833,11.361811,14.711788,18.061766,18.862167,19.662569,20.462973,21.263374,22.063778,22.098917,22.13796,22.1731,22.212145,22.251188,21.439074,20.623053,19.810938,18.998821,18.186707,18.41316,18.635712,18.862167,19.088623,19.311174,19.20185,19.088623,18.975395,18.862167,18.74894,16.937298,15.125654,13.314012,11.498465,9.686822,9.737579,9.788337,9.839094,9.885946,9.936704,8.1992445,6.461786,4.7243266,2.9868677,1.2494087,1.4485333,1.6515622,1.8506867,2.0498111,2.2489357,2.2137961,2.174752,2.135708,2.1005683,2.0615244,3.6506162,5.2358036,6.824895,8.413987,9.999174,8.226576,6.4500723,4.6735697,2.900971,1.1244678,0.9136301,0.698888,0.48805028,0.27330816,0.062470436,3.1508527,2.815074,2.4792955,2.1435168,1.8116426,1.475864,1.9209659,2.366068,2.8111696,3.2562714,3.7013733,4.9546866,6.211904,7.465217,8.718531,9.975748,8.246098,6.5164475,4.786797,3.0532427,1.3235924,1.9092526,2.4910088,3.0727646,3.6545205,4.2362766,7.5159745,10.795672,14.079274,17.358973,20.63867,23.004738,25.370806,27.740778,30.106846,32.476818,28.615364,24.75391,20.89636,17.034906,13.173453,12.064603,10.955752,9.846903,8.734148,7.6252975,10.006983,12.388668,14.774258,17.155943,19.537628,19.330696,19.123762,18.916828,18.705992,18.499058,16.324306,14.145649,11.966993,9.788337,7.6135845,6.5633,5.5169206,4.4705405,3.4241607,2.3738766,2.67842,2.9868677,3.2914112,3.5959544,3.900498,3.7599394,3.619381,3.4788225,3.338264,3.2016098,3.4280653,3.6545205,3.8809757,4.1113358,4.337791,6.3134184,8.289046,10.260769,12.236397,14.212025,11.639023,9.066022,6.493021,3.9239242,1.3509232,1.53443,1.7218413,1.9053483,2.0888553,2.2762666,2.87364,3.474918,4.0761957,4.6735697,5.2748475,4.388548,3.4983444,2.612045,1.7257458,0.8394465,1.8663043,2.8970666,3.9278288,4.958591,5.989353,5.423215,4.8570766,4.290938,3.7287042,3.1625657,4.7516575,6.3407493,7.9337454,9.522837,11.111929,12.771299,14.426766,16.086138,17.741604,19.400974,18.038338,16.679607,15.320874,13.958238,12.599506,12.076316,11.549222,11.0260315,10.498938,9.975748,8.995743,8.019642,7.043542,6.0635366,5.087436,4.2167544,3.3421683,2.4714866,1.5969005,0.7262188,0.679366,0.62860876,0.58175594,0.5349031,0.48805028,0.6520352,0.8160201,0.98390937,1.1478943,1.3118792,1.0580931,0.80821127,0.5544251,0.30063897,0.05075723,0.6559396,1.261122,1.8663043,2.4714866,3.076669,2.4792955,1.8858263,1.2884527,0.6949836,0.10151446,0.19131571,0.28502136,0.37872702,0.46852827,0.5622339,2.5964274,4.630621,6.6687193,8.702912,10.737106,10.295909,9.858616,9.4174185,8.976221,8.538928,7.363703,6.1884775,5.0132523,3.8380275,2.6628022,2.4480603,2.2372224,2.0263848,1.8116426,1.6008049,1.2884527,0.98000497,0.6715572,0.359205,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.09761006,0.19522011,0.29283017,0.39044023,0.48805028,0.39434463,0.30063897,0.21083772,0.11713207,0.023426414,0.031235218,0.03513962,0.039044023,0.046852827,0.05075723,0.12103647,0.19522011,0.26940376,0.339683,0.41386664,0.3357786,0.25769055,0.1796025,0.10151446,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10541886,0.15617609,0.21083772,0.26159495,0.26549935,0.26940376,0.26940376,0.27330816,0.27330816,0.21864653,0.1639849,0.10932326,0.05466163,0.0,0.0,0.0,0.0,0.0,0.0,0.13665408,0.26940376,0.40605783,0.5388075,0.6754616,0.9956226,1.319688,1.6437533,1.9639144,2.2879796,1.8389735,1.3938715,0.94486535,0.4958591,0.05075723,0.26940376,0.48414588,0.7027924,0.92143893,1.1361811,1.0541886,0.96829176,0.8823949,0.79649806,0.7106012,0.6442264,0.57785153,0.5114767,0.44119745,0.37482262,0.3631094,0.3513962,0.3357786,0.3240654,0.31235218,0.41386664,0.5192855,0.62079996,0.7223144,0.8238289,1.6827974,2.541766,3.39683,4.2557983,5.1108627,4.126953,3.1430438,2.1591344,1.1713207,0.18741131,0.32016098,0.45291066,0.58566034,0.71841,0.8511597,0.94876975,1.0502841,1.1517987,1.2494087,1.3509232,1.7686942,2.1864653,2.6042364,3.018103,3.435874,3.9083066,4.380739,4.853172,5.3256044,5.801942,5.380266,4.958591,4.5408196,4.1191444,3.7013733,3.0298162,2.358259,1.6906061,1.0190489,0.3513962,0.76916724,1.1908426,1.6086137,2.0302892,2.4480603,3.174279,3.900498,4.6267166,5.349031,6.0752497,6.001066,5.930787,5.8566036,5.786324,5.7121406,5.9464045,6.1767645,6.4110284,6.6413884,6.8756523,5.704332,4.5369153,3.3655949,2.194274,1.0268579,1.6086137,2.1903696,2.7721257,3.3538816,3.9395418,3.2367494,2.533957,1.8311646,1.1283722,0.42557985,2.6042364,4.786797,6.9654536,9.14411,11.326671,9.288573,7.2543793,5.2201858,3.1859922,1.1517987,3.506153,5.860508,8.214863,10.569217,12.923572,13.09927,13.271063,13.442857,13.614651,13.786445,14.376009,14.969479,15.559043,16.148607,16.738173,18.74894,20.76361,22.774378,24.78905,26.799816,24.906181,23.01645,21.122816,19.229181,17.335546,16.457056,15.578565,14.69617,13.817679,12.939189,14.446288,15.957292,17.468296,18.9793,20.486399,19.553246,18.61619,17.683039,16.745981,15.812829,14.735214,13.657599,12.579984,11.502369,10.424754,10.600452,10.77615,10.951848,11.123642,11.29934,11.603884,11.904523,12.209065,12.509705,12.814248,12.330102,11.845957,11.365715,10.881569,10.401327,9.456462,8.511597,7.5667315,6.621866,5.6730967,5.368553,5.0601053,4.7516575,4.4432096,4.138666,3.9863946,3.8380275,3.6857557,3.5373883,3.3890212,3.5100577,3.631094,3.7560349,3.8770714,3.998108,4.3065557,4.6150036,4.9234514,5.2318993,5.5364423,6.46569,7.3910336,8.320281,9.245625,10.174872,9.187058,8.1992445,7.211431,6.223617,5.2358036,6.688241,8.140678,9.597021,11.0494585,12.501896,12.076316,11.654641,11.232965,10.81129,10.38571,10.268578,10.151445,10.034314,9.917182,9.80005,11.23687,12.6697855,14.106606,15.539521,16.976341,13.610746,10.2451515,6.8795567,3.513962,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19912452,0.39824903,0.60127795,0.80040246,0.999527,0.80040246,0.60127795,0.39824903,0.19912452,0.0,0.14836729,0.30063897,0.44900626,0.60127795,0.74964523,2.5612879,4.376835,6.1884775,8.00012,9.811763,8.706817,7.5979667,6.4891167,5.3841705,4.2753205,6.3329406,8.39056,10.44818,12.5058,14.56342,15.570756,16.578093,17.585428,18.592764,19.6001,19.443924,19.283842,19.127666,18.97149,18.81141,19.596195,20.38098,21.165764,21.954454,22.739239,21.989594,21.243853,20.494207,19.748466,18.998821,18.48344,17.96806,17.456583,16.941202,16.42582,15.473146,14.524376,13.575606,12.626837,11.674163,11.326671,10.979179,10.631687,10.284196,9.936704,8.324185,6.7116675,5.099149,3.4866312,1.8741131,1.9561055,2.0341935,2.1161861,2.194274,2.2762666,2.2957885,2.3153105,2.3348327,2.3543546,2.3738766,3.7989833,5.2201858,6.6413884,8.066495,9.487698,7.8361354,6.1884775,4.5369153,2.8892577,1.2376955,0.999527,0.76135844,0.5231899,0.28892577,0.05075723,2.612045,2.4792955,2.3465457,2.2137961,2.0810463,1.9482968,3.0415294,4.1308575,5.2201858,6.309514,7.3988423,7.6721506,7.9454584,8.218767,8.488171,8.761478,7.3012323,5.840986,4.380739,2.9243972,1.4641509,2.6042364,3.7443218,4.884407,6.0205884,7.1606736,9.058213,10.955752,12.853292,14.750832,16.64837,19.846077,23.043781,26.241488,29.439194,32.636898,28.205402,23.773905,19.338505,14.907008,10.475512,10.303718,10.135828,9.964035,9.796145,9.6243515,13.364769,17.105186,20.845604,24.586021,28.326439,26.522604,24.718771,22.91884,21.115007,19.311174,16.683512,14.051944,11.424281,8.792714,6.1611466,5.3295093,4.4978714,3.6662338,2.8306916,1.999054,2.1981785,2.3933985,2.592523,2.7916477,2.9868677,3.193801,3.4007344,3.611572,3.8185053,4.025439,3.9434462,3.8614538,3.775557,3.6935644,3.611572,5.610626,7.6135845,9.612638,11.611692,13.610746,11.268105,8.921559,6.578918,4.2323723,1.8858263,2.05762,2.2294137,2.397303,2.5690966,2.736986,3.0376248,3.338264,3.638903,3.9356375,4.2362766,3.5881457,2.9361105,2.2879796,1.6359446,0.9878138,2.2098918,3.4319696,4.6540475,5.8761253,7.098203,6.5437784,5.989353,5.434928,4.8805027,4.3260775,5.7316628,7.1333427,8.538928,9.944512,11.350098,12.365242,13.380386,14.395531,15.410676,16.42582,15.469242,14.508759,13.55218,12.595602,11.639023,12.0489855,12.4628525,12.8767185,13.286681,13.700547,12.431617,11.166591,9.897659,8.628729,7.363703,6.1299114,4.8961205,3.6662338,2.4324427,1.1986516,1.116659,1.0346665,0.95267415,0.8706817,0.78868926,1.116659,1.4485333,1.7765031,2.1083772,2.436347,1.9561055,1.475864,0.9956226,0.5192855,0.039044023,0.9956226,1.9561055,2.9165885,3.8770714,4.8375545,3.8848803,2.9322062,1.979532,1.0268579,0.07418364,0.26159495,0.44510186,0.62860876,0.8160201,0.999527,2.5573835,4.11524,5.6730967,7.230953,8.78881,9.030883,9.276859,9.522837,9.768814,10.010887,8.6131115,7.211431,5.813655,4.4119744,3.0141985,2.7486992,2.4871042,2.2255092,1.9639144,1.698415,1.3782539,1.0580931,0.7418364,0.42167544,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.15617609,0.31625658,0.47243267,0.62860876,0.78868926,0.64032197,0.49195468,0.3435874,0.19912452,0.05075723,0.046852827,0.046852827,0.042948425,0.039044023,0.039044023,0.19522011,0.3513962,0.5114767,0.6676528,0.8238289,0.6715572,0.5153811,0.359205,0.20693332,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10541886,0.21083772,0.31625658,0.42167544,0.5231899,0.5036679,0.48414588,0.46462387,0.44510186,0.42557985,0.339683,0.25378615,0.1717937,0.08589685,0.0,0.0,0.0,0.0,0.0,0.0,0.24597734,0.48805028,0.7340276,0.98000497,1.2259823,1.3314011,1.4407244,1.5461433,1.6554666,1.7608855,1.4172981,1.0737107,0.7262188,0.38263142,0.039044023,0.23426414,0.43338865,0.62860876,0.8277333,1.0268579,0.9917182,0.96048295,0.92924774,0.8941081,0.8628729,0.78868926,0.71841,0.6442264,0.57394713,0.4997635,0.4997635,0.4997635,0.4997635,0.4997635,0.4997635,0.60518235,0.7106012,0.8160201,0.92143893,1.0268579,1.6008049,2.1786566,2.7565079,3.3343596,3.912211,3.1664703,2.4207294,1.678893,0.93315214,0.18741131,0.27721256,0.3670138,0.45681506,0.5466163,0.63641757,0.7262188,0.81211567,0.9019169,0.9878138,1.0737107,1.4485333,1.8194515,2.194274,2.5651922,2.9361105,3.49444,4.0527697,4.6110992,5.169429,5.7238536,5.2592297,4.794606,4.3299823,3.8653584,3.4007344,2.8111696,2.2216048,1.6281357,1.038571,0.44900626,0.80430686,1.1557031,1.5070993,1.8584955,2.2137961,2.7252727,3.2367494,3.7482262,4.263607,4.775084,4.9663997,5.1616197,5.3529353,5.5442514,5.735567,6.9771667,8.218767,9.456462,10.698062,11.935758,9.96013,7.984503,6.0049706,4.029343,2.0498111,3.213323,4.380739,5.5442514,6.7116675,7.8751793,6.446168,5.0132523,3.5842414,2.15523,0.7262188,3.6349986,6.5437784,9.456462,12.365242,15.274021,12.392572,9.511124,6.6257706,3.7443218,0.8628729,2.736986,4.607195,6.481308,8.351517,10.22563,13.396004,16.56638,19.736753,22.903223,26.073599,23.492788,20.911978,18.327265,15.746454,13.16174,15.348206,17.538574,5052.0,21.911505,24.101875,22.188719,20.279465,18.370213,16.46096,14.551707,14.313539,14.079274,13.845011,13.610746,13.376482,13.833297,14.2901125,14.746927,15.203742,15.660558,16.531239,17.398016,18.264793,19.13157,19.998348,17.831406,15.664462,13.497519,11.330575,9.163632,9.761005,10.362284,10.963562,11.560935,12.162213,12.455043,12.747873,13.040704,13.333533,13.626364,12.923572,12.220779,11.517986,10.815194,10.112402,9.386183,8.65606,7.929841,7.2036223,6.473499,6.321227,6.168956,6.016684,5.8644123,5.7121406,5.4856853,5.263134,5.036679,4.814128,4.5876727,4.7087092,4.825841,4.9468775,5.067914,5.1889505,5.239708,5.2943697,5.3451266,5.395884,5.4505453,6.3173227,7.1841,8.050878,8.921559,9.788337,9.249529,8.710721,8.175818,7.6370106,7.098203,8.355421,9.608734,10.865952,12.119265,13.376482,12.693212,12.009941,11.326671,10.6434,9.964035,10.354475,10.741011,11.131451,11.521891,11.912332,12.732256,13.55218,14.372105,15.192029,16.011953,12.83377,9.651682,6.473499,3.2914112,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14836729,0.30063897,0.44900626,0.60127795,0.74964523,0.60127795,0.44900626,0.30063897,0.14836729,0.0,0.113227665,0.22645533,0.3357786,0.44900626,0.5622339,1.9248703,3.2875066,4.650143,6.012779,7.375416,7.348085,7.320754,7.2934237,7.266093,7.238762,8.0040245,8.769287,9.530646,10.295909,11.061172,12.2793455,13.493614,14.707883,15.9221525,17.136421,16.785025,16.43363,16.07833,15.726933,15.375536,17.757221,20.138906,22.524496,24.906181,27.287867,25.566027,23.84809,22.126247,20.40831,18.68647,17.768934,16.8514,15.933866,15.016331,14.098797,14.012899,13.923099,13.837202,13.751305,13.661504,12.915763,12.173926,11.428185,10.682445,9.936704,8.449126,6.9615493,5.473972,3.9863946,2.4988174,2.4597735,2.4207294,2.3816853,2.338737,2.2996929,2.377781,2.455869,2.533957,2.6081407,2.6862288,3.9434462,5.2045684,6.461786,7.719003,8.976221,7.4495993,5.9229784,4.4002614,2.87364,1.3509232,1.0893283,0.8238289,0.5622339,0.30063897,0.039044023,2.0732377,2.1435168,2.2137961,2.2840753,2.3543546,2.4246337,4.1581883,5.8956475,7.629202,9.366661,11.100216,10.389614,9.679013,8.968412,8.261715,7.551114,6.3602715,5.169429,3.978586,2.7916477,1.6008049,3.2992198,4.9937305,6.6921453,8.39056,10.088976,10.604357,11.115833,11.631214,12.146595,12.661977,16.69132,20.716759,24.746101,28.77154,32.800884,27.795439,22.789995,17.784552,12.779109,7.773665,8.546737,9.315904,10.085071,10.8542385,11.623405,16.722555,21.821705,26.916948,32.016098,37.111343,33.71451,30.317684,26.920853,23.524023,20.12329,17.042715,13.958238,10.877665,7.793187,4.7126136,4.095718,3.4788225,2.8619268,2.241127,1.6242313,1.7140326,1.8038338,1.893635,1.9834363,2.0732377,2.631567,3.1859922,3.7404175,4.2948427,4.8492675,4.4588275,4.0644827,3.6740425,3.279698,2.8892577,4.911738,6.9381227,8.964508,10.986988,13.013372,10.893282,8.777096,6.66091,4.5408196,2.4246337,2.5808098,2.7330816,2.8892577,3.0454338,3.2016098,3.2016098,3.2016098,3.2016098,3.2016098,3.2016098,2.787743,2.3738766,1.9639144,1.5500476,1.1361811,2.5534792,3.9668727,5.3841705,6.7975645,8.210958,7.6682463,7.1216297,6.578918,6.0323014,5.4856853,6.707763,7.9259367,9.148014,10.366188,11.588266,11.959184,12.334006,12.704925,13.075843,13.450665,12.89624,12.341816,11.783486,11.229061,10.674636,12.025558,13.376482,14.723501,16.074425,17.425346,15.867491,14.309634,12.751778,11.193921,9.636065,8.043069,6.453977,4.860981,3.2679846,1.6749885,1.5578566,1.4407244,1.3235924,1.2064602,1.0893283,1.5812829,2.077142,2.5730011,3.06886,3.5608149,2.854118,2.1474214,1.4407244,0.7340276,0.023426414,1.33921,2.6549935,3.970777,5.2865605,6.5984397,5.290465,3.978586,2.6706111,1.358732,0.05075723,0.3279698,0.60518235,0.8823949,1.1596074,1.43682,2.5183394,3.5959544,4.677474,5.758993,6.8366084,7.7658563,8.699008,9.628256,10.557504,11.486752,9.86252,8.238289,6.6140575,4.985922,3.3616903,3.049338,2.736986,2.4246337,2.1122816,1.7999294,1.4680552,1.1400855,0.80821127,0.48024148,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.21864653,0.43338865,0.6520352,0.8706817,1.0893283,0.8862993,0.6832704,0.48024148,0.27721256,0.07418364,0.06637484,0.05466163,0.046852827,0.03513962,0.023426414,0.26940376,0.5114767,0.75354964,0.9956226,1.2376955,1.0034313,0.77307165,0.5388075,0.30844778,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15617609,0.31625658,0.47243267,0.62860876,0.78868926,0.74574083,0.7027924,0.659844,0.61689556,0.57394713,0.46071947,0.3435874,0.23035973,0.113227665,0.0,0.0,0.0,0.0,0.0,0.0,0.3553006,0.7106012,1.0659018,1.4212024,1.7765031,1.6671798,1.5617609,1.4524376,1.3431144,1.2376955,0.9956226,0.75354964,0.5114767,0.26940376,0.023426414,0.20302892,0.37872702,0.5583295,0.7340276,0.9136301,0.93315214,0.95267415,0.97219616,0.9917182,1.0112402,0.93315214,0.8589685,0.78088045,0.7027924,0.62470436,0.63641757,0.6481308,0.6637484,0.6754616,0.6871748,0.79649806,0.9019169,1.0112402,1.116659,1.2259823,1.5227169,1.8194515,2.1161861,2.416825,2.7135596,2.2059872,1.7023194,1.1986516,0.6910792,0.18741131,0.23426414,0.28111696,0.3318742,0.37872702,0.42557985,0.4997635,0.57394713,0.6481308,0.7262188,0.80040246,1.1283722,1.456342,1.7843118,2.1083772,2.436347,3.0805733,3.7208953,4.365122,5.009348,5.64967,5.138193,4.630621,4.1191444,3.611572,3.1000953,2.5886188,2.0810463,1.5695697,1.0580931,0.5505207,0.8355421,1.1205635,1.4055848,1.6906061,1.9756275,2.2762666,2.5769055,2.87364,3.174279,3.474918,3.9317331,4.388548,4.8492675,5.3060827,5.7628975,8.011833,10.256865,12.5058,14.750832,16.999767,14.215929,11.428185,8.644346,5.860508,3.076669,4.8219366,6.571109,8.316377,10.065549,11.810817,9.655587,7.4964523,5.3412223,3.182088,1.0268579,4.6657605,8.304664,11.943566,15.586374,19.225277,15.4965725,11.763964,8.03526,4.3065557,0.57394713,1.9639144,3.3538816,4.743849,6.133816,7.523783,13.692739,19.861694,26.026745,32.1957,38.360752,32.605663,26.854479,21.095486,15.344301,9.589212,11.951375,14.313539,16.675701,19.037865,21.400028,19.471254,17.546383,15.617609,13.688834,11.763964,12.173926,12.583888,12.993851,13.403813,13.813775,13.216402,12.622932,12.025558,11.43209,10.838621,13.509232,16.175938,18.84655,21.51716,24.187773,20.931501,17.671324,14.415053,11.158782,7.898606,8.925464,9.948417,10.975275,11.998228,13.025085,13.306203,13.591225,13.872341,14.153459,14.438479,13.513136,12.591698,11.6702585,10.748819,9.823476,9.315904,8.804427,8.296855,7.785378,7.2739015,7.277806,7.28171,7.28171,7.2856145,7.2856145,6.98888,6.688241,6.387602,6.086963,5.786324,5.903456,6.0205884,6.141625,6.2587566,6.375889,6.17286,5.969831,5.7668023,5.563773,5.3607445,6.168956,6.9771667,7.785378,8.59359,9.4018,9.311999,9.226103,9.136301,9.050405,8.960603,10.018696,11.076789,12.134882,13.192975,14.251068,13.306203,12.365242,11.424281,10.479416,9.538455,10.436467,11.330575,12.228588,13.1266,14.024612,14.231546,14.434575,14.641508,14.844538,15.051471,12.05289,9.058213,6.0635366,3.06886,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,1.2884527,2.1981785,3.1118085,4.025439,4.939069,5.989353,7.043542,8.093826,9.148014,10.198298,9.671205,9.14411,8.617016,8.089922,7.562827,8.98403,10.409137,11.8303385,13.251541,14.676648,14.126127,13.579511,13.032895,12.486279,11.935758,15.918248,19.896833,23.879324,27.85791,31.836496,29.146362,26.452326,23.758287,21.068155,18.374117,17.054428,15.734741,14.415053,13.095366,11.775677,12.548749,13.325725,14.098797,14.875772,15.648844,14.508759,13.364769,12.220779,11.080693,9.936704,8.574067,7.211431,5.8487945,4.4861584,3.1235218,2.9634414,2.803361,2.6432803,2.4831998,2.3231194,2.4597735,2.5964274,2.7291772,2.8658314,2.998581,4.0918136,5.185046,6.278279,7.3715115,8.460839,7.0630636,5.661383,4.263607,2.8619268,1.4641509,1.175225,0.8862993,0.60127795,0.31235218,0.023426414,1.5383345,1.8116426,2.0810463,2.3543546,2.6276627,2.900971,5.278752,7.660437,10.0382185,12.419904,14.801589,13.107079,11.416472,9.721962,8.031356,6.336845,5.4193106,4.4978714,3.5764325,2.6588979,1.737459,3.9942036,6.2470436,8.503788,10.756628,13.013372,12.146595,11.275913,10.409137,9.542359,8.675582,13.532659,18.389734,23.24681,28.103888,32.960964,27.385477,21.806087,16.2306,10.651209,5.0757227,6.785851,8.495979,10.206107,11.916236,13.626364,20.080341,26.534317,32.9922,39.446175,45.900154,40.90642,35.916595,30.922867,25.929136,20.93931,17.40192,13.868437,10.331048,6.7975645,3.2640803,2.8619268,2.455869,2.0537157,1.6515622,1.2494087,1.2337911,1.2142692,1.1986516,1.1791295,1.1635119,2.0654287,2.9673457,3.8692627,4.7711797,5.6730967,4.9742084,4.271416,3.5686235,2.8658314,2.1630387,4.21285,6.262661,8.312472,10.362284,12.412095,10.522364,8.632633,6.7429028,4.853172,2.9634414,3.1039999,3.240654,3.3812122,3.521771,3.6623292,3.3616903,3.0610514,2.7643168,2.463678,2.1630387,1.9873407,1.8116426,1.6359446,1.4641509,1.2884527,2.893162,4.5017757,6.1103897,7.719003,9.323712,8.78881,8.253906,7.719003,7.1841,6.649197,7.6838636,8.718531,9.753197,10.791768,11.826434,11.553126,11.283723,11.014318,10.744915,10.475512,10.323239,10.170968,10.018696,9.866425,9.714153,11.998228,14.286208,16.574188,18.862167,21.150146,19.303364,17.456583,15.605896,13.759113,11.912332,9.96013,8.007929,6.055728,4.1035266,2.1513257,1.999054,1.8467822,1.6906061,1.5383345,1.3860629,2.0459068,2.7057507,3.3655949,4.029343,4.689187,3.7521305,2.8189783,1.8819219,0.94876975,0.011713207,1.6827974,3.3538816,5.0210614,6.6921453,8.36323,6.6960497,5.02887,3.3616903,1.6906061,0.023426414,0.39434463,0.76526284,1.1361811,1.5031948,1.8741131,2.4792955,3.0805733,3.6818514,4.283129,4.8883114,6.5008297,8.117252,9.733675,11.346193,12.962616,11.111929,9.261242,7.4105554,5.563773,3.7130866,3.349977,2.9868677,2.6237583,2.260649,1.901444,1.5617609,1.2181735,0.8784905,0.5388075,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.27721256,0.5544251,0.8316377,1.1088502,1.3860629,1.1283722,0.8706817,0.61689556,0.359205,0.10151446,0.08199245,0.06637484,0.046852827,0.031235218,0.011713207,0.339683,0.6676528,0.9956226,1.3235924,1.6515622,1.33921,1.0307622,0.71841,0.40996224,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21083772,0.42167544,0.62860876,0.8394465,1.0502841,0.98390937,0.92143893,0.8550641,0.78868926,0.7262188,0.58175594,0.43338865,0.28892577,0.14446288,0.0,0.0,0.0,0.0,0.0,0.0,0.46462387,0.92924774,1.3938715,1.8584955,2.3231194,2.0029583,1.678893,1.358732,1.0346665,0.7106012,0.57394713,0.43338865,0.29283017,0.15227169,0.011713207,0.1717937,0.3279698,0.48414588,0.6442264,0.80040246,0.8706817,0.94486535,1.0190489,1.0893283,1.1635119,1.0815194,0.9956226,0.9136301,0.8316377,0.74964523,0.77307165,0.80040246,0.8238289,0.8511597,0.8745861,0.98390937,1.0932326,1.2064602,1.3157835,1.4251068,1.4407244,1.4602464,1.475864,1.4953861,1.5110037,1.2494087,0.98390937,0.71841,0.45291066,0.18741131,0.19131571,0.19912452,0.20302892,0.20693332,0.21083772,0.27330816,0.3357786,0.39824903,0.46071947,0.5231899,0.80821127,1.0893283,1.3743496,1.6554666,1.9365835,2.6667068,3.3929255,4.1191444,4.8492675,5.575486,5.0210614,4.466636,3.9083066,3.3538816,2.7994564,2.3699722,1.9404879,1.5110037,1.0815194,0.6481308,0.8667773,1.0854238,1.3040704,1.5188124,1.737459,1.8233559,1.9131571,1.999054,2.0888553,2.174752,2.8970666,3.619381,4.3416953,5.0640097,5.786324,9.042596,12.298867,15.551234,18.807507,22.063778,18.471727,14.875772,11.283723,7.6916723,4.0996222,6.4305506,8.761478,11.088503,13.419431,15.750359,12.8650055,9.979652,7.094299,4.2089458,1.3235924,5.6965227,10.065549,14.434575,18.8036,23.176533,18.596668,14.020708,9.440845,4.8648853,0.28892577,1.1947471,2.1005683,3.0102942,3.9161155,4.825841,13.989473,23.153105,32.32064,41.484276,50.65181,41.722443,32.796978,23.86761,14.938243,6.012779,8.550641,11.088503,13.626364,16.164225,18.698183,16.75379,14.809398,12.8650055,10.920613,8.976221,10.03041,11.084598,12.138786,13.196879,14.251068,12.603411,10.955752,9.308095,7.660437,6.012779,10.48332,14.957765,19.428307,23.90275,28.373291,24.02769,19.682093,15.332587,10.983084,6.6374836,8.086017,9.538455,10.986988,12.439425,13.887959,14.161267,14.430671,14.703979,14.977287,15.250595,14.106606,12.96652,11.82253,10.67854,9.538455,9.245625,8.952794,8.659965,8.367134,8.074304,8.234385,8.39056,8.546737,8.706817,8.862993,8.488171,8.113348,7.7385254,7.363703,6.98888,7.1021075,7.2192397,7.3324676,7.445695,7.562827,7.1060123,6.649197,6.1884775,5.7316628,5.2748475,6.0244927,6.7702336,7.5159745,8.265619,9.01136,9.37447,9.737579,10.100689,10.4637985,10.826907,11.685876,12.544845,13.403813,14.2666855,15.125654,13.923099,12.720543,11.517986,10.315431,9.112875,10.518459,11.924045,13.325725,14.73131,16.136894,15.726933,15.31697,14.907008,14.4970455,14.087084,11.275913,8.468649,5.657479,2.8463092,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.6481308,1.1127546,1.5734742,2.0380979,2.4988174,4.6345253,6.7663293,8.898132,11.029937,13.16174,11.342289,9.522837,7.703386,5.883934,4.0605783,5.6926184,7.320754,8.952794,10.58093,12.212971,11.471134,10.729298,9.983557,9.24172,8.499884,14.079274,19.65476,25.234152,30.809639,36.38903,32.722794,29.056562,25.394232,21.727999,18.061766,16.339924,14.618082,12.89624,11.174399,9.448653,11.088503,12.724447,14.364296,16.00024,17.636185,16.09785,14.555612,13.017277,11.478943,9.936704,8.699008,7.461313,6.223617,4.985922,3.7482262,3.4710135,3.1898966,2.9087796,2.631567,2.35045,2.541766,2.7330816,2.9283018,3.1196175,3.310933,4.240181,5.169429,6.094772,7.0240197,7.9493628,6.676528,5.3997884,4.123049,2.8502135,1.5734742,1.261122,0.94876975,0.63641757,0.3240654,0.011713207,0.999527,1.475864,1.9482968,2.4246337,2.900971,3.3734035,6.3993154,9.425227,12.4511385,15.473146,18.499058,15.824542,13.150026,10.475512,7.800996,5.12648,4.474445,3.8263142,3.174279,2.5261483,1.8741131,4.689187,7.5003567,10.311526,13.1266,15.93777,13.688834,11.435994,9.187058,6.9381227,4.689187,10.373997,16.062712,21.751425,27.436235,33.12495,26.975515,20.826082,14.676648,8.52331,2.3738766,5.024966,7.676055,10.323239,12.974329,15.625418,23.438128,31.250835,39.063545,46.876255,54.68896,48.09833,41.511604,34.924877,28.338152,21.751425,17.761126,13.774731,9.788337,5.7980375,1.8116426,1.6242313,1.43682,1.2494087,1.0619974,0.8745861,0.74964523,0.62470436,0.4997635,0.37482262,0.24988174,1.4992905,2.7486992,3.998108,5.251421,6.5008297,5.4856853,4.474445,3.4632049,2.4480603,1.43682,3.513962,5.5871997,7.6643414,9.737579,11.810817,10.151445,8.488171,6.824895,5.1616197,3.4983444,3.6232853,3.7482262,3.873167,3.998108,4.123049,3.5256753,2.9243972,2.3231194,1.7257458,1.1244678,1.1869383,1.2494087,1.3118792,1.3743496,1.43682,3.2367494,5.036679,6.8366084,8.636538,10.436467,9.913278,9.386183,8.862993,8.335898,7.812709,8.663869,9.511124,10.362284,11.213444,12.0606985,11.150972,10.237343,9.323712,8.413987,7.5003567,7.7502384,8.00012,8.250002,8.499884,8.749765,11.974802,15.199838,18.424873,21.64991,24.874947,22.739239,20.599627,18.463919,16.324306,14.188598,11.873287,9.561881,7.250475,4.939069,2.6237583,2.436347,2.2489357,2.0615244,1.8741131,1.6867018,2.514435,3.338264,4.1620927,4.985922,5.813655,4.650143,3.4866312,2.3231194,1.1635119,0.0,2.0263848,4.0488653,6.0752497,8.101635,10.124115,8.101635,6.0752497,4.0488653,2.0263848,0.0,0.46071947,0.92534333,1.3860629,1.8506867,2.3114061,2.436347,2.5612879,2.6862288,2.8111696,2.9361105,5.2358036,7.535496,9.839094,12.138786,14.438479,12.361338,10.2881,8.210958,6.13772,4.0605783,3.6506162,3.2367494,2.8267872,2.4129205,1.999054,1.6515622,1.3001659,0.94876975,0.60127795,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.3357786,0.6754616,1.0112402,1.3509232,1.6867018,1.3743496,1.0619974,0.74964523,0.43729305,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.41386664,0.8238289,1.2376955,1.6515622,2.0615244,1.6749885,1.2884527,0.9019169,0.5114767,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26159495,0.5231899,0.78868926,1.0502841,1.3118792,1.2259823,1.1361811,1.0502841,0.96438736,0.8745861,0.698888,0.5231899,0.3513962,0.1756981,0.0,0.0,0.0,0.0,0.0,0.0,0.57394713,1.1517987,1.7257458,2.2996929,2.87364,2.338737,1.7999294,1.261122,0.7262188,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.13665408,0.27330816,0.41386664,0.5505207,0.6871748,0.81211567,0.93705654,1.0619974,1.1869383,1.3118792,1.2259823,1.1361811,1.0502841,0.96438736,0.8745861,0.9136301,0.94876975,0.9878138,1.0268579,1.0619974,1.175225,1.2884527,1.4016805,1.5110037,1.6242313,1.3626363,1.1010414,0.8355421,0.57394713,0.31235218,0.28892577,0.26159495,0.23816854,0.21083772,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.48805028,0.7262188,0.96438736,1.1986516,1.43682,2.2489357,3.0610514,3.873167,4.689187,5.5013027,4.900025,4.298747,3.7013733,3.1000953,2.4988174,2.1513257,1.7999294,1.4485333,1.1010414,0.74964523,0.9019169,1.0502841,1.1986516,1.3509232,1.4992905,1.3743496,1.2494087,1.1244678,0.999527,0.8745861,1.8623998,2.8502135,3.8380275,4.825841,5.813655,10.073358,14.336966,18.600573,22.86418,27.123882,22.723621,18.32336,13.923099,9.526741,5.12648,8.039165,10.951848,13.864532,16.773312,19.685997,16.074425,12.4628525,8.85128,5.2358036,1.6242313,6.7233806,11.826434,16.925583,22.024733,27.123882,21.700668,16.273548,10.850334,5.423215,0.0,0.42557985,0.8511597,1.2767396,1.698415,2.1239948,14.2901125,26.448421,38.61454,50.776752,62.938965,50.835316,38.73948,26.635832,14.53609,2.436347,5.1499066,7.8634663,10.577025,13.286681,16.00024,14.036326,12.076316,10.112402,8.148487,6.1884775,7.8868923,9.589212,11.287627,12.986042,14.688361,11.986515,9.288573,6.5867267,3.8887846,1.1869383,7.461313,13.735687,20.013966,26.28834,32.562714,27.123882,21.688955,16.250122,10.81129,5.376362,7.250475,9.124588,10.998701,12.8767185,14.750832,15.012426,15.274021,15.535617,15.801116,16.062712,14.700074,13.337439,11.974802,10.612165,9.249529,9.175345,9.101162,9.023073,8.94889,8.874706,9.187058,9.499411,9.811763,10.124115,10.436467,9.987461,9.538455,9.085544,8.636538,8.187531,8.300759,8.413987,8.52331,8.636538,8.749765,8.039165,7.3246584,6.6140575,5.899552,5.1889505,5.8761253,6.5633,7.250475,7.9376497,8.624825,9.43694,10.249056,11.061172,11.873287,12.689307,13.349152,14.012899,14.676648,15.336493,16.00024,14.53609,13.075843,11.611692,10.151445,8.687295,10.600452,12.513609,14.426766,16.33602,18.249176,17.226223,16.199366,15.176412,14.149553,13.1266,10.498938,7.8751793,5.251421,2.6237583,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,3.2757936,6.4891167,9.698535,12.911859,16.125181,13.013372,9.901564,6.785851,3.6740425,0.5622339,2.4012074,4.2362766,6.0752497,7.914223,9.749292,8.812236,7.8751793,6.9381227,6.001066,5.0640097,12.236397,19.412687,26.58898,33.761368,40.937656,36.29923,31.660797,27.026272,22.387842,17.749413,15.625418,13.501423,11.373524,9.249529,7.125534,9.6243515,12.127073,14.625891,17.124708,19.623526,17.686943,15.750359,13.813775,11.873287,9.936704,8.823949,7.7111945,6.5984397,5.4856853,4.376835,3.9746814,3.5764325,3.174279,2.77603,2.3738766,2.6237583,2.87364,3.1235218,3.3734035,3.6232853,4.388548,5.1499066,5.911265,6.676528,7.437886,6.2860875,5.138193,3.9863946,2.8385005,1.6867018,1.3509232,1.0112402,0.6754616,0.3357786,0.0,1.261122,1.7843118,2.3035975,2.822883,3.3421683,3.8614538,6.0713453,8.277332,10.48332,12.693212,14.899199,12.740065,10.58093,8.421796,6.2587566,4.0996222,3.68966,3.279698,2.8697357,2.4597735,2.0498111,4.298747,6.551587,8.800523,11.0494585,13.298394,11.838148,10.381805,8.921559,7.461313,6.001066,10.651209,15.3013525,19.951496,24.601639,29.251781,23.992552,18.733322,13.477997,8.218767,2.9634414,5.185046,7.406651,9.628256,11.8537655,14.07537,20.010061,25.944754,31.879444,37.814137,43.74883,38.595016,33.441204,28.28349,23.129679,17.975868,14.735214,11.49456,8.253906,5.0132523,1.7765031,1.7062237,1.639849,1.5734742,1.5031948,1.43682,1.2533131,1.0659018,0.8823949,0.698888,0.5114767,1.475864,2.4441557,3.408543,4.3729305,5.337318,4.618908,3.9044023,3.1859922,2.4675822,1.7491722,3.2992198,4.845363,6.3915067,7.941554,9.487698,8.277332,7.066968,5.8566036,4.646239,3.435874,3.8106966,4.1894236,4.564246,4.939069,5.3138914,4.942973,4.572055,4.2011366,3.8341231,3.4632049,3.174279,2.8892577,2.6003318,2.3114061,2.0263848,3.4514916,4.8765984,6.3017054,7.726812,9.151918,8.722435,8.296855,7.8673706,7.4417906,7.012306,7.7892823,8.566258,9.343235,10.124115,10.901091,10.05774,9.21439,8.371038,7.531592,6.688241,6.89127,7.098203,7.3012323,7.5081654,7.7111945,10.256865,12.802535,15.348206,17.893875,20.435642,19.026152,17.616663,16.207174,14.797685,13.388195,11.478943,9.565785,7.656533,5.74728,3.8380275,3.6349986,3.4319696,3.2289407,3.0259118,2.8267872,3.2992198,3.775557,4.251894,4.7243266,5.2006636,4.173806,3.1508527,2.1239948,1.1010414,0.07418364,1.6827974,3.2914112,4.8961205,6.504734,8.113348,6.4891167,4.8687897,3.2445583,1.6242313,0.0,0.37872702,0.76135844,1.1400855,1.5188124,1.901444,2.135708,2.3699722,2.6042364,2.8385005,3.076669,4.9468775,6.8209906,8.691199,10.565312,12.435521,11.217348,9.999174,8.777096,7.558923,6.336845,5.610626,4.884407,4.154284,3.4280653,2.7018464,2.2216048,1.7452679,1.2689307,0.78868926,0.31235218,0.30063897,0.28892577,0.27330816,0.26159495,0.24988174,0.46852827,0.6910792,0.9097257,1.1283722,1.3509232,1.1713207,0.9917182,0.80821127,0.62860876,0.44900626,0.359205,0.26940376,0.1796025,0.08980125,0.0,0.3318742,0.659844,0.9917182,1.319688,1.6515622,1.33921,1.0307622,0.71841,0.40996224,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.24597734,0.45681506,0.6676528,0.8784905,1.0893283,1.0112402,0.93315214,0.8550641,0.77697605,0.698888,0.5583295,0.42167544,0.28111696,0.14055848,0.0,0.0,0.0,0.0,0.0,0.0,0.46071947,0.92143893,1.3782539,1.8389735,2.2996929,1.8741131,1.4446288,1.0190489,0.58956474,0.1639849,0.13274968,0.10151446,0.07418364,0.042948425,0.011713207,0.12494087,0.23816854,0.3513962,0.46071947,0.57394713,0.6832704,0.79649806,0.9058213,1.0151446,1.1244678,1.0737107,1.0190489,0.96829176,0.9136301,0.8628729,0.97610056,1.0932326,1.2064602,1.3235924,1.43682,1.5500476,1.6632754,1.7765031,1.8858263,1.999054,1.6632754,1.3314011,0.9956226,0.659844,0.3240654,0.3513962,0.37872702,0.40605783,0.43338865,0.46071947,0.37872702,0.29673457,0.21474212,0.13274968,0.05075723,0.10932326,0.1639849,0.22255093,0.28111696,0.3357786,0.5036679,0.6715572,0.8394465,1.0073358,1.175225,1.8194515,2.463678,3.1118085,3.7560349,4.4002614,3.9239242,3.4514916,2.9751544,2.4988174,2.0263848,1.7452679,1.4641509,1.183034,0.9058213,0.62470436,0.78868926,0.94876975,1.1127546,1.2767396,1.43682,1.4016805,1.3626363,1.3235924,1.2884527,1.2494087,1.9365835,2.6237583,3.310933,3.998108,4.689187,8.101635,11.514082,14.92653,18.338978,21.751425,18.885593,16.019762,13.153932,10.2881,7.426173,10.202203,12.978233,15.758167,18.534197,21.314133,17.56981,13.829392,10.085071,6.3407493,2.6003318,6.4188375,10.241247,14.059752,17.878258,21.700668,17.37459,13.048512,8.726339,4.4002614,0.07418364,0.42557985,0.78088045,1.1322767,1.4836729,1.8389735,11.541413,21.247757,30.954102,40.65654,50.362885,40.726818,31.090755,21.458595,11.82253,2.1864653,4.337791,6.4891167,8.636538,10.787864,12.939189,13.887959,14.836729,15.789403,16.738173,17.686943,16.835783,15.984623,15.129559,14.278399,13.423335,11.521891,9.620447,7.719003,5.813655,3.912211,8.410083,12.907954,17.405825,21.903696,26.401567,22.875893,19.350218,15.824542,12.298867,8.773191,9.913278,11.0494585,12.185639,13.325725,14.461906,14.551707,14.641508,14.73131,14.821111,14.9109125,13.825488,12.743969,11.6585455,10.573121,9.487698,9.351044,9.21439,9.073831,8.937177,8.800523,9.081639,9.366661,9.647778,9.928895,10.213917,9.772718,9.331521,8.894228,8.453031,8.011833,8.800523,9.589212,10.373997,11.162686,11.951375,11.045554,10.139732,9.2339115,8.331994,7.426173,7.9454584,8.464745,8.98403,9.503315,10.0265045,10.436467,10.850334,11.2642,11.674163,12.08803,12.607315,13.1266,13.645885,14.169076,14.688361,13.591225,12.494087,11.393045,10.295909,9.198771,10.920613,12.63855,14.360392,16.07833,17.800169,16.640562,15.484859,14.329156,13.169549,12.013845,9.608734,7.2075267,4.806319,2.4012074,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,2.619854,5.1889505,7.7619514,10.331048,12.900145,10.48332,8.070399,5.6535745,3.240654,0.8238289,2.533957,4.2440853,5.9542136,7.6643414,9.37447,8.324185,7.2739015,6.223617,5.173333,4.123049,9.956225,15.789403,21.62258,27.455757,33.288933,30.762785,28.240541,25.718298,23.196054,20.67381,18.12814,15.586374,13.040704,10.495033,7.9493628,9.741484,11.533605,13.325725,15.12175,16.91387,15.617609,14.321347,13.028991,11.732729,10.436467,9.2221985,8.007929,6.79366,5.579391,4.3612175,3.998108,3.631094,3.2679846,2.900971,2.5378613,2.787743,3.0376248,3.2875066,3.5373883,3.78727,4.4119744,5.0327744,5.6535745,6.278279,6.899079,5.8175592,4.73604,3.6506162,2.5690966,1.4875772,1.1908426,0.8941081,0.59346914,0.29673457,0.0,1.5266213,2.0888553,2.6549935,3.2211318,3.7833657,4.349504,5.7394714,7.1294384,8.519405,9.909373,11.29934,9.655587,8.011833,6.364176,4.7204223,3.076669,2.9048753,2.7330816,2.5651922,2.3933985,2.2255092,3.912211,5.5989127,7.2856145,8.976221,10.662923,9.991365,9.323712,8.652155,7.9805984,7.3129454,10.924518,14.53609,18.151566,21.763138,25.37471,21.009588,16.644466,12.2793455,7.914223,3.5491016,5.3451266,7.141152,8.933272,10.729298,12.525322,16.581997,20.63867,24.69925,28.755922,32.812595,29.091702,25.366901,21.646006,17.921206,14.200311,11.709302,9.21439,6.7233806,4.2284675,1.737459,1.7882162,1.8428779,1.893635,1.9482968,1.999054,1.7530766,1.5110037,1.2650263,1.0190489,0.77307165,1.456342,2.135708,2.815074,3.49444,4.173806,3.7521305,3.330455,2.9087796,2.4831998,2.0615244,3.0805733,4.1035266,5.1225758,6.141625,7.1606736,6.4032197,5.645766,4.8883114,4.1308575,3.3734035,3.998108,4.6267166,5.251421,5.8761253,6.5008297,6.3602715,6.2197127,6.0791545,5.938596,5.801942,5.1616197,4.5252023,3.8887846,3.2484627,2.612045,3.6623292,4.7126136,5.7628975,6.813182,7.8634663,7.531592,7.2036223,6.871748,6.5437784,6.211904,6.918601,7.621393,8.32809,9.030883,9.737579,8.964508,8.191436,7.4183645,6.649197,5.8761253,6.036206,6.196286,6.356367,6.5164475,6.676528,8.538928,10.405232,12.271536,14.133936,16.00024,15.31697,14.633699,13.954333,13.271063,12.587793,11.080693,9.573594,8.066495,6.559396,5.0483923,4.83365,4.6150036,4.396357,4.181615,3.9629683,4.087909,4.21285,4.337791,4.462732,4.5876727,3.7013733,2.8111696,1.9248703,1.038571,0.14836729,1.33921,2.5300527,3.7208953,4.911738,6.098676,4.8805027,3.6584249,2.4402514,1.2181735,0.0,0.29673457,0.59346914,0.8941081,1.1908426,1.4875772,1.8311646,2.1786566,2.522244,2.8658314,3.213323,4.657952,6.1025805,7.5472097,8.991838,10.436467,10.073358,9.706344,9.343235,8.976221,8.6131115,7.570636,6.5281606,5.4856853,4.4432096,3.4007344,2.795552,2.1903696,1.5851873,0.98000497,0.37482262,0.39824903,0.42557985,0.44900626,0.47633708,0.4997635,0.60127795,0.7066968,0.80821127,0.9097257,1.0112402,0.96438736,0.91753453,0.8706817,0.8238289,0.77307165,0.62079996,0.46462387,0.30844778,0.15617609,0.0,0.24597734,0.4958591,0.7418364,0.9917182,1.2376955,1.0034313,0.77307165,0.5388075,0.30844778,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.23426414,0.39044023,0.5466163,0.7066968,0.8628729,0.79649806,0.7262188,0.659844,0.59346914,0.5231899,0.42167544,0.31625658,0.21083772,0.10541886,0.0,0.0,0.0,0.0,0.0,0.0,0.3435874,0.6910792,1.0346665,1.3782539,1.7257458,1.4055848,1.0893283,0.77307165,0.45681506,0.13665408,0.113227665,0.093705654,0.07027924,0.046852827,0.023426414,0.113227665,0.19912452,0.28892577,0.37482262,0.46071947,0.5583295,0.6520352,0.74574083,0.8433509,0.93705654,0.92143893,0.9019169,0.8862993,0.8667773,0.8511597,1.0424755,1.2337911,1.4290112,1.620327,1.8116426,1.9248703,2.0380979,2.1513257,2.260649,2.3738766,1.9678187,1.5617609,1.1517987,0.74574083,0.3357786,0.41777104,0.4958591,0.57785153,0.6559396,0.737932,0.60908675,0.48414588,0.3553006,0.22645533,0.10151446,0.1639849,0.23035973,0.29673457,0.359205,0.42557985,0.5231899,0.62079996,0.71841,0.8160201,0.9136301,1.3899672,1.8663043,2.3465457,2.822883,3.2992198,2.951728,2.6003318,2.2489357,1.901444,1.5500476,1.33921,1.1283722,0.92143893,0.7106012,0.4997635,0.6754616,0.8511597,1.0268579,1.1986516,1.3743496,1.4251068,1.475864,1.5266213,1.5734742,1.6242313,2.0107672,2.4012074,2.787743,3.174279,3.5608149,6.126007,8.687295,11.248583,13.813775,16.375063,15.043662,13.716166,12.384764,11.053363,9.725866,12.369146,15.008522,17.651802,20.295082,22.938364,19.065197,15.192029,11.318862,7.445695,3.5764325,6.114294,8.65606,11.193921,13.735687,16.273548,13.048512,9.823476,6.5984397,3.3734035,0.14836729,0.42948425,0.7106012,0.9917182,1.2689307,1.5500476,8.796618,16.043188,23.293663,30.540234,37.786804,30.618322,23.445936,16.277452,9.108971,1.9365835,3.5256753,5.1108627,6.699954,8.289046,9.874233,13.739592,17.601046,21.4625,25.323954,29.189312,25.780767,22.37613,18.97149,15.566852,12.162213,11.057267,9.952321,8.847376,7.7424297,6.6374836,9.358852,12.076316,14.797685,17.519053,20.236517,18.623999,17.01148,15.398962,13.786445,12.173926,12.576079,12.974329,13.376482,13.774731,14.176885,14.090988,14.008995,13.927003,13.845011,13.763018,12.954806,12.146595,11.338385,10.534078,9.725866,9.526741,9.323712,9.124588,8.925464,8.726339,8.976221,9.230007,9.483793,9.733675,9.987461,9.557977,9.128492,8.699008,8.265619,7.8361354,9.300286,10.760532,12.224684,13.688834,15.14908,14.051944,12.954806,11.85767,10.760532,9.663396,10.0147915,10.366188,10.721489,11.072885,11.424281,11.435994,11.4516115,11.4633255,11.475039,11.486752,11.8654785,12.244205,12.619028,12.997755,13.376482,12.642454,11.908427,11.178304,10.444276,9.714153,11.240774,12.767395,14.294017,15.820638,17.351164,16.058807,14.770353,13.481901,12.189544,10.901091,8.718531,6.5398736,4.3612175,2.1786566,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,1.9639144,3.892689,5.8214636,7.746334,9.675109,7.957172,6.239235,4.521298,2.803361,1.0893283,2.6706111,4.251894,5.833177,7.4183645,8.999647,7.8361354,6.676528,5.5130157,4.349504,3.1859922,7.676055,12.166118,16.65618,21.146242,25.636305,25.230247,24.82419,24.414227,24.00817,23.598207,20.634766,17.671324,14.703979,11.740538,8.773191,9.858616,10.944039,12.029464,13.114887,14.200311,13.548276,12.89624,12.244205,11.588266,10.936231,9.620447,8.300759,6.984976,5.6691923,4.349504,4.0215344,3.68966,3.3616903,3.0298162,2.7018464,2.951728,3.2016098,3.4514916,3.7013733,3.951255,4.4314966,4.9156423,5.395884,5.8800297,6.364176,5.349031,4.3338866,3.3187418,2.3035975,1.2884527,1.0307622,0.77307165,0.5153811,0.25769055,0.0,1.7882162,2.397303,3.0063896,3.619381,4.2284675,4.8375545,5.4115014,5.9815445,6.5554914,7.1294384,7.699481,6.571109,5.4388323,4.31046,3.1781836,2.0498111,2.1200905,2.1903696,2.260649,2.330928,2.4012074,3.5256753,4.650143,5.774611,6.899079,8.023546,8.144583,8.265619,8.386656,8.503788,8.624825,11.20173,13.774731,16.351637,18.924637,21.501543,18.026625,14.555612,11.080693,7.60968,4.138666,5.505207,6.871748,8.238289,9.608734,10.975275,13.153932,15.336493,17.515148,19.693806,21.876366,19.584482,17.296501,15.004618,12.716639,10.424754,8.679486,6.9342184,5.1889505,3.4436827,1.698415,1.8741131,2.0459068,2.2177005,2.3894942,2.5612879,2.2567444,1.9522011,1.6476578,1.3431144,1.038571,1.4329157,1.8272603,2.2216048,2.6159496,3.0141985,2.8853533,2.7565079,2.631567,2.5027218,2.3738766,2.8658314,3.3616903,3.853645,4.3455997,4.8375545,4.533011,4.2284675,3.9239242,3.619381,3.310933,4.1894236,5.0640097,5.938596,6.813182,7.687768,7.7775693,7.8673706,7.957172,8.046973,8.136774,7.1489606,6.1611466,5.173333,4.1894236,3.2016098,3.873167,4.548629,5.22409,5.899552,6.575013,6.3407493,6.1103897,5.8761253,5.645766,5.4115014,6.044015,6.676528,7.309041,7.941554,8.574067,7.871275,7.168483,6.46569,5.7668023,5.0640097,5.1772375,5.2943697,5.407597,5.520825,5.6379566,6.8209906,8.007929,9.190963,10.377901,11.560935,11.607788,11.650736,11.697589,11.744442,11.787391,10.682445,9.577498,8.472553,7.367607,6.262661,6.028397,5.7980375,5.563773,5.3334136,5.099149,4.8765984,4.650143,4.423688,4.2011366,3.9746814,3.2250361,2.475391,1.7257458,0.97610056,0.22645533,0.9956226,1.7686942,2.541766,3.3148375,4.087909,3.2718892,2.4519646,1.6359446,0.8160201,0.0,0.21474212,0.42948425,0.6442264,0.8589685,1.0737107,1.5305257,1.9834363,2.4402514,2.893162,3.349977,4.369026,5.3841705,6.4032197,7.4183645,8.437413,8.929368,9.4174185,9.909373,10.397423,10.889378,9.530646,8.171914,6.813182,5.4583545,4.0996222,3.3655949,2.6354716,1.901444,1.1713207,0.43729305,0.4997635,0.5622339,0.62470436,0.6871748,0.74964523,0.7340276,0.71841,0.7066968,0.6910792,0.6754616,0.76135844,0.8433509,0.92924774,1.0151446,1.1010414,0.8784905,0.659844,0.44119745,0.21864653,0.0,0.1639849,0.3318742,0.4958591,0.659844,0.8238289,0.6715572,0.5153811,0.359205,0.20693332,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.21864653,0.3240654,0.42557985,0.5309987,0.63641757,0.58175594,0.5231899,0.46462387,0.40605783,0.3513962,0.28111696,0.21083772,0.14055848,0.07027924,0.0,0.0,0.0,0.0,0.0,0.0,0.23035973,0.46071947,0.6910792,0.92143893,1.1517987,0.94096094,0.7340276,0.5270943,0.32016098,0.113227665,0.09761006,0.08199245,0.06637484,0.05075723,0.039044023,0.10151446,0.1639849,0.22645533,0.28892577,0.3513962,0.42948425,0.5114767,0.58956474,0.6715572,0.74964523,0.76916724,0.78478485,0.80430686,0.8199245,0.8394465,1.1088502,1.3782539,1.6476578,1.9170616,2.1864653,2.2996929,2.4129205,2.5261483,2.639376,2.7486992,2.2684577,1.7882162,1.3118792,0.8316377,0.3513962,0.48414588,0.61689556,0.74574083,0.8784905,1.0112402,0.8394465,0.6676528,0.4958591,0.3240654,0.14836729,0.22255093,0.29673457,0.3670138,0.44119745,0.5114767,0.5388075,0.5661383,0.59346914,0.62079996,0.6481308,0.96048295,1.2689307,1.5812829,1.8897307,2.1981785,1.9756275,1.7491722,1.5266213,1.3001659,1.0737107,0.93315214,0.79649806,0.6559396,0.5153811,0.37482262,0.5622339,0.74964523,0.93705654,1.1244678,1.3118792,1.4485333,1.5890918,1.7257458,1.8623998,1.999054,2.0888553,2.174752,2.260649,2.35045,2.436347,4.1503797,5.8644123,7.57454,9.288573,10.998701,11.205634,11.408664,11.615597,11.818625,12.025558,14.532186,17.03881,19.549341,22.05597,24.562595,20.560583,16.55857,12.556558,8.550641,4.548629,5.8097506,7.0708723,8.331994,9.589212,10.850334,8.726339,6.5984397,4.474445,2.35045,0.22645533,0.43338865,0.64032197,0.8472553,1.0541886,1.261122,6.0518236,10.8425255,15.633226,20.423927,25.210726,20.50592,15.801116,11.096312,6.3915067,1.6867018,2.7135596,3.736513,4.7633705,5.786324,6.813182,13.58732,20.361458,27.1395,33.91364,40.687775,34.729656,28.77154,22.813423,16.85921,10.901091,10.592644,10.284196,9.975748,9.671205,9.362757,10.303718,11.248583,12.189544,13.134409,14.07537,14.376009,14.676648,14.973383,15.274021,15.57466,15.238882,14.899199,14.56342,14.223738,13.887959,13.634172,13.376482,13.122696,12.86891,12.611219,12.084125,11.553126,11.022127,10.491129,9.964035,9.698535,9.43694,9.175345,8.913751,8.648251,8.870802,9.093353,9.315904,9.538455,9.761005,9.343235,8.921559,8.503788,8.082112,7.6643414,9.80005,11.935758,14.07537,16.211079,18.35069,17.058334,15.76988,14.481428,13.189071,11.900618,12.084125,12.271536,12.455043,12.63855,12.825961,12.435521,12.0489855,11.66245,11.275913,10.889378,11.123642,11.357906,11.592171,11.826434,12.0606985,11.693685,11.326671,10.959657,10.592644,10.22563,11.560935,12.89624,14.231546,15.566852,16.898252,15.477051,14.055848,12.630741,11.209538,9.788337,7.8283267,5.872221,3.9161155,1.9561055,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,1.3118792,2.5964274,3.8809757,5.165524,6.4500723,5.4310236,4.4119744,3.3890212,2.3699722,1.3509232,2.803361,4.2597027,5.716045,7.168483,8.624825,7.348085,6.0752497,4.7985106,3.5256753,2.2489357,5.395884,8.546737,11.693685,14.840633,17.987581,19.693806,21.403933,23.110157,24.816381,26.526508,23.141392,19.756275,16.371159,12.986042,9.600925,9.975748,10.354475,10.733202,11.111929,11.486752,11.478943,11.46723,11.45942,11.447707,11.435994,10.018696,8.597494,7.1762915,5.758993,4.337791,4.041056,3.7482262,3.4514916,3.1586614,2.8619268,3.1118085,3.3616903,3.611572,3.8614538,4.1113358,4.454923,4.7985106,5.138193,5.481781,5.825368,4.8765984,3.9317331,2.9829633,2.0341935,1.0893283,0.8706817,0.6520352,0.43338865,0.21864653,0.0,2.0498111,2.7057507,3.3616903,4.0137253,4.6696653,5.3256044,5.0796275,4.83365,4.591577,4.3455997,4.0996222,3.4866312,2.8697357,2.2567444,1.639849,1.0268579,1.3353056,1.6437533,1.9561055,2.2645533,2.5769055,3.1391394,3.7013733,4.263607,4.825841,5.388075,6.297801,7.2075267,8.117252,9.026978,9.936704,11.475039,13.013372,14.551707,16.086138,17.624472,15.043662,12.466757,9.885946,7.3051367,4.7243266,5.6652875,6.606249,7.5433054,8.484266,9.425227,9.725866,10.03041,10.331048,10.6355915,10.936231,10.081166,9.2221985,8.36323,7.5081654,6.649197,5.6535745,4.6540475,3.6584249,2.6588979,1.6632754,1.9561055,2.2489357,2.541766,2.8306916,3.1235218,2.7604125,2.3933985,2.0302892,1.6632754,1.3001659,1.4094892,1.5188124,1.6281357,1.7413634,1.8506867,2.018576,2.1864653,2.3543546,2.5183394,2.6862288,2.6510892,2.6159496,2.5808098,2.5456703,2.5105307,2.6588979,2.8072653,2.9556324,3.1039999,3.2484627,4.376835,5.5013027,6.6257706,7.7502384,8.874706,9.194867,9.515028,9.835189,10.155351,10.475512,9.136301,7.800996,6.461786,5.12648,3.78727,4.087909,4.388548,4.689187,4.985922,5.2865605,5.153811,5.017157,4.884407,4.747753,4.6110992,5.173333,5.7316628,6.2938967,6.852226,7.4105554,6.7780423,6.1494336,5.5130157,4.884407,4.251894,4.318269,4.388548,4.4588275,4.5291066,4.5993857,5.1030536,5.610626,6.114294,6.621866,7.125534,7.898606,8.671678,9.440845,10.213917,10.986988,10.284196,9.581403,8.878611,8.175818,7.47693,7.2270484,6.9810715,6.7311897,6.4852123,6.239235,5.661383,5.087436,4.513489,3.9356375,3.3616903,2.7486992,2.135708,1.5266213,0.9136301,0.30063897,0.6559396,1.0112402,1.3665408,1.7218413,2.0732377,1.6593709,1.2455044,0.8316377,0.41386664,0.0,0.13274968,0.26549935,0.39824903,0.5309987,0.6637484,1.2259823,1.7921207,2.358259,2.9243972,3.4866312,4.0761957,4.6657605,5.2592297,5.8487945,6.4383593,7.7814736,9.128492,10.471607,11.818625,13.16174,11.490656,9.815667,8.144583,6.473499,4.7985106,3.9395418,3.0805733,2.2216048,1.358732,0.4997635,0.60127795,0.698888,0.80040246,0.9019169,0.999527,0.8667773,0.7340276,0.60127795,0.46852827,0.3357786,0.5544251,0.77307165,0.9917182,1.2064602,1.4251068,1.1400855,0.8550641,0.5700427,0.28502136,0.0,0.08199245,0.1639849,0.24597734,0.3318742,0.41386664,0.3357786,0.25769055,0.1796025,0.10151446,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.20302892,0.25378615,0.30844778,0.359205,0.41386664,0.3631094,0.31625658,0.26940376,0.22255093,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.0,0.0,0.0,0.0,0.0,0.113227665,0.23035973,0.3435874,0.46071947,0.57394713,0.47633708,0.37872702,0.28111696,0.1835069,0.08589685,0.078088045,0.07418364,0.06637484,0.058566034,0.05075723,0.08589685,0.12494087,0.1639849,0.19912452,0.23816854,0.30063897,0.3670138,0.43338865,0.4958591,0.5622339,0.61689556,0.6676528,0.71841,0.77307165,0.8238289,1.1713207,1.5188124,1.8663043,2.2137961,2.5612879,2.6745155,2.787743,2.900971,3.0141985,3.1235218,2.5730011,2.018576,1.4680552,0.9136301,0.3631094,0.5466163,0.7340276,0.91753453,1.1010414,1.2884527,1.0698062,0.8511597,0.63641757,0.41777104,0.19912452,0.28111696,0.359205,0.44119745,0.5192855,0.60127795,0.5583295,0.5153811,0.47243267,0.42948425,0.38653582,0.5309987,0.6715572,0.8160201,0.95657855,1.1010414,0.999527,0.9019169,0.80040246,0.698888,0.60127795,0.5309987,0.46071947,0.39044023,0.32016098,0.24988174,0.44900626,0.6481308,0.8511597,1.0502841,1.2494087,1.475864,1.698415,1.9248703,2.1513257,2.3738766,2.1630387,1.9482968,1.737459,1.5266213,1.3118792,2.174752,3.0376248,3.900498,4.7633705,5.6262436,7.363703,9.105066,10.84643,12.583888,14.325252,16.69913,19.069101,21.442978,23.816854,26.186827,22.05597,17.921206,13.790349,9.655587,5.5247293,5.505207,5.4856853,5.466163,5.446641,5.423215,4.4002614,3.3734035,2.35045,1.3235924,0.30063897,0.43338865,0.5700427,0.7066968,0.8394465,0.97610056,3.3070288,5.6379566,7.9727893,10.303718,12.63855,10.397423,8.156297,5.919074,3.677947,1.43682,1.901444,2.3621633,2.8267872,3.2875066,3.7482262,13.438952,23.125774,32.812595,42.49942,52.18624,43.678547,35.16695,26.655354,18.147661,9.636065,10.128019,10.61607,11.108025,11.596075,12.08803,11.252487,10.416945,9.581403,8.745861,7.914223,10.124115,12.337912,14.551707,16.761599,18.975395,17.901684,16.82407,15.750359,14.676648,13.599033,13.173453,12.743969,12.318389,11.888905,11.4633255,11.209538,10.955752,10.705871,10.452085,10.198298,9.874233,9.550168,9.226103,8.898132,8.574067,8.769287,8.960603,9.151918,9.343235,9.538455,9.128492,8.718531,8.308568,7.898606,7.4886436,10.299813,13.110983,15.926057,18.737226,21.548395,20.068628,18.584955,17.101282,15.621513,14.13784,14.153459,14.17298,14.188598,14.208119,14.223738,13.438952,12.650263,11.861574,11.076789,10.2881,10.381805,10.471607,10.565312,10.6590185,10.748819,10.748819,10.744915,10.741011,10.741011,10.737106,11.881096,13.021181,14.165172,15.309161,16.449247,14.895294,13.341343,11.783486,10.229534,8.675582,6.9381227,5.2045684,3.4710135,1.7335546,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.6559396,1.2962615,1.9404879,2.5808098,3.2250361,2.900971,2.5808098,2.2567444,1.9365835,1.6125181,2.9400148,4.267512,5.5950084,6.9225054,8.250002,6.8639393,5.473972,4.087909,2.7018464,1.3118792,3.1157131,4.9234514,6.727285,8.531119,10.338858,14.161267,17.983677,21.806087,25.628496,29.450907,25.644114,21.841227,18.034433,14.231546,10.424754,10.096785,9.76491,9.433036,9.105066,8.773191,9.405705,10.0382185,10.670732,11.303245,11.935758,10.413041,8.894228,7.3715115,5.8487945,4.3260775,4.0644827,3.8067923,3.5451972,3.2836022,3.0259118,3.2757936,3.5256753,3.775557,4.025439,4.2753205,4.478349,4.6813784,4.884407,5.083532,5.2865605,4.40807,3.5256753,2.6471848,1.7686942,0.8862993,0.7106012,0.5309987,0.3553006,0.1756981,0.0,2.3114061,3.0141985,3.7130866,4.4119744,5.1108627,5.813655,4.7516575,3.6857557,2.6237583,1.5617609,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.5505207,1.1010414,1.6515622,2.1981785,2.7486992,2.7486992,2.7486992,2.7486992,2.7486992,2.7486992,4.4510183,6.1494336,7.8517528,9.550168,11.248583,11.748346,12.24811,12.751778,13.251541,13.751305,12.0606985,10.373997,8.687295,7.000593,5.3138914,5.825368,6.336845,6.8483214,7.363703,7.8751793,6.3017054,4.7243266,3.1508527,1.5734742,0.0,0.57394713,1.1517987,1.7257458,2.2996929,2.87364,2.6237583,2.3738766,2.1239948,1.8741131,1.6242313,2.0380979,2.4480603,2.8619268,3.2757936,3.6857557,3.2640803,2.8385005,2.4129205,1.9873407,1.5617609,1.3860629,1.2142692,1.038571,0.8628729,0.6871748,1.1517987,1.6125181,2.0732377,2.5378613,2.998581,2.436347,1.8741131,1.3118792,0.74964523,0.18741131,0.78868926,1.3860629,1.9873407,2.5886188,3.1859922,4.564246,5.938596,7.3129454,8.687295,10.061645,10.612165,11.162686,11.713207,12.263727,12.814248,11.123642,9.43694,7.7502384,6.0635366,4.376835,4.298747,4.224563,4.1503797,4.0761957,3.998108,3.9629683,3.9239242,3.8887846,3.8497405,3.8106966,4.298747,4.786797,5.2748475,5.7628975,6.250948,5.688714,5.12648,4.564246,3.998108,3.435874,3.4632049,3.4866312,3.513962,3.5373883,3.5608149,3.3890212,3.213323,3.0376248,2.8619268,2.6862288,4.1894236,5.688714,7.1880045,8.687295,10.186585,9.885946,9.589212,9.288573,8.987934,8.687295,8.4257,8.164105,7.898606,7.6370106,7.375416,6.4500723,5.5247293,4.5993857,3.6740425,2.7486992,2.2762666,1.7999294,1.3235924,0.8511597,0.37482262,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.92534333,1.6008049,2.2762666,2.951728,3.6232853,3.78727,3.951255,4.1113358,4.2753205,4.4393053,6.6374836,8.835662,11.037745,13.235924,15.438006,13.450665,11.4633255,9.475985,7.4886436,5.5013027,4.513489,3.5256753,2.5378613,1.5500476,0.5622339,0.698888,0.8394465,0.97610056,1.1127546,1.2494087,0.999527,0.74964523,0.4997635,0.24988174,0.0,0.3513962,0.698888,1.0502841,1.4016805,1.7491722,1.4016805,1.0502841,0.698888,0.3513962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.1756981,0.22645533,0.27330816,0.3240654,0.37482262,0.46071947,0.5505207,0.63641757,0.7262188,0.81211567,1.2376955,1.6632754,2.0888553,2.514435,2.9361105,3.049338,3.1625657,3.2757936,3.3890212,3.4983444,2.87364,2.2489357,1.6242313,0.999527,0.37482262,0.61299115,0.8511597,1.0893283,1.3235924,1.5617609,1.3001659,1.038571,0.77307165,0.5114767,0.24988174,0.3357786,0.42557985,0.5114767,0.60127795,0.6871748,0.57394713,0.46071947,0.3513962,0.23816854,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.3357786,0.5505207,0.76135844,0.97610056,1.1869383,1.4992905,1.8116426,2.1239948,2.436347,2.7486992,2.2372224,1.7257458,1.2142692,0.698888,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,3.5256753,6.801469,10.073358,13.349152,16.624945,18.862167,21.09939,23.336613,25.573835,27.811058,23.551353,19.287746,15.024139,10.760532,6.5008297,5.2006636,3.900498,2.6003318,1.3001659,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.43729305,0.4997635,0.5622339,0.62470436,0.6871748,0.5622339,0.43729305,0.31235218,0.18741131,0.062470436,0.28892577,0.5114767,0.737932,0.96438736,1.1869383,1.0893283,0.9878138,0.8862993,0.78868926,0.6871748,13.286681,25.886187,38.489597,51.089104,63.68861,52.623535,41.562363,30.50119,19.436115,8.374943,9.663396,10.951848,12.236397,13.524849,14.813302,12.201257,9.589212,6.9732623,4.3612175,1.7491722,5.8761253,9.999174,14.126127,18.249176,22.37613,20.560583,18.74894,16.937298,15.125654,13.314012,12.712734,12.111456,11.514082,10.912805,10.311526,10.338858,10.362284,10.38571,10.413041,10.436467,10.049932,9.663396,9.276859,8.886419,8.499884,8.663869,8.823949,8.987934,9.151918,9.311999,8.913751,8.511597,8.113348,7.7111945,7.3129454,10.799577,14.286208,17.776743,21.263374,24.750006,23.075018,21.400028,5052.0,18.05005,16.375063,16.226696,16.074425,15.926057,15.773785,15.625418,14.438479,13.251541,12.0606985,10.87376,9.686822,9.636065,9.589212,9.538455,9.487698,9.43694,9.80005,10.163159,10.526268,10.889378,11.248583,12.201257,13.150026,14.098797,15.051471,16.00024,14.313539,12.626837,10.936231,9.249529,7.562827,6.0518236,4.5369153,3.0259118,1.5110037,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.37482262,0.74964523,1.1244678,1.4992905,1.8741131,3.076669,4.2753205,5.473972,6.676528,7.8751793,6.375889,4.8765984,3.3734035,1.8741131,0.37482262,0.8394465,1.3001659,1.7608855,2.2255092,2.6862288,8.624825,14.56342,20.502016,26.436708,32.375305,28.15074,23.926178,19.701614,15.477051,11.248583,10.213917,9.175345,8.136774,7.098203,6.0635366,7.336372,8.6131115,9.885946,11.162686,12.439425,10.81129,9.187058,7.562827,5.938596,4.3143644,4.087909,3.8614538,3.638903,3.4124475,3.1859922,3.435874,3.6857557,3.9356375,4.1894236,4.4393053,4.5017757,4.564246,4.6267166,4.689187,4.7516575,3.9356375,3.1235218,2.3114061,1.4992905,0.6871748,0.5505207,0.41386664,0.27330816,0.13665408,0.0,1.8506867,2.4090161,2.97125,3.5295796,4.0918136,4.650143,4.3612175,4.068387,3.7794614,3.4905357,3.2016098,3.506153,3.814601,4.123049,4.4314966,4.73604,4.970304,5.2006636,5.434928,5.6691923,5.899552,6.364176,6.824895,7.289519,7.7502384,8.210958,9.60483,10.998701,12.388668,13.78254,15.176412,14.34087,13.505327,12.6697855,11.834243,10.998701,9.655587,8.308568,6.9654536,5.618435,4.2753205,4.6852827,5.095245,5.505207,5.9151692,6.3251314,5.3060827,4.290938,3.2718892,2.2567444,1.2376955,1.4953861,1.7530766,2.0107672,2.2684577,2.5261483,2.280171,2.0341935,1.7882162,1.5461433,1.3001659,1.6281357,1.9600099,2.2918842,2.619854,2.951728,2.9829633,3.0141985,3.049338,3.0805733,3.1118085,2.6042364,2.0927596,1.5812829,1.0737107,0.5622339,1.0737107,1.5812829,2.0927596,2.6042364,3.1118085,2.631567,2.1474214,1.6632754,1.183034,0.698888,1.0932326,1.4836729,1.8780174,2.2684577,2.6628022,3.814601,4.9663997,6.1181984,7.2739015,8.4257,8.894228,9.358852,9.82738,10.295909,10.760532,9.612638,8.460839,7.3129454,6.1611466,5.0132523,5.02887,5.040583,5.056201,5.0718184,5.087436,5.2592297,5.4271193,5.5989127,5.7668023,5.938596,6.0713453,6.2079997,6.3407493,6.477403,6.6140575,6.3017054,5.9932575,5.6809053,5.3724575,5.0640097,4.93126,4.802415,4.6735697,4.5408196,4.4119744,3.998108,3.5842414,3.1664703,2.7526035,2.338737,3.5725281,4.806319,6.044015,7.277806,8.511597,8.261715,8.007929,7.7541428,7.504261,7.250475,7.363703,7.480835,7.5940623,7.7111945,7.824422,7.152865,6.481308,5.805846,5.134289,4.462732,3.8106966,3.1586614,2.5066261,1.8506867,1.1986516,1.0698062,0.94096094,0.80821127,0.679366,0.5505207,0.46071947,0.3709182,0.28111696,0.19131571,0.10151446,0.14446288,0.19131571,0.23426414,0.28111696,0.3240654,0.9058213,1.4836729,2.0654287,2.6432803,3.2250361,3.3812122,3.541293,3.697469,3.853645,4.0137253,5.8956475,7.7814736,9.6673,11.553126,13.438952,11.931853,10.4286585,8.921559,7.4183645,5.911265,4.8765984,3.8380275,2.7994564,1.7608855,0.7262188,0.8238289,0.92534333,1.0268579,1.1244678,1.2259823,0.98390937,0.7418364,0.4958591,0.25378615,0.011713207,0.339683,0.6676528,0.9956226,1.3235924,1.6515622,1.3860629,1.1244678,0.8628729,0.60127795,0.3357786,0.26940376,0.20302892,0.13665408,0.06637484,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.14836729,0.14836729,0.14836729,0.14836729,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.058566034,0.07027924,0.078088045,0.08980125,0.10151446,0.14836729,0.19522011,0.24207294,0.28892577,0.3357786,0.6520352,0.96829176,1.2806439,1.5969005,1.9131571,2.0341935,2.1591344,2.280171,2.4012074,2.5261483,2.6237583,2.7252727,2.8267872,2.9243972,3.0259118,2.4792955,1.9365835,1.3899672,0.8433509,0.30063897,0.48805028,0.679366,0.8706817,1.0580931,1.2494087,1.0463798,0.8394465,0.63641757,0.42948425,0.22645533,0.29283017,0.359205,0.42557985,0.4958591,0.5622339,0.47243267,0.38263142,0.29283017,0.20302892,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.10151446,0.10541886,0.10932326,0.10932326,0.113227665,0.30063897,0.49195468,0.6832704,0.8706817,1.0619974,1.3040704,1.542239,1.7843118,2.0224805,2.260649,1.8389735,1.4172981,0.9956226,0.57394713,0.14836729,0.16008049,0.1717937,0.1796025,0.19131571,0.19912452,2.8189783,5.4388323,8.058686,10.67854,13.298394,15.223265,17.148134,19.07691,21.00178,22.926651,19.561056,16.195461,12.829865,9.464272,6.098676,4.8805027,3.6584249,2.4402514,1.2181735,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.3513962,0.39824903,0.44900626,0.4997635,0.5505207,0.45291066,0.3553006,0.25769055,0.16008049,0.062470436,0.24597734,0.42557985,0.60908675,0.79259366,0.97610056,1.1713207,1.3665408,1.5617609,1.7530766,1.9482968,12.154405,22.360512,32.56662,42.76882,52.97493,43.76835,34.565674,25.359093,16.156416,6.949836,8.117252,9.284669,10.452085,11.619501,12.786918,14.774258,16.761599,18.74894,20.73628,22.723621,22.247284,21.767042,21.2868,20.80656,20.326319,19.162806,17.999294,16.835783,15.676175,14.512663,13.696643,12.8767185,12.0606985,11.240774,10.424754,10.292005,10.159255,10.0265045,9.893755,9.761005,9.190963,8.617016,8.043069,7.473026,6.899079,7.1880045,7.473026,7.7619514,8.050878,8.335898,8.140678,7.941554,7.746334,7.5472097,7.348085,10.229534,13.110983,15.988527,18.869976,21.751425,20.498112,19.244799,17.991486,16.738173,15.488764,15.262308,15.035853,14.813302,14.586847,14.364296,13.645885,12.93138,12.216875,11.502369,10.787864,10.791768,10.791768,10.795672,10.795672,10.799577,11.057267,11.314958,11.572648,11.8303385,12.08803,12.236397,12.380859,12.529227,12.677594,12.825961,11.510178,10.194394,8.878611,7.5667315,6.250948,5.001539,3.7482262,2.4988174,1.2494087,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07027924,0.14055848,0.21083772,0.28111696,0.3513962,0.28111696,0.21083772,0.14055848,0.07027924,0.0,0.0,0.0,0.0,0.0,0.0,0.30063897,0.60127795,0.9019169,1.1986516,1.4992905,2.6081407,3.7130866,4.8219366,5.930787,7.0357327,5.786324,4.5369153,3.2875066,2.0380979,0.78868926,1.0580931,1.3314011,1.6047094,1.8780174,2.1513257,7.008402,11.869383,16.730364,21.591345,26.448421,23.906654,21.360985,18.815315,16.269644,13.723974,12.181735,10.639496,9.097258,7.5550184,6.012779,7.3012323,8.59359,9.882042,11.170495,12.4628525,10.756628,9.0465,7.3402762,5.6340523,3.9239242,3.6623292,3.4007344,3.1391394,2.87364,2.612045,2.8306916,3.049338,3.2640803,3.4827268,3.7013733,3.7208953,3.7404175,3.7599394,3.7794614,3.7989833,3.1508527,2.4988174,1.8506867,1.1986516,0.5505207,0.44119745,0.3318742,0.21864653,0.10932326,0.0,1.3860629,1.8077383,2.2294137,2.6471848,3.06886,3.4866312,3.970777,4.4510183,4.9351645,5.4193106,5.899552,6.6140575,7.328563,8.046973,8.761478,9.475985,9.390087,9.304191,9.218294,9.136301,9.050405,9.975748,10.901091,11.826434,12.751778,13.673217,14.75864,15.844065,16.92949,18.014912,19.100336,16.92949,14.75864,12.591698,10.42085,8.250002,7.2465706,6.2431393,5.2436123,4.240181,3.2367494,3.5451972,3.853645,4.1581883,4.466636,4.775084,4.3143644,3.853645,3.39683,2.9361105,2.475391,2.416825,2.3543546,2.2957885,2.233318,2.174752,1.9365835,1.6945106,1.456342,1.2142692,0.97610056,1.2220778,1.4680552,1.717937,1.9639144,2.2137961,2.7018464,3.193801,3.6818514,4.173806,4.661856,3.8185053,2.97125,2.1278992,1.2806439,0.43729305,0.9956226,1.5539521,2.1083772,2.6667068,3.2250361,2.822883,2.4207294,2.018576,1.6164225,1.2142692,1.397776,1.5812829,1.7686942,1.9522011,2.135708,3.06886,3.998108,4.927356,5.8566036,6.785851,7.172387,7.558923,7.941554,8.32809,8.710721,8.101635,7.4886436,6.8756523,6.262661,5.64967,5.755089,5.860508,5.9659266,6.0713453,6.1767645,6.551587,6.930314,7.309041,7.6838636,8.062591,7.843944,7.629202,7.4105554,7.191909,6.9732623,6.918601,6.860035,6.801469,6.746807,6.688241,6.4032197,6.1181984,5.833177,5.548156,5.263134,4.607195,3.951255,3.2992198,2.6432803,1.9873407,2.9556324,3.9278288,4.8961205,5.8683167,6.8366084,6.6335793,6.426646,6.223617,6.016684,5.813655,6.3056097,6.7975645,7.289519,7.7814736,8.273428,7.8556576,7.433982,7.016211,6.5945354,6.1767645,5.3451266,4.513489,3.6857557,2.854118,2.0263848,1.8272603,1.6281357,1.4329157,1.2337911,1.038571,0.8706817,0.7027924,0.5349031,0.3670138,0.19912452,0.23816854,0.28111696,0.32016098,0.359205,0.39824903,0.8862993,1.3704453,1.8545911,2.338737,2.8267872,2.979059,3.1313305,3.2836022,3.435874,3.5881457,5.1577153,6.727285,8.296855,9.866425,11.435994,10.416945,9.393991,8.371038,7.348085,6.3251314,5.2358036,4.1503797,3.0610514,1.9756275,0.8862993,0.94876975,1.0112402,1.0737107,1.1361811,1.1986516,0.96438736,0.7301232,0.4958591,0.26159495,0.023426414,0.3318742,0.63641757,0.94096094,1.2455044,1.5500476,1.3743496,1.1986516,1.0268579,0.8511597,0.6754616,0.5388075,0.40605783,0.26940376,0.13665408,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.113227665,0.113227665,0.113227665,0.113227665,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.046852827,0.05075723,0.058566034,0.06637484,0.07418364,0.12103647,0.1639849,0.21083772,0.25378615,0.30063897,0.8433509,1.3860629,1.9287747,2.4714866,3.0141985,2.8306916,2.6510892,2.4714866,2.2918842,2.1122816,2.1981785,2.2879796,2.3738766,2.463678,2.5495746,2.084951,1.620327,1.1557031,0.6910792,0.22645533,0.3670138,0.5114767,0.6520352,0.79649806,0.93705654,0.78868926,0.6442264,0.4958591,0.3474918,0.19912452,0.24597734,0.29673457,0.3435874,0.39044023,0.43729305,0.3709182,0.30063897,0.23426414,0.1678893,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.078088045,0.08589685,0.08980125,0.093705654,0.10151446,0.26940376,0.43338865,0.60127795,0.76916724,0.93705654,1.1049459,1.2728351,1.4407244,1.6086137,1.7765031,1.4407244,1.1088502,0.77697605,0.44510186,0.113227665,0.12103647,0.12884527,0.13665408,0.14055848,0.14836729,2.1161861,4.0801005,6.044015,8.011833,9.975748,11.588266,13.200784,14.813302,16.42582,18.038338,15.570756,13.103174,10.6355915,8.16801,5.700427,4.560342,3.4202564,2.280171,1.1400855,0.0,0.046852827,0.08980125,0.13665408,0.1796025,0.22645533,0.26159495,0.30063897,0.3357786,0.37482262,0.41386664,0.3435874,0.27330816,0.20302892,0.13274968,0.062470436,0.20302892,0.3435874,0.48414588,0.62079996,0.76135844,1.2533131,1.7413634,2.233318,2.7213683,3.213323,11.022127,18.830933,26.64364,34.452446,42.26125,34.913166,27.568985,20.2209,12.872814,5.5247293,6.571109,7.621393,8.667773,9.714153,10.764437,17.351164,23.937891,30.524616,37.111343,43.701973,38.61454,33.531006,28.443571,23.360039,18.276506,17.761126,17.24965,16.738173,16.226696,15.711315,14.676648,13.641981,12.607315,11.572648,10.537982,10.249056,9.956225,9.6673,9.378374,9.085544,8.32809,7.570636,6.813182,6.055728,5.298274,5.7121406,6.126007,6.5359693,6.949836,7.363703,7.367607,7.3715115,7.37932,7.3832245,7.387129,9.659492,11.931853,14.204215,16.476578,18.74894,17.921206,17.08957,16.261835,15.430198,14.59856,14.301826,14.001186,13.700547,13.399908,13.09927,12.857197,12.615124,12.373051,12.130978,11.888905,11.943566,11.998228,12.05289,12.107552,12.162213,12.314485,12.466757,12.619028,12.771299,12.923572,12.271536,11.615597,10.959657,10.303718,9.651682,8.706817,7.7658563,6.8209906,5.8800297,4.939069,3.951255,2.9634414,1.9756275,0.9878138,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14055848,0.28111696,0.42167544,0.5583295,0.698888,0.5583295,0.42167544,0.28111696,0.14055848,0.0,0.0,0.0,0.0,0.0,0.0,0.22645533,0.44900626,0.6754616,0.9019169,1.1244678,2.1396124,3.154757,4.169902,5.185046,6.2001905,5.2006636,4.2011366,3.2016098,2.1981785,1.1986516,1.2806439,1.3665408,1.4485333,1.5305257,1.6125181,5.395884,9.17925,12.958711,16.742077,20.525442,19.658665,18.795792,17.929016,17.066143,16.199366,14.153459,12.103647,10.05774,8.011833,5.9620223,7.266093,8.574067,9.878138,11.182208,12.486279,10.698062,8.905942,7.1177254,5.3295093,3.5373883,3.2367494,2.9361105,2.639376,2.338737,2.0380979,2.2216048,2.4090161,2.592523,2.77603,2.9634414,2.9400148,2.9165885,2.893162,2.87364,2.8502135,2.3621633,1.8741131,1.3860629,0.9019169,0.41386664,0.3318742,0.24597734,0.1639849,0.08199245,0.0,0.92534333,1.2064602,1.4836729,1.7647898,2.0459068,2.3231194,3.5803368,4.83365,6.0908675,7.3441806,8.601398,9.721962,10.84643,11.966993,13.091461,14.212025,13.809871,13.407718,13.005564,12.603411,12.201257,13.58732,14.973383,16.36335,17.749413,19.13938,19.916355,20.693333,21.470308,22.247284,23.02426,19.518106,16.015858,12.509705,9.0035515,5.5013027,4.841459,4.181615,3.521771,2.8619268,2.1981785,2.4051118,2.6081407,2.815074,3.018103,3.2250361,3.3226464,3.4202564,3.5178664,3.6154766,3.7130866,3.3343596,2.9556324,2.5808098,2.2020829,1.8233559,1.5890918,1.3548276,1.1205635,0.8862993,0.6481308,0.8160201,0.98000497,1.1439898,1.3118792,1.475864,2.4207294,3.3694992,4.318269,5.263134,6.211904,5.0327744,3.853645,2.6706111,1.4914817,0.31235218,0.91753453,1.5227169,2.1278992,2.7330816,3.338264,3.0141985,2.6940374,2.3699722,2.0459068,1.7257458,1.7023194,1.678893,1.6593709,1.6359446,1.6125181,2.3192148,3.0259118,3.736513,4.4432096,5.1499066,5.45445,5.755089,6.055728,6.3602715,6.66091,6.5867267,6.5125427,6.4383593,6.364176,6.2860875,6.481308,6.676528,6.871748,7.066968,7.262188,7.8478484,8.433509,9.019169,9.600925,10.186585,9.616543,9.0465,8.476458,7.9064145,7.336372,7.531592,7.726812,7.9220324,8.117252,8.312472,7.871275,7.433982,6.9927845,6.551587,6.114294,5.2162814,4.322173,3.4280653,2.533957,1.6359446,2.3426414,3.049338,3.7521305,4.4588275,5.1616197,5.0054436,4.8492675,4.689187,4.533011,4.376835,5.2436123,6.114294,6.984976,7.8556576,8.726339,8.55845,8.39056,8.2226715,8.054782,7.8868923,6.8795567,5.872221,4.8648853,3.8575494,2.8502135,2.5847144,2.3192148,2.0537157,1.7882162,1.5266213,1.2806439,1.0346665,0.78868926,0.5466163,0.30063897,0.3357786,0.3709182,0.40605783,0.44119745,0.47633708,0.8667773,1.2533131,1.6437533,2.0341935,2.4246337,2.5730011,2.7213683,2.8658314,3.0141985,3.1625657,4.415879,5.6730967,6.9264097,8.183627,9.43694,8.898132,8.359325,7.816613,7.277806,6.7389984,5.5989127,4.462732,3.3265507,2.1864653,1.0502841,1.0737107,1.1010414,1.1244678,1.1517987,1.175225,0.94876975,0.71841,0.49195468,0.26549935,0.039044023,0.32016098,0.60127795,0.8862993,1.1674163,1.4485333,1.3626363,1.2767396,1.1869383,1.1010414,1.0112402,0.80821127,0.60908675,0.40605783,0.20302892,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.031235218,0.03513962,0.039044023,0.046852827,0.05075723,0.093705654,0.13665408,0.1756981,0.21864653,0.26159495,1.0307622,1.8038338,2.5730011,3.3421683,4.1113358,3.631094,3.1469483,2.6667068,2.182561,1.698415,1.7765031,1.8506867,1.9248703,1.999054,2.0732377,1.6906061,1.3040704,0.92143893,0.5349031,0.14836729,0.24597734,0.339683,0.43338865,0.5309987,0.62470436,0.5349031,0.44510186,0.3553006,0.26549935,0.1756981,0.20302892,0.23035973,0.25769055,0.28502136,0.31235218,0.26940376,0.22255093,0.1756981,0.13274968,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.058566034,0.06637484,0.07418364,0.078088045,0.08589685,0.23426414,0.37872702,0.5231899,0.6676528,0.81211567,0.9058213,1.0034313,1.097137,1.1908426,1.2884527,1.0463798,0.80430686,0.5583295,0.31625658,0.07418364,0.078088045,0.08589685,0.08980125,0.093705654,0.10151446,1.4094892,2.7213683,4.029343,5.3412223,6.649197,7.9493628,9.249529,10.549695,11.849861,13.150026,11.580457,10.010887,8.441318,6.871748,5.298274,4.240181,3.1781836,2.1200905,1.0580931,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.1756981,0.19912452,0.22645533,0.24988174,0.27330816,0.23426414,0.19131571,0.14836729,0.10541886,0.062470436,0.16008049,0.25769055,0.3553006,0.45291066,0.5505207,1.3353056,2.1200905,2.9048753,3.68966,4.474445,9.889851,15.305257,20.720663,26.136068,31.551476,26.057981,20.568392,15.078801,9.589212,4.0996222,5.02887,5.9542136,6.883461,7.8088045,8.738052,19.924164,31.110277,42.300293,53.48641,64.67642,54.9857,45.29497,35.604244,25.913517,16.226696,16.36335,16.500004,16.636658,16.773312,16.91387,15.660558,14.407245,13.153932,11.900618,10.651209,10.202203,9.753197,9.308095,8.859089,8.413987,7.4691215,6.5281606,5.5832953,4.6423345,3.7013733,4.2362766,4.775084,5.3138914,5.8487945,6.387602,6.5945354,6.801469,7.008402,7.2192397,7.426173,9.089449,10.756628,12.419904,14.0831785,15.750359,15.344301,14.934339,14.528281,14.118319,13.712261,13.337439,12.962616,12.587793,12.212971,11.838148,12.068507,12.298867,12.529227,12.755682,12.986042,13.095366,13.200784,13.310107,13.419431,13.524849,13.571702,13.618555,13.6693125,13.716166,13.763018,12.306676,10.84643,9.390087,7.9337454,6.473499,5.903456,5.3334136,4.7633705,4.193328,3.6232853,2.900971,2.174752,1.4485333,0.7262188,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21083772,0.42167544,0.62860876,0.8394465,1.0502841,0.8394465,0.62860876,0.42167544,0.21083772,0.0,0.0,0.0,0.0,0.0,0.0,0.14836729,0.30063897,0.44900626,0.60127795,0.74964523,1.6710842,2.5964274,3.5178664,4.4393053,5.3607445,4.6110992,3.8614538,3.1118085,2.3621633,1.6125181,1.5031948,1.397776,1.2884527,1.183034,1.0737107,3.7794614,6.4852123,9.190963,11.896713,14.59856,15.41458,16.2306,17.04662,17.858736,18.674755,16.121277,13.567798,11.018223,8.464745,5.911265,7.230953,8.554545,9.874233,11.193921,12.513609,10.639496,8.765383,6.8951745,5.0210614,3.1508527,2.8111696,2.475391,2.135708,1.7999294,1.4641509,1.6164225,1.7686942,1.9209659,2.0732377,2.2255092,2.1591344,2.096664,2.0302892,1.9639144,1.901444,1.5734742,1.2494087,0.92534333,0.60127795,0.27330816,0.21864653,0.1639849,0.10932326,0.05466163,0.0,0.46071947,0.60127795,0.7418364,0.8823949,1.0229534,1.1635119,3.1898966,5.2162814,7.2465706,9.272955,11.29934,12.829865,14.360392,15.890917,17.421442,18.95197,18.229654,17.511244,16.788929,16.07052,15.348206,17.198893,19.049578,20.900265,22.750952,24.601639,25.070168,25.538694,26.011127,26.479656,26.948185,22.11063,17.26917,12.431617,7.590158,2.7486992,2.4324427,2.1161861,1.796025,1.4797685,1.1635119,1.2650263,1.3665408,1.4680552,1.5734742,1.6749885,2.330928,2.9868677,3.638903,4.2948427,4.950782,4.2557983,3.5608149,2.8658314,2.1708477,1.475864,1.2455044,1.0151446,0.78478485,0.5544251,0.3240654,0.40605783,0.48805028,0.57394713,0.6559396,0.737932,2.1435168,3.5491016,4.950782,6.356367,7.7619514,6.2470436,4.732136,3.2172275,1.7023194,0.18741131,0.8394465,1.4914817,2.1435168,2.7994564,3.4514916,3.2094188,2.9634414,2.7213683,2.4792955,2.2372224,2.0068626,1.7765031,1.5461433,1.3157835,1.0893283,1.5734742,2.05762,2.541766,3.0259118,3.513962,3.7326086,3.951255,4.173806,4.3924527,4.6110992,5.0757227,5.5364423,6.001066,6.461786,6.9264097,7.211431,7.4964523,7.7814736,8.066495,8.351517,9.14411,9.936704,10.729298,11.521891,12.314485,11.389141,10.467703,9.546264,8.62092,7.699481,8.148487,8.59359,9.042596,9.491602,9.936704,9.343235,8.745861,8.152391,7.558923,6.9615493,5.8292727,4.6930914,3.5569105,2.4207294,1.2884527,1.7257458,2.1669433,2.6081407,3.049338,3.4866312,3.377308,3.2679846,3.1586614,3.049338,2.9361105,4.185519,5.4310236,6.6804323,7.9259367,9.175345,9.261242,9.343235,9.4291315,9.515028,9.600925,8.413987,7.230953,6.044015,4.860981,3.6740425,3.3421683,3.0102942,2.67842,2.3465457,2.0107672,1.6906061,1.3665408,1.0463798,0.7223144,0.39824903,0.42948425,0.46071947,0.48805028,0.5192855,0.5505207,0.8433509,1.1400855,1.43682,1.7296503,2.0263848,2.1669433,2.3114061,2.4519646,2.5964274,2.736986,3.677947,4.618908,5.5559645,6.4969254,7.437886,7.37932,7.320754,7.266093,7.2075267,7.1489606,5.9620223,4.775084,3.5881457,2.4012074,1.2142692,1.1986516,1.1869383,1.175225,1.1635119,1.1517987,0.92924774,0.7106012,0.48805028,0.26940376,0.05075723,0.30844778,0.5700427,0.8316377,1.0893283,1.3509232,1.3509232,1.3509232,1.3509232,1.3509232,1.3509232,1.0815194,0.80821127,0.5388075,0.26940376,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.015617609,0.015617609,0.019522011,0.023426414,0.023426414,0.06637484,0.10541886,0.14446288,0.1835069,0.22645533,1.2220778,2.2216048,3.2172275,4.2167544,5.212377,4.4275923,3.6428072,2.8580225,2.0732377,1.2884527,1.3509232,1.4133936,1.475864,1.5383345,1.6008049,1.2962615,0.9917182,0.6832704,0.37872702,0.07418364,0.12103647,0.1717937,0.21864653,0.26549935,0.31235218,0.28111696,0.24597734,0.21474212,0.1835069,0.14836729,0.15617609,0.1639849,0.1717937,0.1796025,0.18741131,0.1639849,0.14055848,0.12103647,0.09761006,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.03513962,0.046852827,0.05466163,0.06637484,0.07418364,0.19912452,0.32016098,0.44119745,0.5661383,0.6871748,0.7106012,0.7340276,0.75354964,0.77697605,0.80040246,0.6481308,0.4958591,0.3435874,0.19131571,0.039044023,0.039044023,0.042948425,0.046852827,0.046852827,0.05075723,0.7066968,1.358732,2.0146716,2.6706111,3.3265507,4.3143644,5.298274,6.2860875,7.2739015,8.261715,7.590158,6.918601,6.2431393,5.571582,4.900025,3.9200199,2.9400148,1.9600099,0.98000497,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.13665408,0.12103647,0.10932326,0.093705654,0.078088045,0.062470436,0.11713207,0.1717937,0.22645533,0.28111696,0.3357786,1.4172981,2.4988174,3.5764325,4.657952,5.7394714,8.757574,11.775677,14.797685,17.815788,20.837795,17.202797,13.571702,9.940608,6.3056097,2.6745155,3.4827268,4.290938,5.099149,5.903456,6.7116675,22.50107,38.286568,54.07597,69.86147,85.65087,71.35295,57.058933,42.76492,28.470901,14.176885,14.96167,15.750359,16.539047,17.323833,18.112522,16.640562,15.172507,13.700547,12.232492,10.764437,10.159255,9.554072,8.94889,8.343708,7.7385254,6.610153,5.481781,4.3534083,3.2289407,2.1005683,2.7643168,3.4241607,4.087909,4.7516575,5.4115014,5.8214636,6.2314262,6.6413884,7.0513506,7.461313,8.519405,9.577498,10.6355915,11.693685,12.751778,12.763491,12.779109,12.794726,12.810344,12.825961,12.373051,11.924045,11.475039,11.0260315,10.573121,11.275913,11.978706,12.681499,13.384291,14.087084,14.247164,14.407245,14.567325,14.727406,14.8874855,14.828919,14.774258,14.7156925,14.657126,14.59856,12.337912,10.081166,7.8205175,5.559869,3.2992198,3.1039999,2.9048753,2.7057507,2.5105307,2.3114061,1.8506867,1.3860629,0.92534333,0.46071947,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28111696,0.5583295,0.8394465,1.1205635,1.4016805,1.1205635,0.8394465,0.5583295,0.28111696,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,1.2064602,2.0341935,2.8658314,3.6935644,4.5252023,4.025439,3.5256753,3.0259118,2.5261483,2.0263848,1.7257458,1.4290112,1.1322767,0.8355421,0.5388075,2.1669433,3.7911747,5.4193106,7.0474463,8.675582,11.170495,13.665408,16.16032,18.655233,21.150146,18.093,15.035853,11.978706,8.921559,5.8644123,7.195813,8.531119,9.866425,11.20173,12.537036,10.58093,8.628729,6.6726236,4.716518,2.7643168,2.3855898,2.0107672,1.6359446,1.261122,0.8862993,1.0073358,1.1283722,1.2494087,1.3665408,1.4875772,1.3782539,1.2728351,1.1635119,1.0580931,0.94876975,0.78868926,0.62470436,0.46071947,0.30063897,0.13665408,0.10932326,0.08199245,0.05466163,0.027330816,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.7994564,5.5989127,8.398369,11.20173,14.001186,15.93777,17.874353,19.810938,21.751425,23.68801,22.649437,21.610867,20.5762,19.537628,18.499058,20.81437,23.125774,25.437181,27.748587,30.063898,30.223978,30.387962,30.551949,30.712029,30.876013,24.69925,18.526388,12.349625,6.1767645,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,1.33921,2.5495746,3.7638438,4.9742084,6.1884775,5.173333,4.1620927,3.1508527,2.135708,1.1244678,0.9019169,0.6754616,0.44900626,0.22645533,0.0,0.0,0.0,0.0,0.0,0.0,1.8623998,3.7247996,5.5871997,7.4495993,9.311999,7.461313,5.610626,3.7638438,1.9131571,0.062470436,0.76135844,1.4641509,2.1630387,2.8619268,3.5608149,3.4007344,3.2367494,3.076669,2.912684,2.7486992,2.3114061,1.8741131,1.43682,0.999527,0.5622339,0.8238289,1.0893283,1.3509232,1.6125181,1.8741131,2.0107672,2.1513257,2.2879796,2.4246337,2.5612879,3.5608149,4.564246,5.563773,6.5633,7.562827,7.9376497,8.312472,8.687295,9.062118,9.43694,10.436467,11.435994,12.439425,13.438952,14.438479,13.16174,11.888905,10.612165,9.339331,8.062591,8.761478,9.464272,10.163159,10.862047,11.560935,10.81129,10.061645,9.311999,8.562354,7.812709,6.4383593,5.0640097,3.6857557,2.3114061,0.93705654,1.1127546,1.2884527,1.4641509,1.6359446,1.8116426,1.7491722,1.6867018,1.6242313,1.5617609,1.4992905,3.1235218,4.7516575,6.375889,8.00012,9.6243515,9.964035,10.299813,10.6355915,10.975275,11.311053,9.948417,8.58578,7.223144,5.8644123,4.5017757,4.0996222,3.7013733,3.2992198,2.900971,2.4988174,2.1005683,1.698415,1.3001659,0.9019169,0.4997635,0.5231899,0.5505207,0.57394713,0.60127795,0.62470436,0.8238289,1.0268579,1.2259823,1.4251068,1.6242313,1.7608855,1.901444,2.0380979,2.174752,2.3114061,2.9361105,3.5608149,4.1894236,4.814128,5.4388323,5.8644123,6.2860875,6.7116675,7.137247,7.562827,6.3251314,5.087436,3.8497405,2.612045,1.3743496,1.3235924,1.2767396,1.2259823,1.175225,1.1244678,0.9136301,0.698888,0.48805028,0.27330816,0.062470436,0.30063897,0.5388075,0.77307165,1.0112402,1.2494087,1.33921,1.4251068,1.5110037,1.6008049,1.6867018,1.3509232,1.0112402,0.6754616,0.3357786,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,1.4133936,2.639376,3.8614538,5.087436,6.3134184,5.22409,4.138666,3.049338,1.9639144,0.8745861,0.92534333,0.97610056,1.0268579,1.0737107,1.1244678,0.9019169,0.6754616,0.44900626,0.22645533,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.1639849,0.26159495,0.3631094,0.46071947,0.5622339,0.5114767,0.46071947,0.41386664,0.3631094,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6754616,1.3509232,2.0263848,2.7018464,3.3734035,3.5998588,3.8263142,4.0488653,4.2753205,4.5017757,3.5998588,2.7018464,1.7999294,0.9019169,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,1.4992905,2.87364,4.251894,5.6262436,7.000593,7.6252975,8.250002,8.874706,9.499411,10.124115,8.351517,6.575013,4.7985106,3.0259118,1.2494087,1.9365835,2.6237583,3.310933,3.998108,4.689187,25.077976,45.46286,65.85165,86.236534,106.62532,87.72411,68.826805,49.92559,31.02438,12.123169,13.563893,15.000713,16.437534,17.874353,19.311174,17.624472,15.93777,14.251068,12.564366,10.87376,10.112402,9.351044,8.58578,7.824422,7.0630636,5.7511845,4.4393053,3.1235218,1.8116426,0.4997635,1.2884527,2.0732377,2.8619268,3.6506162,4.4393053,5.0483923,5.661383,6.2743745,6.8873653,7.5003567,7.9493628,8.398369,8.85128,9.300286,9.749292,10.186585,10.6238785,11.061172,11.498465,11.935758,11.412568,10.889378,10.362284,9.839094,9.311999,10.487225,11.66245,12.837675,14.012899,15.188125,15.398962,15.613705,15.824542,16.039284,16.250122,16.086138,15.926057,15.762072,15.598087,15.438006,12.373051,9.311999,6.250948,3.1859922,0.12494087,0.30063897,0.47633708,0.6481308,0.8238289,0.999527,0.80040246,0.60127795,0.39824903,0.19912452,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3513962,0.698888,1.0502841,1.4016805,1.7491722,1.4016805,1.0502841,0.698888,0.3513962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.737932,1.475864,2.2137961,2.951728,3.6857557,3.435874,3.1859922,2.9361105,2.6862288,2.436347,1.9482968,1.4641509,0.97610056,0.48805028,0.0,0.5505207,1.1010414,1.6515622,2.1981785,2.7486992,6.9264097,11.100216,15.274021,19.447828,23.625538,20.06082,16.500004,12.939189,9.37447,5.813655,7.1606736,8.511597,9.86252,11.213444,12.564366,10.526268,8.488171,6.4500723,4.4119744,2.3738766,1.9639144,1.5500476,1.1361811,0.7262188,0.31235218,0.39824903,0.48805028,0.57394713,0.6637484,0.74964523,0.60127795,0.44900626,0.30063897,0.14836729,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.260649,4.5252023,6.785851,9.050405,11.311053,14.215929,17.1169,20.021774,22.922745,25.823717,23.851994,21.88027,19.908546,17.936825,15.961197,17.581524,19.197947,20.81437,22.430792,24.051117,24.179964,24.30881,24.441559,24.570404,24.69925,19.908546,15.113941,10.323239,5.5286336,0.737932,0.98000497,1.2220778,1.4641509,1.7062237,1.9482968,2.0029583,2.0537157,2.1083772,2.1591344,2.2137961,2.8463092,3.4827268,4.1191444,4.7516575,5.388075,4.493967,3.6037633,2.7096553,1.815547,0.92534333,0.76135844,0.60127795,0.43729305,0.27330816,0.113227665,0.10932326,0.10151446,0.09761006,0.093705654,0.08589685,1.9209659,3.7521305,5.5832953,7.4183645,9.249529,7.47693,5.700427,3.9239242,2.1513257,0.37482262,1.0073358,1.639849,2.2723622,2.9048753,3.5373883,3.5608149,3.5881457,3.611572,3.638903,3.6623292,3.213323,2.7643168,2.3114061,1.8623998,1.4133936,1.5656652,1.717937,1.8702087,2.0224805,2.174752,2.3465457,2.5183394,2.6940374,2.8658314,3.0376248,3.8419318,4.6423345,5.446641,6.2470436,7.0513506,7.504261,7.9610763,8.413987,8.870802,9.323712,9.940608,10.553599,11.170495,11.783486,12.400381,11.342289,10.284196,9.226103,8.16801,7.113821,7.832231,8.550641,9.272955,9.991365,10.71368,9.917182,9.120684,8.32809,7.531592,6.7389984,5.591104,4.4432096,3.2953155,2.1474214,0.999527,1.1908426,1.3782539,1.5695697,1.7608855,1.9482968,1.8663043,1.7804074,1.6945106,1.6086137,1.5266213,2.9087796,4.2948427,5.6809053,7.0630636,8.449126,8.870802,9.288573,9.710248,10.131924,10.549695,9.351044,8.156297,6.957645,5.758993,4.564246,4.1035266,3.6467118,3.1898966,2.7330816,2.2762666,1.9522011,1.6281357,1.3079748,0.98390937,0.6637484,0.6949836,0.7262188,0.76135844,0.79259366,0.8238289,1.0112402,1.1947471,1.3782539,1.5656652,1.7491722,1.8116426,1.8702087,1.9287747,1.9912452,2.0498111,2.6159496,3.1781836,3.7443218,4.31046,4.8765984,5.4271193,5.9815445,6.532065,7.08649,7.6370106,6.5633,5.493494,4.4197836,3.3460727,2.2762666,2.1083772,1.9443923,1.7804074,1.6164225,1.4485333,1.2689307,1.0854238,0.9019169,0.71841,0.5388075,0.6637484,0.79259366,0.92143893,1.0463798,1.175225,1.3235924,1.475864,1.6242313,1.7765031,1.9248703,1.5969005,1.2689307,0.94096094,0.61689556,0.28892577,0.23035973,0.1717937,0.113227665,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.21083772,0.42557985,0.63641757,0.8511597,1.0619974,2.1435168,3.2211318,4.3026514,5.3841705,6.461786,5.3334136,4.2089458,3.0805733,1.9522011,0.8238289,0.8433509,0.8667773,0.8862993,0.9058213,0.92534333,0.7418364,0.5583295,0.37872702,0.19522011,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.06637484,0.12884527,0.19522011,0.26159495,0.3240654,0.3240654,0.32016098,0.31625658,0.31625658,0.31235218,0.26940376,0.22645533,0.1835069,0.14055848,0.10151446,0.14055848,0.1796025,0.21864653,0.26159495,0.30063897,0.26159495,0.22645533,0.18741131,0.14836729,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.14446288,0.23816854,0.3357786,0.42948425,0.5231899,0.48414588,0.44119745,0.39824903,0.3553006,0.31235218,0.25378615,0.19912452,0.14055848,0.08199245,0.023426414,0.38653582,0.74574083,1.1049459,1.4641509,1.8233559,1.4602464,1.0932326,0.7301232,0.3631094,0.0,0.5505207,1.1010414,1.6515622,2.1981785,2.7486992,2.9243972,3.096191,3.2679846,3.4397783,3.611572,3.2016098,2.787743,2.3738766,1.9639144,1.5500476,1.3509232,1.1517987,0.94876975,0.74964523,0.5505207,0.47633708,0.39824903,0.3240654,0.24988174,0.1756981,0.14836729,0.12494087,0.10151446,0.07418364,0.05075723,0.08589685,0.12103647,0.15617609,0.19131571,0.22645533,1.3001659,2.3738766,3.4514916,4.5252023,5.5989127,6.434455,7.266093,8.097731,8.929368,9.761005,8.98403,8.203149,7.422269,6.6413884,5.8644123,6.4422636,7.0240197,7.601871,8.183627,8.761478,24.69925,40.633114,56.56698,72.50085,88.438614,73.80492,59.171215,44.537518,29.90772,15.274021,16.874826,18.475632,20.076437,21.673336,23.274141,21.118912,18.959778,16.800642,14.645412,12.486279,11.631214,10.77615,9.921086,9.066022,8.210958,6.7897553,5.368553,3.9434462,2.522244,1.1010414,1.7843118,2.463678,3.1469483,3.8302186,4.513489,5.040583,5.571582,6.1025805,6.6335793,7.1606736,7.3324676,7.504261,7.6721506,7.843944,8.011833,8.531119,9.0465,9.565785,10.081166,10.600452,10.194394,9.788337,9.386183,8.980125,8.574067,9.811763,11.0494585,12.287154,13.524849,14.762545,14.606369,14.454097,14.297921,14.141745,13.985569,13.661504,13.337439,13.013372,12.689307,12.361338,9.909373,7.4574084,5.0054436,2.5534792,0.10151446,0.23816854,0.37872702,0.5192855,0.659844,0.80040246,0.64032197,0.48024148,0.32016098,0.16008049,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28111696,0.5583295,0.8394465,1.1205635,1.4016805,1.1205635,0.8394465,0.5583295,0.28111696,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.58956474,1.1791295,1.7686942,2.358259,2.951728,2.7565079,2.5612879,2.366068,2.1708477,1.9756275,1.5812829,1.183034,0.78868926,0.39434463,0.0,0.59346914,1.1908426,1.7843118,2.3816853,2.9751544,6.2158084,9.456462,12.693212,15.933866,19.174519,16.515621,13.860628,11.20173,8.546737,5.8878384,6.8678436,7.8478484,8.827853,9.807858,10.787864,9.921086,9.058213,8.191436,7.328563,6.461786,5.852699,5.2436123,4.630621,4.0215344,3.4124475,2.8892577,2.366068,1.8467822,1.3235924,0.80040246,0.71841,0.64032197,0.5583295,0.48024148,0.39824903,0.32016098,0.23816854,0.16008049,0.078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.7257458,3.4514916,5.173333,6.899079,8.624825,12.494087,16.359446,20.228708,24.094067,27.96333,25.05455,22.14577,19.240894,16.332115,13.423335,14.348679,15.270117,16.191557,17.1169,18.038338,18.135948,18.233559,18.33117,18.42878,18.526388,15.113941,11.705398,8.292951,4.884407,1.475864,1.9365835,2.3933985,2.854118,3.3148375,3.775557,3.8809757,3.9863946,4.0918136,4.193328,4.298747,4.357313,4.415879,4.474445,4.5291066,4.5876727,3.814601,3.0415294,2.2684577,1.4992905,0.7262188,0.62470436,0.5231899,0.42557985,0.3240654,0.22645533,0.21474212,0.20693332,0.19522011,0.1835069,0.1756981,1.9756275,3.7794614,5.5832953,7.3832245,9.187058,7.4886436,5.786324,4.087909,2.3855898,0.6871748,1.2533131,1.815547,2.3816853,2.9478238,3.513962,3.7247996,3.9356375,4.1503797,4.3612175,4.575959,4.1113358,3.6506162,3.1859922,2.7252727,2.260649,2.3035975,2.3465457,2.3894942,2.4324427,2.475391,2.6823244,2.8892577,3.096191,3.3031244,3.513962,4.1191444,4.7243266,5.3256044,5.930787,6.5359693,7.0708723,7.605776,8.140678,8.675582,9.21439,9.440845,9.671205,9.901564,10.131924,10.362284,9.522837,8.683391,7.843944,7.000593,6.1611466,6.902983,7.6409154,8.382751,9.120684,9.86252,9.023073,8.183627,7.3441806,6.5008297,5.661383,4.743849,3.8224099,2.900971,1.9834363,1.0619974,1.2689307,1.4719596,1.678893,1.8819219,2.0888553,1.979532,1.8741131,1.7647898,1.6593709,1.5500476,2.6940374,3.8380275,4.985922,6.1299114,7.2739015,7.7775693,8.281238,8.781001,9.284669,9.788337,8.75367,7.7229075,6.688241,5.657479,4.6267166,4.1113358,3.5959544,3.0805733,2.5651922,2.0498111,1.8038338,1.5617609,1.3157835,1.0698062,0.8238289,0.8667773,0.9058213,0.94486535,0.98390937,1.0268579,1.1947471,1.3665408,1.53443,1.7062237,1.8741131,1.8584955,1.8389735,1.8233559,1.8038338,1.7882162,2.2918842,2.795552,3.3031244,3.8067923,4.3143644,4.9937305,5.6730967,6.3524623,7.0318284,7.7111945,6.805373,5.8956475,4.989826,4.084005,3.174279,2.893162,2.6159496,2.3348327,2.0537157,1.7765031,1.6242313,1.4719596,1.3157835,1.1635119,1.0112402,1.0307622,1.0463798,1.0659018,1.0815194,1.1010414,1.3118792,1.5266213,1.737459,1.9482968,2.1630387,1.8467822,1.5266213,1.2103647,0.8941081,0.57394713,0.46071947,0.3435874,0.23035973,0.113227665,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.38653582,0.77307165,1.1635119,1.5500476,1.9365835,2.87364,3.8067923,4.743849,5.677001,6.6140575,5.446641,4.279225,3.1118085,1.9443923,0.77307165,0.76526284,0.75354964,0.74574083,0.7340276,0.7262188,0.58566034,0.44510186,0.30454338,0.1639849,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.10541886,0.21083772,0.31625658,0.42167544,0.5231899,0.5309987,0.5388075,0.5466163,0.5544251,0.5622339,0.47633708,0.39434463,0.30844778,0.22255093,0.13665408,0.23035973,0.3240654,0.41386664,0.5075723,0.60127795,0.5231899,0.44900626,0.37482262,0.30063897,0.22645533,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.12884527,0.21864653,0.30844778,0.39824903,0.48805028,0.45291066,0.41777104,0.38263142,0.3474918,0.31235218,0.26159495,0.20693332,0.15617609,0.10151446,0.05075723,0.76916724,1.4914817,2.2098918,2.9283018,3.6506162,2.920493,2.1903696,1.4602464,0.7301232,0.0,0.42557985,0.8511597,1.2767396,1.698415,2.1239948,2.2450314,2.366068,2.4831998,2.6042364,2.7252727,2.7994564,2.87364,2.951728,3.0259118,3.1000953,2.7018464,2.2996929,1.901444,1.4992905,1.1010414,0.94876975,0.80040246,0.6481308,0.4997635,0.3513962,0.28892577,0.22645533,0.1639849,0.10151446,0.039044023,0.093705654,0.15227169,0.21083772,0.26940376,0.3240654,1.1010414,1.8741131,2.6510892,3.4241607,4.2011366,5.239708,6.278279,7.320754,8.359325,9.4018,9.616543,9.8312845,10.046027,10.260769,10.475512,10.947944,11.420377,11.892809,12.365242,12.837675,24.320522,35.803368,47.286217,58.769062,70.24801,59.885723,49.519535,39.153347,28.791061,18.424873,20.18576,21.95055,23.711435,25.476225,27.23711,24.609447,21.981785,19.354122,16.72646,14.098797,13.153932,12.205161,11.256392,10.311526,9.362757,7.8283267,6.297801,4.7633705,3.232845,1.698415,2.2762666,2.854118,3.4319696,4.009821,4.5876727,5.036679,5.481781,5.930787,6.375889,6.824895,6.715572,6.606249,6.4969254,6.3836975,6.2743745,6.871748,7.4691215,8.066495,8.663869,9.261242,8.976221,8.691199,8.406178,8.121157,7.8361354,9.136301,10.436467,11.736633,13.036799,14.336966,13.813775,13.2905855,12.771299,12.24811,11.72492,11.23687,10.748819,10.260769,9.776623,9.288573,7.445695,5.602817,3.7599394,1.9170616,0.07418364,0.1796025,0.28502136,0.39044023,0.4958591,0.60127795,0.48024148,0.359205,0.23816854,0.12103647,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21083772,0.42167544,0.62860876,0.8394465,1.0502841,0.8394465,0.62860876,0.42167544,0.21083772,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.44119745,0.8862993,1.3274968,1.7686942,2.2137961,2.0732377,1.9326792,1.7921207,1.6515622,1.5110037,1.2103647,0.9058213,0.60518235,0.30063897,0.0,0.64032197,1.2806439,1.9209659,2.5612879,3.2016098,5.505207,7.8088045,10.116306,12.419904,14.723501,12.970425,11.221252,9.468176,7.715099,5.9620223,6.571109,7.1841,7.793187,8.402273,9.01136,9.319808,9.628256,9.936704,10.241247,10.549695,9.741484,8.933272,8.128965,7.320754,6.5125427,5.380266,4.2479897,3.1157131,1.9834363,0.8511597,0.8394465,0.8316377,0.8199245,0.80821127,0.80040246,0.64032197,0.48024148,0.32016098,0.16008049,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1869383,2.3738766,3.5608149,4.7516575,5.938596,10.768341,15.601992,20.435642,25.26929,30.099037,26.257105,22.415173,18.573242,14.73131,10.889378,11.115833,11.342289,11.568744,11.799104,12.025558,12.091934,12.154405,12.220779,12.28325,12.349625,10.323239,8.296855,6.266566,4.240181,2.2137961,2.8892577,3.5686235,4.2440853,4.9234514,5.5989127,5.758993,5.9151692,6.0713453,6.2314262,6.387602,5.8683167,5.349031,4.825841,4.3065557,3.78727,3.135235,2.4831998,1.8311646,1.1791295,0.5231899,0.48805028,0.44900626,0.41386664,0.37482262,0.3357786,0.3240654,0.30844778,0.29283017,0.27721256,0.26159495,2.0341935,3.8067923,5.579391,7.3519893,9.124588,7.5003567,5.8761253,4.251894,2.6237583,0.999527,1.4992905,1.9951496,2.4910088,2.9907722,3.4866312,3.8887846,4.2870336,4.689187,5.087436,5.4856853,5.0132523,4.5369153,4.0605783,3.5881457,3.1118085,3.0454338,2.979059,2.9087796,2.8424048,2.77603,3.018103,3.260176,3.5022488,3.7443218,3.9863946,4.396357,4.802415,5.2084727,5.618435,6.0244927,6.6413884,7.2543793,7.871275,8.484266,9.101162,8.944985,8.78881,8.636538,8.480362,8.324185,7.703386,7.0786815,6.4578815,5.833177,5.212377,5.9737353,6.7311897,7.492548,8.253906,9.01136,8.128965,7.2426662,6.356367,5.473972,4.5876727,3.8965936,3.2016098,2.5105307,1.815547,1.1244678,1.3431144,1.5656652,1.7843118,2.0068626,2.2255092,2.096664,1.9639144,1.8350691,1.7062237,1.5734742,2.4792955,3.3851168,4.290938,5.196759,6.098676,6.6843367,7.269997,7.8556576,8.441318,9.023073,8.156297,7.289519,6.422742,5.5559645,4.689187,4.11524,3.541293,2.97125,2.397303,1.8233559,1.6593709,1.4914817,1.3235924,1.1557031,0.9878138,1.0346665,1.0815194,1.1283722,1.1791295,1.2259823,1.3782539,1.53443,1.6906061,1.8467822,1.999054,1.9053483,1.8116426,1.7140326,1.620327,1.5266213,1.9717231,2.416825,2.8619268,3.3031244,3.7482262,4.5564375,5.364649,6.17286,6.9810715,7.7892823,7.043542,6.3017054,5.559869,4.8180323,4.0761957,3.6818514,3.2836022,2.8892577,2.494913,2.1005683,1.9756275,1.8545911,1.7335546,1.6086137,1.4875772,1.3938715,1.3040704,1.2103647,1.116659,1.0268579,1.3001659,1.5734742,1.8506867,2.1239948,2.4012074,2.0927596,1.7843118,1.475864,1.1713207,0.8628729,0.6910792,0.5192855,0.3435874,0.1717937,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.5622339,1.1244678,1.6867018,2.2489357,2.8111696,3.6037633,4.3924527,5.181142,5.9737353,6.7624245,5.5559645,4.3455997,3.1391394,1.9326792,0.7262188,0.6832704,0.6442264,0.60518235,0.5661383,0.5231899,0.42557985,0.3318742,0.23426414,0.13665408,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.14446288,0.28892577,0.43338865,0.58175594,0.7262188,0.7418364,0.76135844,0.77697605,0.79649806,0.81211567,0.6832704,0.5583295,0.42948425,0.30063897,0.1756981,0.32016098,0.46462387,0.60908675,0.75354964,0.9019169,0.78868926,0.6754616,0.5622339,0.44900626,0.3357786,0.27330816,0.21083772,0.14836729,0.08589685,0.023426414,0.10932326,0.19522011,0.28111696,0.3631094,0.44900626,0.42167544,0.39434463,0.3670138,0.339683,0.31235218,0.26549935,0.21864653,0.1717937,0.12103647,0.07418364,1.1557031,2.233318,3.3148375,4.396357,5.473972,4.380739,3.2836022,2.1903696,1.0932326,0.0,0.30063897,0.60127795,0.9019169,1.1986516,1.4992905,1.5656652,1.6359446,1.7023194,1.7686942,1.8389735,2.4012074,2.9634414,3.5256753,4.087909,4.650143,4.0488653,3.4514916,2.8502135,2.2489357,1.6515622,1.4251068,1.1986516,0.97610056,0.74964523,0.5231899,0.42557985,0.3240654,0.22645533,0.12494087,0.023426414,0.10541886,0.1835069,0.26549935,0.3435874,0.42557985,0.9019169,1.3743496,1.8506867,2.3231194,2.7994564,4.0488653,5.2943697,6.5437784,7.7892823,9.0386915,10.249056,11.455516,12.665881,13.8762455,15.086611,15.453624,15.816733,16.183748,16.546856,16.91387,23.941795,30.973623,38.00155,45.033375,52.0613,45.966526,39.86785,33.769176,27.670498,21.575727,23.500597,25.425468,27.350338,29.275208,31.200079,28.103888,25.003792,21.9076,18.81141,15.711315,14.672744,13.634172,12.591698,11.553126,10.510651,8.870802,7.2270484,5.5832953,3.9434462,2.2996929,2.7721257,3.2445583,3.716991,4.1894236,4.661856,5.02887,5.3919797,5.758993,6.1221027,6.4891167,6.098676,5.708236,5.3177958,4.927356,4.5369153,5.2162814,5.891743,6.571109,7.2465706,7.9259367,7.7619514,7.5940623,7.4300776,7.266093,7.098203,8.460839,9.823476,11.186112,12.548749,13.911386,13.021181,12.130978,11.240774,10.350571,9.464272,8.812236,8.164105,7.5120697,6.8639393,6.211904,4.9781127,3.7482262,2.514435,1.2806439,0.05075723,0.12103647,0.19131571,0.26159495,0.3318742,0.39824903,0.32016098,0.23816854,0.16008049,0.078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14055848,0.28111696,0.42167544,0.5583295,0.698888,0.5583295,0.42167544,0.28111696,0.14055848,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29673457,0.58956474,0.8862993,1.1791295,1.475864,1.3899672,1.3040704,1.2181735,1.1361811,1.0502841,0.8394465,0.62860876,0.42167544,0.21083772,0.0,0.6832704,1.3704453,2.0537157,2.7408905,3.4241607,4.794606,6.165051,7.535496,8.905942,10.276386,9.4291315,8.577971,7.7307167,6.883461,6.036206,6.278279,6.5164475,6.75852,6.996689,7.238762,8.718531,10.198298,11.678067,13.157836,14.637604,13.634172,12.626837,11.623405,10.61607,9.612638,7.871275,6.126007,4.3846436,2.6432803,0.9019169,0.96048295,1.0190489,1.0815194,1.1400855,1.1986516,0.96048295,0.71841,0.48024148,0.23816854,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6481308,1.3001659,1.9482968,2.6003318,3.2484627,9.0465,14.844538,20.642574,26.440613,32.23865,27.459661,22.684578,17.905588,13.1266,8.351517,7.882988,7.4144597,6.9459314,6.481308,6.012779,6.044015,6.0791545,6.1103897,6.141625,6.1767645,5.5286336,4.884407,4.240181,3.5959544,2.951728,3.8458362,4.7399445,5.6340523,6.5281606,7.426173,7.633106,7.843944,8.054782,8.265619,8.476458,7.37932,6.278279,5.181142,4.084005,2.9868677,2.455869,1.9209659,1.3899672,0.8589685,0.3240654,0.3513962,0.37482262,0.39824903,0.42557985,0.44900626,0.42948425,0.40996224,0.39044023,0.3709182,0.3513962,2.0927596,3.8341231,5.579391,7.320754,9.062118,7.5120697,5.9620223,4.4119744,2.8619268,1.3118792,1.7413634,2.1708477,2.6042364,3.0337205,3.4632049,4.0488653,4.6384296,5.22409,5.813655,6.3993154,5.911265,5.423215,4.939069,4.4510183,3.9629683,3.7833657,3.6076677,3.4280653,3.252367,3.076669,3.3538816,3.631094,3.9083066,4.185519,4.462732,4.6735697,4.884407,5.0913405,5.3021784,5.5130157,6.2079997,6.902983,7.5979667,8.292951,8.987934,8.449126,7.9064145,7.367607,6.8287997,6.2860875,5.883934,5.477876,5.0718184,4.6657605,4.263607,5.040583,5.8214636,6.602344,7.3832245,8.164105,7.230953,6.3017054,5.3724575,4.4432096,3.513962,3.049338,2.5808098,2.1161861,1.6515622,1.1869383,1.4212024,1.6593709,1.893635,2.1278992,2.3621633,2.2098918,2.05762,1.9053483,1.7530766,1.6008049,2.2645533,2.9283018,3.5959544,4.2597027,4.9234514,5.591104,6.2587566,6.9264097,7.5940623,8.261715,7.558923,6.8561306,6.153338,5.4505453,4.7516575,4.1191444,3.4905357,2.8619268,2.2294137,1.6008049,1.5110037,1.4212024,1.3314011,1.2415999,1.1517987,1.2064602,1.261122,1.3157835,1.3704453,1.4251068,1.5656652,1.7062237,1.8467822,1.9834363,2.1239948,1.9522011,1.7804074,1.6086137,1.43682,1.261122,1.6476578,2.0341935,2.416825,2.803361,3.1859922,4.123049,5.056201,5.9932575,6.9264097,7.8634663,7.2856145,6.707763,6.1299114,5.55206,4.9742084,4.466636,3.9551594,3.4436827,2.9361105,2.4246337,2.330928,2.241127,2.1474214,2.0537157,1.9639144,1.7608855,1.5578566,1.3548276,1.1517987,0.94876975,1.2884527,1.6242313,1.9639144,2.2996929,2.639376,2.338737,2.0420024,1.7452679,1.4485333,1.1517987,0.92143893,0.6910792,0.46071947,0.23035973,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.737932,1.475864,2.2137961,2.951728,3.6857557,4.3338866,4.9781127,5.6223392,6.266566,6.910792,5.6652875,4.415879,3.1703746,1.9209659,0.6754616,0.60518235,0.5349031,0.46462387,0.39434463,0.3240654,0.26940376,0.21474212,0.16008049,0.10541886,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.1835069,0.3709182,0.5544251,0.7418364,0.92534333,0.95267415,0.98000497,1.0073358,1.0346665,1.0619974,0.8941081,0.7223144,0.5544251,0.38263142,0.21083772,0.40996224,0.60908675,0.80430686,1.0034313,1.1986516,1.0502841,0.9019169,0.74964523,0.60127795,0.44900626,0.3631094,0.27330816,0.18741131,0.10151446,0.011713207,0.093705654,0.1717937,0.25378615,0.3318742,0.41386664,0.39434463,0.3709182,0.3513962,0.3318742,0.31235218,0.26940376,0.22645533,0.1835069,0.14055848,0.10151446,1.5383345,2.979059,4.4197836,5.860508,7.3012323,5.840986,4.380739,2.920493,1.4602464,0.0,0.1756981,0.3513962,0.5231899,0.698888,0.8745861,0.8902037,0.9058213,0.92143893,0.93315214,0.94876975,1.999054,3.049338,4.0996222,5.1499066,6.2001905,5.3997884,4.5993857,3.7989833,2.998581,2.1981785,1.901444,1.6008049,1.3001659,0.999527,0.698888,0.5622339,0.42557985,0.28892577,0.14836729,0.011713207,0.113227665,0.21864653,0.32016098,0.42167544,0.5231899,0.698888,0.8745861,1.0502841,1.2259823,1.4016805,2.854118,4.31046,5.7668023,7.2192397,8.675582,10.881569,13.083652,15.289639,17.495626,19.701614,19.959305,20.216995,20.470781,20.728472,20.986162,23.566973,26.143877,28.720783,31.297688,33.874596,32.04343,30.21617,28.385004,26.55384,24.72658,26.811531,28.900385,30.98924,33.074192,35.163048,31.594423,28.025799,24.46108,20.892456,17.323833,16.191557,15.059279,13.927003,12.794726,11.66245,9.909373,8.156297,6.4032197,4.6540475,2.900971,3.2679846,3.6349986,4.0020123,4.369026,4.73604,5.0210614,5.3021784,5.5832953,5.8683167,6.1494336,5.481781,4.8102236,4.138666,3.4710135,2.7994564,3.5569105,4.3143644,5.0718184,5.8292727,6.5867267,6.5437784,6.4969254,6.453977,6.407124,6.364176,7.7892823,9.21439,10.6355915,12.0606985,13.4858055,12.228588,10.971371,9.714153,8.456935,7.1997175,6.387602,5.575486,4.7633705,3.951255,3.1391394,2.514435,1.893635,1.2689307,0.6481308,0.023426414,0.058566034,0.093705654,0.12884527,0.1639849,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07027924,0.14055848,0.21083772,0.28111696,0.3513962,0.28111696,0.21083772,0.14055848,0.07027924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14836729,0.29673457,0.44119745,0.58956474,0.737932,0.7066968,0.679366,0.6481308,0.61689556,0.58566034,0.46852827,0.3513962,0.23426414,0.11713207,0.0,0.7301232,1.4602464,2.1903696,2.920493,3.6506162,4.084005,4.521298,4.9546866,5.388075,5.825368,5.883934,5.938596,5.997162,6.055728,6.114294,5.9815445,5.852699,5.7238536,5.591104,5.462259,8.113348,10.768341,13.419431,16.07052,18.725513,17.522957,16.320402,15.117846,13.91529,12.712734,10.358379,8.007929,5.6535745,3.3031244,0.94876975,1.0815194,1.2103647,1.33921,1.4680552,1.6008049,1.2806439,0.96048295,0.64032197,0.32016098,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.113227665,0.22645533,0.3357786,0.44900626,0.5622339,7.3246584,14.087084,20.849508,27.611933,34.37436,28.662216,22.950077,17.237936,11.525795,5.813655,4.650143,3.4866312,2.3231194,1.1635119,0.0,0.0,0.0,0.0,0.0,0.0,0.737932,1.475864,2.2137961,2.951728,3.6857557,4.7985106,5.911265,7.0240197,8.136774,9.249529,9.511124,9.776623,10.0382185,10.299813,10.561408,8.886419,7.211431,5.5364423,3.8614538,2.1864653,1.7765031,1.3626363,0.94876975,0.5388075,0.12494087,0.21083772,0.30063897,0.38653582,0.47633708,0.5622339,0.5388075,0.5114767,0.48805028,0.46071947,0.43729305,2.1513257,3.8614538,5.575486,7.2856145,8.999647,7.523783,6.0518236,4.575959,3.1000953,1.6242313,1.9873407,2.35045,2.7135596,3.076669,3.435874,4.21285,4.985922,5.7628975,6.5359693,7.3129454,6.813182,6.3134184,5.813655,5.3138914,4.814128,4.5252023,4.2362766,3.951255,3.6623292,3.3734035,3.6857557,3.998108,4.3143644,4.6267166,4.939069,4.950782,4.9624953,4.9742084,4.985922,5.001539,5.774611,6.551587,7.3246584,8.101635,8.874706,7.9493628,7.0240197,6.098676,5.173333,4.251894,4.0605783,3.873167,3.6857557,3.4983444,3.310933,4.1113358,4.911738,5.7121406,6.5125427,7.3129454,6.336845,5.3607445,4.388548,3.4124475,2.436347,2.1981785,1.9639144,1.7257458,1.4875772,1.2494087,1.4992905,1.7491722,1.999054,2.2489357,2.4988174,2.3231194,2.1513257,1.9756275,1.7999294,1.6242313,2.0498111,2.475391,2.900971,3.3265507,3.7482262,4.5017757,5.251421,6.001066,6.7507114,7.5003567,6.9615493,6.426646,5.8878384,5.349031,4.814128,4.126953,3.435874,2.7486992,2.0615244,1.3743496,1.3626363,1.3509232,1.33921,1.3235924,1.3118792,1.3743496,1.43682,1.4992905,1.5617609,1.6242313,1.7491722,1.8741131,1.999054,2.1239948,2.2489357,1.999054,1.7491722,1.4992905,1.2494087,0.999527,1.3235924,1.6515622,1.9756275,2.2996929,2.6237583,3.6857557,4.7516575,5.813655,6.8756523,7.9376497,7.523783,7.113821,6.699954,6.2860875,5.8761253,5.251421,4.6267166,3.998108,3.3734035,2.7486992,2.6862288,2.6237583,2.5612879,2.4988174,2.436347,2.1239948,1.8116426,1.4992905,1.1869383,0.8745861,1.2767396,1.6749885,2.0732377,2.475391,2.87364,2.5886188,2.2996929,2.0107672,1.7257458,1.43682,1.1517987,0.8628729,0.57394713,0.28892577,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.9136301,1.8233559,2.736986,3.6506162,4.564246,5.0640097,5.563773,6.0635366,6.5633,7.0630636,5.774611,4.4861584,3.2016098,1.9131571,0.62470436,0.5231899,0.42557985,0.3240654,0.22645533,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.22645533,0.44900626,0.6754616,0.9019169,1.1244678,1.1635119,1.1986516,1.2376955,1.2767396,1.3118792,1.1010414,0.8862993,0.6754616,0.46071947,0.24988174,0.4997635,0.74964523,0.999527,1.2494087,1.4992905,1.3118792,1.1244678,0.93705654,0.74964523,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.3631094,0.3513962,0.3357786,0.3240654,0.31235218,0.27330816,0.23816854,0.19912452,0.1639849,0.12494087,1.9248703,3.7247996,5.5247293,7.3246584,9.124588,7.3012323,5.473972,3.6506162,1.8233559,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,1.6008049,3.1391394,4.6735697,6.211904,7.7502384,6.7507114,5.7511845,4.7516575,3.7482262,2.7486992,2.3738766,1.999054,1.6242313,1.2494087,0.8745861,0.698888,0.5231899,0.3513962,0.1756981,0.0,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.0,1.6632754,3.3265507,4.985922,6.649197,8.312472,11.514082,14.711788,17.913397,21.111103,24.312714,24.46108,24.613352,24.761719,24.91399,25.062359,23.188246,21.314133,19.436115,17.562002,15.687888,18.124235,20.560583,23.000834,25.437181,27.873528,30.126368,32.375305,34.62424,36.873177,39.126015,35.088863,31.051712,27.010654,22.973503,18.936352,17.714273,16.48829,15.262308,14.036326,12.814248,10.947944,9.089449,7.223144,5.3607445,3.4983444,3.7638438,4.025439,4.2870336,4.548629,4.814128,5.0132523,5.212377,5.4115014,5.610626,5.813655,4.860981,3.912211,2.9634414,2.0107672,1.0619974,1.901444,2.736986,3.5764325,4.4119744,5.251421,5.3256044,5.3997884,5.473972,5.548156,5.6262436,7.113821,8.601398,10.088976,11.576552,13.06413,11.435994,9.811763,8.187531,6.5633,4.939069,3.9629683,2.9868677,2.0107672,1.038571,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.77697605,1.5500476,2.3231194,3.1000953,3.873167,3.3734035,2.87364,2.3738766,1.8741131,1.3743496,2.338737,3.2992198,4.263607,5.22409,6.1884775,5.688714,5.1889505,4.689187,4.1894236,3.6857557,7.5120697,11.338385,15.160794,18.987108,22.813423,21.411741,20.013966,18.612286,17.21451,15.812829,12.849388,9.885946,6.9264097,3.9629683,0.999527,1.1986516,1.4016805,1.6008049,1.7999294,1.999054,1.6008049,1.1986516,0.80040246,0.39824903,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14446288,0.28892577,0.43338865,0.58175594,0.7262188,6.2353306,11.744442,17.253553,22.76657,28.27568,23.570877,18.869976,14.169076,9.464272,4.7633705,3.8224099,2.8814487,1.9443923,1.0034313,0.062470436,0.05466163,0.046852827,0.039044023,0.031235218,0.023426414,0.60908675,1.1947471,1.7804074,2.366068,2.951728,3.8380275,4.728231,5.618435,6.5086384,7.3988423,7.60968,7.8205175,8.031356,8.238289,8.449126,7.297328,6.1455293,4.9937305,3.8419318,2.6862288,2.1708477,1.6593709,1.1439898,0.62860876,0.113227665,0.7106012,1.3118792,1.9131571,2.514435,3.1118085,2.67842,2.2489357,1.815547,1.3821584,0.94876975,2.35045,3.7482262,5.1499066,6.551587,7.9493628,6.813182,5.6730967,4.5369153,3.4007344,2.260649,2.514435,2.7682211,3.018103,3.2718892,3.5256753,4.095718,4.6657605,5.2358036,5.805846,6.375889,5.9815445,5.5832953,5.1889505,4.794606,4.4002614,4.0918136,3.7833657,3.4788225,3.1703746,2.8619268,3.4319696,4.0020123,4.572055,5.142098,5.7121406,5.989353,6.266566,6.5437784,6.8209906,7.098203,7.773665,8.449126,9.124588,9.80005,10.475512,9.597021,8.718531,7.843944,6.9654536,6.086963,5.700427,5.3138914,4.9234514,4.5369153,4.1503797,4.646239,5.1460023,5.6418614,6.141625,6.6374836,5.7824197,4.927356,4.0722914,3.2172275,2.3621633,2.1083772,1.8506867,1.5969005,1.3431144,1.0893283,1.3431144,1.6008049,1.8584955,2.1161861,2.3738766,2.25284,2.1318035,2.0068626,1.8858263,1.7608855,2.084951,2.4090161,2.7291772,3.0532427,3.3734035,4.0605783,4.7516575,5.4388323,6.126007,6.813182,6.395411,5.9776397,5.559869,5.142098,4.7243266,4.1308575,3.541293,2.9478238,2.3543546,1.7608855,1.7140326,1.6632754,1.6125181,1.5617609,1.5110037,1.5305257,1.5461433,1.5656652,1.5812829,1.6008049,1.737459,1.8741131,2.0107672,2.1513257,2.2879796,2.0615244,1.8389735,1.6125181,1.3860629,1.1635119,1.5812829,2.0029583,2.4207294,2.8424048,3.2640803,4.2362766,5.2084727,6.180669,7.152865,8.125061,7.676055,7.230953,6.7819467,6.336845,5.8878384,5.462259,5.036679,4.6110992,4.1894236,3.7638438,3.5608149,3.357786,3.154757,2.951728,2.7486992,2.5534792,2.358259,2.1669433,1.9717231,1.7765031,1.999054,2.2255092,2.4519646,2.6745155,2.900971,2.612045,2.3231194,2.0380979,1.7491722,1.4641509,1.1713207,0.8823949,0.59346914,0.30063897,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.08589685,0.12103647,0.15617609,0.19131571,0.22645533,1.0034313,1.7843118,2.5651922,3.3460727,4.123049,4.806319,5.4895897,6.17286,6.8561306,7.5394006,6.141625,4.743849,3.3460727,1.9482968,0.5505207,0.46852827,0.38653582,0.30063897,0.21864653,0.13665408,0.12103647,0.10151446,0.08589685,0.06637484,0.05075723,0.15227169,0.25378615,0.359205,0.46071947,0.5622339,0.62860876,0.698888,0.76526284,0.8316377,0.9019169,0.9878138,1.0737107,1.1635119,1.2494087,1.33921,1.1088502,0.8823949,0.6559396,0.42557985,0.19912452,0.39824903,0.60127795,0.80040246,0.999527,1.1986516,1.0502841,0.9019169,0.74964523,0.60127795,0.44900626,0.3709182,0.28892577,0.21083772,0.12884527,0.05075723,0.10932326,0.1717937,0.23035973,0.28892577,0.3513962,0.3318742,0.31625658,0.29673457,0.28111696,0.26159495,0.25378615,0.24597734,0.23816854,0.23426414,0.22645533,1.6554666,3.084478,4.513489,5.9464045,7.375416,5.903456,4.4314966,2.9556324,1.4836729,0.011713207,0.05466163,0.09761006,0.14055848,0.1835069,0.22645533,0.19912452,0.1756981,0.14836729,0.12494087,0.10151446,2.455869,4.814128,7.172387,9.530646,11.888905,9.987461,8.086017,6.1884775,4.2870336,2.3855898,2.0537157,1.717937,1.3821584,1.0463798,0.7106012,0.74574083,0.77697605,0.80821127,0.8433509,0.8745861,0.80040246,0.7262188,0.6481308,0.57394713,0.4997635,0.5309987,0.5583295,0.58956474,0.62079996,0.6481308,1.9561055,3.260176,4.564246,5.8683167,7.1762915,10.436467,13.700547,16.960724,20.224804,23.488884,22.82904,22.169195,21.509352,20.845604,20.18576,20.006157,19.82265,19.639143,19.455637,19.276033,21.45469,23.633347,25.815908,27.994564,30.173222,31.278166,32.383114,33.491962,34.59691,35.701855,32.387016,29.076084,25.761246,22.450314,19.13938,17.956347,16.777216,15.598087,14.418958,13.235924,11.584361,9.928895,8.273428,6.617962,4.9624953,5.056201,5.153811,5.2475166,5.3412223,5.4388323,5.7316628,6.0205884,6.3134184,6.606249,6.899079,6.094772,5.290465,4.4861584,3.6818514,2.87364,3.5725281,4.271416,4.9663997,5.6652875,6.364176,6.551587,6.7389984,6.9264097,7.113821,7.3012323,8.175818,9.050405,9.924991,10.799577,11.674163,10.877665,10.081166,9.280765,8.484266,7.687768,6.17286,4.657952,3.1430438,1.6281357,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.07418364,0.07027924,0.06637484,0.06637484,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3435874,0.6832704,1.0268579,1.3704453,1.7140326,1.3782539,1.0463798,0.7145056,0.38263142,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.19131571,0.37872702,0.5700427,0.76135844,0.94876975,0.76135844,0.5700427,0.37872702,0.19131571,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.62079996,1.2415999,1.8584955,2.4792955,3.1000953,2.7096553,2.3192148,1.9287747,1.5383345,1.1517987,2.330928,3.5100577,4.689187,5.8683167,7.0513506,6.5359693,6.0244927,5.5130157,5.001539,4.4861584,7.9610763,11.435994,14.9109125,18.38583,21.860748,20.646479,19.428307,18.210133,16.991959,15.773785,12.958711,10.139732,7.320754,4.50568,1.6867018,1.8311646,1.9717231,2.1161861,2.2567444,2.4012074,1.9209659,1.4446288,0.96829176,0.49195468,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1756981,0.3553006,0.5309987,0.7106012,0.8862993,5.1460023,9.4018,13.661504,17.917301,22.1731,18.48344,14.789876,11.096312,7.406651,3.7130866,2.9946766,2.2762666,1.5617609,0.8433509,0.12494087,0.10932326,0.093705654,0.078088045,0.06637484,0.05075723,0.48414588,0.9136301,1.3470187,1.7804074,2.2137961,2.8814487,3.5491016,4.2167544,4.884407,5.548156,5.708236,5.8644123,6.0205884,6.180669,6.336845,5.708236,5.0757227,4.447114,3.8185053,3.1859922,2.5690966,1.9522011,1.3353056,0.71841,0.10151446,1.2142692,2.3231194,3.435874,4.548629,5.661383,4.8219366,3.9824903,3.1430438,2.3035975,1.4641509,2.5495746,3.638903,4.7243266,5.813655,6.899079,6.098676,5.298274,4.5017757,3.7013733,2.900971,3.0415294,3.1859922,3.3265507,3.4710135,3.611572,3.978586,4.3416953,4.7087092,5.0718184,5.4388323,5.1460023,4.8570766,4.5681505,4.279225,3.9863946,3.6584249,3.3343596,3.0063896,2.67842,2.35045,3.1781836,4.0059166,4.83365,5.661383,6.4891167,7.0318284,7.570636,8.113348,8.65606,9.198771,9.776623,10.350571,10.924518,11.498465,12.076316,11.2446785,10.416945,9.585307,8.75367,7.9259367,7.336372,6.7507114,6.1611466,5.575486,4.985922,5.181142,5.376362,5.571582,5.7668023,5.9620223,5.2279944,4.493967,3.7560349,3.0220075,2.2879796,2.0146716,1.7413634,1.4680552,1.1986516,0.92534333,1.1908426,1.456342,1.7218413,1.9834363,2.2489357,2.1786566,2.1083772,2.0380979,1.9717231,1.901444,2.1200905,2.338737,2.5612879,2.7799344,2.998581,3.6232853,4.251894,4.8765984,5.5013027,6.126007,5.8292727,5.5286336,5.2318993,4.9351645,4.6384296,4.138666,3.6428072,3.1430438,2.6471848,2.1513257,2.0615244,1.9756275,1.8858263,1.7999294,1.7140326,1.6867018,1.6593709,1.6281357,1.6008049,1.5734742,1.7257458,1.8741131,2.0263848,2.174752,2.3231194,2.1239948,1.9248703,1.7257458,1.5266213,1.3235924,1.8389735,2.3543546,2.8697357,3.3851168,3.900498,4.7828927,5.6652875,6.547683,7.4300776,8.312472,7.8283267,7.348085,6.8639393,6.3836975,5.899552,5.6730967,5.4505453,5.22409,5.001539,4.775084,4.4314966,4.0918136,3.7482262,3.4046388,3.0610514,2.9868677,2.9087796,2.8306916,2.7526035,2.6745155,2.7252727,2.77603,2.8267872,2.87364,2.9243972,2.639376,2.35045,2.0615244,1.7765031,1.4875772,1.1947471,0.9019169,0.60908675,0.31625658,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.12103647,0.20302892,0.28502136,0.3670138,0.44900626,1.097137,1.7452679,2.3933985,3.0415294,3.6857557,4.552533,5.4193106,6.282183,7.1489606,8.011833,6.504734,4.997635,3.4905357,1.9834363,0.47633708,0.40996224,0.3435874,0.28111696,0.21474212,0.14836729,0.12884527,0.10541886,0.08199245,0.058566034,0.039044023,0.25378615,0.47243267,0.6910792,0.9058213,1.1244678,1.0346665,0.94486535,0.8550641,0.76526284,0.6754616,0.81211567,0.94876975,1.0893283,1.2259823,1.3626363,1.1205635,0.8784905,0.63641757,0.39434463,0.14836729,0.30063897,0.44900626,0.60127795,0.74964523,0.9019169,0.78868926,0.6754616,0.5622339,0.44900626,0.3357786,0.28892577,0.24207294,0.19522011,0.14836729,0.10151446,0.14446288,0.19131571,0.23426414,0.28111696,0.3240654,0.30063897,0.28111696,0.25769055,0.23426414,0.21083772,0.23426414,0.25769055,0.28111696,0.30063897,0.3240654,1.3860629,2.4441557,3.506153,4.564246,5.6262436,4.50568,3.3851168,2.2645533,1.1439898,0.023426414,0.058566034,0.093705654,0.12884527,0.1639849,0.19912452,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,3.3148375,6.493021,9.671205,12.849388,16.023666,13.224211,10.424754,7.6252975,4.825841,2.0263848,1.7296503,1.43682,1.1400855,0.8433509,0.5505207,0.78868926,1.0307622,1.2689307,1.5110037,1.7491722,1.475864,1.1986516,0.92534333,0.6481308,0.37482262,0.5583295,0.74574083,0.92924774,1.116659,1.3001659,2.2489357,3.193801,4.142571,5.0913405,6.036206,9.362757,12.689307,16.011953,19.338505,22.66115,21.193096,19.721136,18.25308,16.78112,15.313066,16.82407,18.33117,19.842173,21.353176,22.86418,24.785145,26.706112,28.630981,30.551949,32.476818,32.43387,32.394825,32.35578,32.31674,32.27379,29.689075,27.100456,24.511837,21.923218,19.338505,18.202324,17.066143,15.933866,14.797685,13.661504,12.212971,10.768341,9.319808,7.871275,6.426646,6.3524623,6.278279,6.2079997,6.133816,6.0635366,6.446168,6.832704,7.2192397,7.601871,7.988407,7.328563,6.6687193,6.008875,5.349031,4.689187,5.2436123,5.801942,6.3602715,6.918601,7.47693,7.773665,8.074304,8.374943,8.675582,8.976221,9.237816,9.499411,9.761005,10.0265045,10.2881,10.319335,10.346666,10.377901,10.409137,10.436467,8.382751,6.329036,4.271416,2.2177005,0.1639849,0.12884527,0.09761006,0.06637484,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.08199245,0.078088045,0.07418364,0.06637484,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6832704,1.3704453,2.0537157,2.7408905,3.4241607,2.7604125,2.096664,1.4290112,0.76526284,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.37872702,0.76135844,1.1400855,1.5188124,1.901444,1.5188124,1.1400855,0.76135844,0.37872702,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.46462387,0.92924774,1.3938715,1.8584955,2.3231194,2.0459068,1.7647898,1.4836729,1.2064602,0.92534333,2.3231194,3.7208953,5.1186714,6.5164475,7.914223,7.387129,6.8639393,6.336845,5.813655,5.2865605,8.413987,11.537509,14.661031,17.788456,20.911978,19.877312,18.842646,17.80798,16.773312,15.738646,13.06413,10.393518,7.719003,5.0483923,2.3738766,2.4597735,2.5456703,2.631567,2.7135596,2.7994564,2.2450314,1.6906061,1.1361811,0.58175594,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21083772,0.42167544,0.62860876,0.8394465,1.0502841,4.056674,7.0591593,10.065549,13.0719385,16.074425,13.392099,10.709775,8.027451,5.3451266,2.6628022,2.1669433,1.6710842,1.1791295,0.6832704,0.18741131,0.1639849,0.14055848,0.12103647,0.09761006,0.07418364,0.3553006,0.63641757,0.9136301,1.1947471,1.475864,1.9209659,2.366068,2.8111696,3.2562714,3.7013733,3.8067923,3.9083066,4.0137253,4.1191444,4.224563,4.1191444,4.009821,3.9044023,3.795079,3.6857557,2.9673457,2.2489357,1.5266213,0.80821127,0.08589685,1.7140326,3.338264,4.9624953,6.5867267,8.210958,6.9654536,5.716045,4.4705405,3.2211318,1.9756275,2.7486992,3.5256753,4.298747,5.0757227,5.8487945,5.388075,4.9234514,4.462732,3.998108,3.5373883,3.5686235,3.6037633,3.6349986,3.6662338,3.7013733,3.8614538,4.0215344,4.181615,4.3416953,4.5017757,4.3143644,4.1308575,3.9434462,3.7599394,3.5764325,3.2289407,2.8814487,2.533957,2.1864653,1.8389735,2.9243972,4.0059166,5.0913405,6.1767645,7.262188,8.070399,8.878611,9.686822,10.491129,11.29934,11.775677,12.24811,12.724447,13.200784,13.673217,12.892336,12.111456,11.326671,10.545791,9.761005,8.976221,8.187531,7.3988423,6.6140575,5.825368,5.716045,5.610626,5.5013027,5.395884,5.2865605,4.6735697,4.056674,3.4436827,2.8267872,2.2137961,1.9209659,1.6320401,1.3431144,1.0541886,0.76135844,1.0346665,1.3079748,1.5812829,1.8506867,2.1239948,2.1083772,2.0888553,2.0732377,2.0537157,2.0380979,2.15523,2.2723622,2.3894942,2.5066261,2.6237583,3.1859922,3.7482262,4.3143644,4.8765984,5.4388323,5.2592297,5.083532,4.903929,4.728231,4.548629,4.1464753,3.7443218,3.3421683,2.9400148,2.5378613,2.4129205,2.2879796,2.1630387,2.0380979,1.9131571,1.8389735,1.7686942,1.6945106,1.6242313,1.5500476,1.7140326,1.8741131,2.0380979,2.1981785,2.3621633,2.1864653,2.0107672,1.8389735,1.6632754,1.4875772,2.096664,2.7057507,3.3187418,3.9278288,4.5369153,5.3295093,6.1221027,6.914696,7.70729,8.499884,7.9805984,7.465217,6.9459314,6.4305506,5.911265,5.8878384,5.8644123,5.8370814,5.813655,5.786324,5.3060827,4.8219366,4.3416953,3.8575494,3.3734035,3.416352,3.455396,3.49444,3.533484,3.5764325,3.4514916,3.3265507,3.2016098,3.076669,2.951728,2.6628022,2.3738766,2.0888553,1.7999294,1.5110037,1.2181735,0.92143893,0.62860876,0.3318742,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.15617609,0.28502136,0.41386664,0.5466163,0.6754616,1.1908426,1.7062237,2.2216048,2.7330816,3.2484627,4.298747,5.3451266,6.3915067,7.4417906,8.488171,6.871748,5.251421,3.6349986,2.018576,0.39824903,0.3513962,0.30454338,0.25769055,0.21083772,0.1639849,0.13665408,0.10932326,0.078088045,0.05075723,0.023426414,0.359205,0.6910792,1.0229534,1.3548276,1.6867018,1.4407244,1.1908426,0.94486535,0.698888,0.44900626,0.63641757,0.8238289,1.0112402,1.1986516,1.3860629,1.1283722,0.8706817,0.61689556,0.359205,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.60127795,0.5231899,0.44900626,0.37482262,0.30063897,0.22645533,0.21083772,0.19522011,0.1796025,0.1639849,0.14836729,0.1796025,0.21083772,0.23816854,0.26940376,0.30063897,0.27330816,0.24597734,0.21864653,0.19131571,0.1639849,0.21474212,0.26940376,0.32016098,0.3709182,0.42557985,1.116659,1.8038338,2.494913,3.1859922,3.873167,3.1079042,2.338737,1.5734742,0.80430686,0.039044023,0.06637484,0.093705654,0.12103647,0.14836729,0.1756981,0.1756981,0.1756981,0.1756981,0.1756981,0.1756981,4.173806,8.16801,12.166118,16.164225,20.162333,16.46096,12.763491,9.062118,5.3607445,1.6632754,1.4055848,1.1517987,0.8980125,0.6442264,0.38653582,0.8355421,1.2806439,1.7296503,2.1786566,2.6237583,2.1513257,1.6749885,1.1986516,0.7262188,0.24988174,0.58956474,0.92924774,1.2689307,1.6086137,1.9482968,2.541766,3.1313305,3.7208953,4.31046,4.900025,8.289046,11.674163,15.063184,18.448301,21.837322,19.557152,17.27698,14.996809,12.716639,10.436467,13.641981,16.843592,20.0452,23.24681,26.448421,28.1156,29.778875,31.446056,33.10933,34.776512,33.589573,32.40654,31.2196,30.036566,28.849628,26.987228,25.124828,23.262428,21.400028,19.537628,18.448301,17.358973,16.26574,15.176412,14.087084,12.845484,11.607788,10.366188,9.128492,7.8868923,7.648724,7.406651,7.168483,6.9264097,6.688241,7.164578,7.6409154,8.121157,8.597494,9.073831,8.55845,8.043069,7.531592,7.016211,6.5008297,6.918601,7.336372,7.7541428,8.171914,8.58578,8.999647,9.413514,9.823476,10.237343,10.651209,10.299813,9.948417,9.600925,9.249529,8.898132,9.757101,10.61607,11.471134,12.330102,13.189071,10.592644,7.996216,5.4036927,2.8072653,0.21083772,0.1717937,0.12884527,0.08589685,0.042948425,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.093705654,0.08589685,0.078088045,0.07027924,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0268579,2.0537157,3.0805733,4.1113358,5.138193,4.138666,3.1430438,2.1435168,1.1478943,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.5700427,1.1400855,1.7101282,2.280171,2.8502135,2.280171,1.7101282,1.1400855,0.5700427,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.30844778,0.62079996,0.92924774,1.2415999,1.5500476,1.3782539,1.2103647,1.038571,0.8706817,0.698888,2.3153105,3.9317331,5.5442514,7.1606736,8.773191,8.238289,7.699481,7.1606736,6.6257706,6.086963,8.862993,11.639023,14.411149,17.18718,19.96321,19.108145,18.256985,17.405825,16.55076,15.699601,13.173453,10.6434,8.117252,5.591104,3.0610514,3.0883822,3.1157131,3.1469483,3.174279,3.2016098,2.5690966,1.9365835,1.3040704,0.6715572,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24207294,0.48414588,0.7262188,0.96829176,1.2142692,2.9634414,4.716518,6.4695945,8.2226715,9.975748,8.300759,6.629675,4.958591,3.2836022,1.6125181,1.33921,1.0659018,0.79649806,0.5231899,0.24988174,0.21864653,0.19131571,0.16008049,0.12884527,0.10151446,0.22645533,0.3553006,0.48414588,0.60908675,0.737932,0.96048295,1.183034,1.4055848,1.6281357,1.8506867,1.901444,1.9561055,2.0068626,2.0615244,2.1122816,2.5261483,2.9439192,3.357786,3.7716527,4.1894236,3.3655949,2.541766,1.7218413,0.8980125,0.07418364,2.2137961,4.349504,6.4891167,8.624825,10.764437,9.108971,7.453504,5.7980375,4.142571,2.4871042,2.951728,3.4124475,3.873167,4.337791,4.7985106,4.6735697,4.548629,4.423688,4.298747,4.173806,4.095718,4.0215344,3.9434462,3.8653584,3.78727,3.7443218,3.697469,3.6506162,3.6076677,3.5608149,3.4827268,3.4007344,3.3226464,3.240654,3.1625657,2.795552,2.4285383,2.0615244,1.6906061,1.3235924,2.6667068,4.009821,5.3529353,6.6960497,8.039165,9.108971,10.182681,11.256392,12.326198,13.399908,13.774731,14.149553,14.524376,14.899199,15.274021,14.539994,13.805966,13.0719385,12.334006,11.599979,10.612165,9.6243515,8.636538,7.648724,6.66091,6.250948,5.840986,5.4310236,5.0210614,4.6110992,4.1191444,3.6232853,3.1274261,2.631567,2.135708,1.8311646,1.5227169,1.2142692,0.9058213,0.60127795,0.8784905,1.1596074,1.4407244,1.7218413,1.999054,2.0341935,2.069333,2.1044729,2.1396124,2.174752,2.1903696,2.2059872,2.2216048,2.233318,2.2489357,2.7486992,3.2484627,3.7482262,4.251894,4.7516575,4.6930914,4.6345253,4.575959,4.521298,4.462732,4.154284,3.8458362,3.541293,3.232845,2.9243972,2.7643168,2.6003318,2.436347,2.2762666,2.1122816,1.9951496,1.8780174,1.7608855,1.6437533,1.5266213,1.698415,1.8741131,2.0498111,2.2255092,2.4012074,2.2489357,2.1005683,1.9482968,1.7999294,1.6515622,2.3543546,3.0610514,3.7638438,4.4705405,5.173333,5.8761253,6.578918,7.28171,7.984503,8.687295,8.136774,7.5823493,7.0318284,6.477403,5.9268827,6.098676,6.2743745,6.4500723,6.6257706,6.801469,6.1767645,5.5559645,4.93126,4.31046,3.6857557,3.8458362,4.0020123,4.1581883,4.318269,4.474445,4.173806,3.873167,3.5764325,3.2757936,2.9751544,2.6862288,2.4012074,2.1122816,1.8233559,1.5383345,1.2415999,0.94096094,0.6442264,0.3474918,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.19131571,0.3670138,0.5466163,0.7223144,0.9019169,1.2806439,1.6632754,2.0459068,2.4285383,2.8111696,4.041056,5.270943,6.5008297,7.7307167,8.960603,7.2348576,5.5091114,3.7794614,2.0537157,0.3240654,0.29673457,0.26549935,0.23426414,0.20693332,0.1756981,0.14055848,0.10932326,0.078088045,0.046852827,0.011713207,0.46071947,0.9058213,1.3548276,1.8038338,2.2489357,1.8467822,1.4407244,1.0346665,0.62860876,0.22645533,0.46071947,0.698888,0.93705654,1.175225,1.4133936,1.1400855,0.8667773,0.59346914,0.3240654,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.30063897,0.26159495,0.22645533,0.18741131,0.14836729,0.113227665,0.12884527,0.14836729,0.1639849,0.1835069,0.19912452,0.21474212,0.23035973,0.24597734,0.26159495,0.27330816,0.24207294,0.21083772,0.1756981,0.14446288,0.113227665,0.19522011,0.27721256,0.359205,0.44119745,0.5231899,0.8433509,1.1635119,1.4836729,1.8038338,2.1239948,1.7101282,1.2962615,0.8784905,0.46462387,0.05075723,0.07027924,0.08980125,0.10932326,0.12884527,0.14836729,0.1639849,0.1756981,0.18741131,0.19912452,0.21083772,5.02887,9.846903,14.664935,19.482967,24.300999,19.701614,15.098324,10.498938,5.899552,1.3001659,1.0854238,0.8706817,0.6559396,0.44119745,0.22645533,0.8784905,1.53443,2.1903696,2.8463092,3.4983444,2.8267872,2.1513257,1.475864,0.80040246,0.12494087,0.62079996,1.116659,1.6086137,2.1044729,2.6003318,2.8306916,3.0649557,3.2992198,3.5295796,3.7638438,7.211431,10.662923,14.114414,17.562002,21.013493,17.921206,14.832824,11.740538,8.652155,5.563773,10.455989,15.35211,20.24823,25.14435,30.036566,31.446056,32.85164,34.26113,35.666714,37.076202,34.745277,32.41435,30.08342,27.756395,25.425468,24.289286,23.1492,22.01302,20.876839,19.736753,18.694279,17.647898,16.601519,15.559043,14.512663,13.477997,12.447234,11.416472,10.381805,9.351044,8.941081,8.535024,8.128965,7.719003,7.3129454,7.882988,8.453031,9.023073,9.593117,10.163159,9.792241,9.421323,9.054309,8.683391,8.312472,8.589685,8.866898,9.14411,9.421323,9.698535,10.22563,10.748819,11.275913,11.799104,12.326198,11.361811,10.401327,9.43694,8.476458,7.5120697,9.198771,10.881569,12.568271,14.251068,15.93777,12.802535,9.6673,6.532065,3.39683,0.26159495,0.21083772,0.15617609,0.10541886,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.10151446,0.093705654,0.08199245,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.3704453,2.7408905,4.1113358,5.481781,6.8483214,5.520825,4.1894236,2.8580225,1.5305257,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.76135844,1.5188124,2.280171,3.0415294,3.7989833,3.0415294,2.280171,1.5188124,0.76135844,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.15617609,0.30844778,0.46462387,0.62079996,0.77307165,0.7145056,0.6559396,0.59346914,0.5349031,0.47633708,2.3075018,4.138666,5.9737353,7.8049,9.636065,9.085544,8.538928,7.988407,7.437886,6.8873653,9.311999,11.736633,14.161267,16.585901,19.010534,18.342882,17.671324,17.003672,16.332115,15.660558,13.2788725,10.897186,8.515501,6.133816,3.7482262,3.7208953,3.68966,3.6584249,3.631094,3.5998588,2.8892577,2.1786566,1.4680552,0.76135844,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.27330816,0.5505207,0.8238289,1.1010414,1.3743496,1.8741131,2.3738766,2.87364,3.3734035,3.873167,3.213323,2.5495746,1.8858263,1.2259823,0.5622339,0.5114767,0.46071947,0.41386664,0.3631094,0.31235218,0.27330816,0.23816854,0.19912452,0.1639849,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.93705654,1.8741131,2.8111696,3.7482262,4.689187,3.7638438,2.8385005,1.9131571,0.9878138,0.062470436,2.7135596,5.3607445,8.011833,10.662923,13.314012,11.248583,9.187058,7.125534,5.0640097,2.998581,3.1508527,3.2992198,3.4514916,3.5998588,3.7482262,3.9629683,4.173806,4.388548,4.5993857,4.814128,4.6267166,4.4393053,4.251894,4.0605783,3.873167,3.6232853,3.3734035,3.1235218,2.87364,2.6237583,2.6510892,2.6745155,2.7018464,2.7252727,2.7486992,2.3621633,1.9756275,1.5890918,1.1986516,0.81211567,2.4129205,4.0137253,5.610626,7.211431,8.812236,10.151445,11.486752,12.825961,14.161267,15.500477,15.773785,16.050997,16.324306,16.601519,16.874826,16.187653,15.500477,14.813302,14.126127,13.438952,12.24811,11.061172,9.874233,8.687295,7.5003567,6.785851,6.0752497,5.3607445,4.650143,3.9356375,3.5608149,3.1859922,2.8111696,2.436347,2.0615244,1.737459,1.4133936,1.0893283,0.76135844,0.43729305,0.7262188,1.0112402,1.3001659,1.5890918,1.8741131,1.9639144,2.0498111,2.135708,2.2255092,2.3114061,2.2255092,2.135708,2.0498111,1.9639144,1.8741131,2.3114061,2.7486992,3.1859922,3.6232853,4.0605783,4.123049,4.1894236,4.251894,4.3143644,4.376835,4.1620927,3.951255,3.736513,3.5256753,3.310933,3.1118085,2.912684,2.7135596,2.514435,2.3114061,2.1513257,1.9873407,1.8233559,1.6632754,1.4992905,1.6867018,1.8741131,2.0615244,2.2489357,2.436347,2.3114061,2.1864653,2.0615244,1.9365835,1.8116426,2.612045,3.4124475,4.21285,5.0132523,5.813655,6.426646,7.0357327,7.648724,8.261715,8.874706,8.289046,7.699481,7.113821,6.524256,5.938596,6.3134184,6.688241,7.0630636,7.437886,7.812709,7.0513506,6.2860875,5.5247293,4.7633705,3.998108,4.2753205,4.548629,4.825841,5.099149,5.376362,4.900025,4.423688,3.951255,3.474918,2.998581,2.7135596,2.4246337,2.135708,1.8506867,1.5617609,1.261122,0.96438736,0.6637484,0.3631094,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22645533,0.44900626,0.6754616,0.9019169,1.1244678,1.3743496,1.6242313,1.8741131,2.1239948,2.3738766,3.78727,5.2006636,6.6140575,8.023546,9.43694,7.601871,5.7628975,3.9239242,2.0888553,0.24988174,0.23816854,0.22645533,0.21083772,0.19912452,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.5622339,1.1244678,1.6867018,2.2489357,2.8111696,2.2489357,1.6867018,1.1244678,0.5622339,0.0,0.28892577,0.57394713,0.8628729,1.1517987,1.43682,1.1517987,0.8628729,0.57394713,0.28892577,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,0.1756981,0.28892577,0.39824903,0.5114767,0.62470436,0.57394713,0.5231899,0.47633708,0.42557985,0.37482262,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.14836729,0.1756981,0.19912452,0.22645533,0.24988174,5.8878384,11.525795,17.163752,22.801708,28.435762,22.938364,17.437061,11.935758,6.4383593,0.93705654,0.76135844,0.58566034,0.41386664,0.23816854,0.062470436,0.92534333,1.7882162,2.6510892,3.513962,4.376835,3.4983444,2.6237583,1.7491722,0.8745861,0.0,0.6481308,1.3001659,1.9482968,2.6003318,3.2484627,3.1235218,2.998581,2.87364,2.7486992,2.6237583,6.13772,9.651682,13.16174,16.675701,20.18576,16.289165,12.388668,8.488171,4.5876727,0.6871748,7.2739015,13.860628,20.45126,27.037985,33.624714,34.776512,35.924404,37.076202,38.2241,39.375896,35.900978,32.42606,28.951143,25.476225,22.001307,21.58744,21.173573,20.76361,20.349745,19.935879,18.936352,17.936825,16.937298,15.93777,14.938243,14.11051,13.286681,12.4628525,11.639023,10.81129,10.237343,9.663396,9.085544,8.511597,7.9376497,8.601398,9.261242,9.924991,10.588739,11.248583,11.0260315,10.799577,10.573121,10.350571,10.124115,10.260769,10.401327,10.537982,10.674636,10.81129,11.4516115,12.08803,12.724447,13.360865,14.001186,12.423808,10.850334,9.276859,7.699481,6.126007,8.636538,11.150972,13.661504,16.175938,18.68647,15.012426,11.338385,7.660437,3.9863946,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.7140326,3.4241607,5.138193,6.8483214,8.562354,6.899079,5.2358036,3.5764325,1.9131571,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.94876975,1.901444,2.8502135,3.7989833,4.7516575,3.7989833,2.8502135,1.901444,0.94876975,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,2.2996929,4.349504,6.3993154,8.449126,10.498938,9.936704,9.37447,8.812236,8.250002,7.687768,9.761005,11.838148,13.911386,15.988527,18.061766,17.573715,17.085665,16.601519,16.113468,15.625418,13.388195,11.150972,8.913751,6.676528,4.4393053,4.349504,4.263607,4.173806,4.087909,3.998108,3.213323,2.4246337,1.6359446,0.8511597,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21864653,0.44119745,0.659844,0.8784905,1.1010414,1.4992905,1.901444,2.2996929,2.7018464,3.1000953,2.5690966,2.0380979,1.5110037,0.98000497,0.44900626,0.40996224,0.3709182,0.3318742,0.28892577,0.24988174,0.24597734,0.23816854,0.23426414,0.23035973,0.22645533,0.57394713,0.92534333,1.2767396,1.6242313,1.9756275,1.7335546,1.4914817,1.2494087,1.0034313,0.76135844,0.60908675,0.45681506,0.30454338,0.15227169,0.0,0.80821127,1.620327,2.4285383,3.240654,4.0488653,3.39683,2.7447948,2.0927596,1.4407244,0.78868926,2.9634414,5.142098,7.320754,9.499411,11.674163,10.006983,8.339804,6.6726236,5.0054436,3.338264,3.6584249,3.978586,4.298747,4.618908,4.939069,4.8883114,4.841459,4.794606,4.747753,4.7009,4.4432096,4.1894236,3.9356375,3.6818514,3.4241607,3.2094188,2.9907722,2.7721257,2.5534792,2.338737,2.3933985,2.4480603,2.5027218,2.5573835,2.612045,2.7447948,2.8775444,3.0102942,3.1430438,3.2757936,4.1308575,4.985922,5.840986,6.6960497,7.551114,8.671678,9.796145,10.916709,12.041177,13.16174,13.458474,13.751305,14.048039,14.34087,14.637604,14.450192,14.262781,14.07537,13.887959,13.700547,12.31058,10.920613,9.530646,8.140678,6.7507114,6.0752497,5.3997884,4.7243266,4.0488653,3.3734035,3.076669,2.77603,2.475391,2.174752,1.8741131,1.678893,1.4797685,1.2806439,1.0854238,0.8862993,1.116659,1.3431144,1.5695697,1.796025,2.0263848,2.0732377,2.1200905,2.1669433,2.2137961,2.260649,2.1708477,2.077142,1.9834363,1.893635,1.7999294,2.1278992,2.455869,2.7838387,3.1118085,3.435874,3.5491016,3.6623292,3.775557,3.8887846,3.998108,3.8497405,3.7013733,3.5491016,3.4007344,3.2484627,3.0532427,2.854118,2.6588979,2.4597735,2.260649,2.1239948,1.9873407,1.8506867,1.7140326,1.5734742,1.698415,1.8194515,1.9443923,2.0654287,2.1864653,2.096664,2.0029583,1.9092526,1.815547,1.7257458,2.5183394,3.310933,4.1035266,4.8961205,5.688714,6.649197,7.6135845,8.574067,9.538455,10.498938,10.034314,9.565785,9.097258,8.628729,8.164105,8.421796,8.679486,8.933272,9.190963,9.448653,9.21439,8.976221,8.738052,8.499884,8.261715,7.758047,7.2543793,6.746807,6.2431393,5.735567,5.1303844,4.521298,3.9161155,3.3070288,2.7018464,2.4792955,2.260649,2.0380979,1.8194515,1.6008049,1.2923572,0.98390937,0.679366,0.3709182,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.1717937,0.19522011,0.21864653,0.23816854,0.26159495,0.21864653,0.1756981,0.13665408,0.093705654,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.1796025,0.359205,0.5388075,0.71841,0.9019169,1.3704453,1.8389735,2.3114061,2.7799344,3.2484627,4.7204223,6.1884775,7.660437,9.128492,10.600452,8.531119,6.46569,4.396357,2.330928,0.26159495,0.23816854,0.21864653,0.19522011,0.1717937,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.44900626,0.9019169,1.3509232,1.7999294,2.2489357,1.7999294,1.3509232,0.9019169,0.44900626,0.0,0.23035973,0.46071947,0.6910792,0.92143893,1.1517987,0.92143893,0.6910792,0.46071947,0.23035973,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.08980125,0.13665408,0.1796025,0.22645533,0.22255093,0.21864653,0.21864653,0.21474212,0.21083772,0.1835069,0.15227169,0.12103647,0.093705654,0.062470436,0.15227169,0.24207294,0.3318742,0.42167544,0.5114767,0.47633708,0.44119745,0.40605783,0.3709182,0.3357786,0.28111696,0.22645533,0.1717937,0.11713207,0.062470436,0.078088045,0.093705654,0.10932326,0.12103647,0.13665408,0.15617609,0.1756981,0.19912452,0.21864653,0.23816854,5.4193106,10.600452,15.785499,20.96664,26.151686,21.083773,16.015858,10.947944,5.8800297,0.81211567,0.6715572,0.5309987,0.39434463,0.25378615,0.113227665,0.78868926,1.4680552,2.1435168,2.822883,3.4983444,2.7994564,2.1005683,1.4016805,0.698888,0.0,0.6637484,1.3235924,1.9873407,2.6510892,3.310933,3.154757,2.998581,2.8385005,2.6823244,2.5261483,7.4964523,12.466757,17.437061,22.40346,27.373764,23.110157,18.84655,14.579038,10.315431,6.0518236,10.498938,14.949956,19.400974,23.84809,28.299107,31.844305,35.385597,38.92689,42.472088,46.013382,40.80491,35.596436,30.387962,25.183395,19.974922,20.205282,20.435642,20.666,20.89636,21.12672,19.639143,18.151566,16.663988,15.176412,13.688834,12.8767185,12.068507,11.256392,10.44818,9.636065,9.194867,8.75367,8.308568,7.8673706,7.426173,8.140678,8.859089,9.577498,10.295909,11.014318,10.729298,10.444276,10.159255,9.874233,9.589212,9.690726,9.792241,9.893755,9.999174,10.100689,11.014318,11.924045,12.837675,13.751305,14.661031,12.845484,11.0260315,9.2104845,7.3910336,5.575486,7.793187,10.0147915,12.236397,14.454097,16.675701,14.130032,11.584361,9.0386915,6.4969254,3.951255,3.2679846,2.5847144,1.901444,1.2181735,0.5388075,0.42948425,0.3240654,0.21474212,0.10932326,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.3743496,2.7486992,4.126953,5.5013027,6.8756523,5.5676775,4.2597027,2.951728,1.6437533,0.3357786,0.27330816,0.21083772,0.14836729,0.08589685,0.023426414,0.79649806,1.5695697,2.3426414,3.1157131,3.8887846,3.1118085,2.330928,1.5539521,0.77697605,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,1.8623998,3.5256753,5.1889505,6.8483214,8.511597,8.320281,8.128965,7.9337454,7.7424297,7.551114,9.21439,10.87376,12.537036,14.200311,15.863586,15.188125,14.516567,13.845011,13.173453,12.497992,11.088503,9.679013,8.269524,6.860035,5.4505453,5.024966,4.5993857,4.173806,3.7482262,3.3265507,2.6706111,2.0146716,1.358732,0.7066968,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1639849,0.3318742,0.4958591,0.659844,0.8238289,1.1244678,1.4251068,1.7257458,2.0263848,2.3231194,1.9287747,1.5305257,1.1322767,0.7340276,0.3357786,0.30844778,0.27721256,0.24597734,0.21864653,0.18741131,0.21474212,0.24207294,0.26940376,0.29673457,0.3240654,1.0502841,1.7765031,2.4988174,3.2250361,3.951255,3.4632049,2.979059,2.494913,2.0107672,1.5266213,1.2181735,0.9136301,0.60908675,0.30454338,0.0,0.6832704,1.3665408,2.0459068,2.7291772,3.4124475,3.0337205,2.6510892,2.2723622,1.893635,1.5110037,3.2172275,4.9234514,6.6257706,8.331994,10.0382185,8.765383,7.492548,6.2197127,4.9468775,3.6740425,4.165997,4.6540475,5.1460023,5.6340523,6.126007,5.8175592,5.5091114,5.2006636,4.8961205,4.5876727,4.263607,3.9434462,3.619381,3.2992198,2.9751544,2.7916477,2.6042364,2.4207294,2.233318,2.0498111,2.135708,2.2216048,2.3035975,2.3894942,2.475391,3.1274261,3.7794614,4.4314966,5.083532,5.735567,5.8487945,5.958118,6.067441,6.1767645,6.2860875,7.195813,8.101635,9.01136,9.917182,10.826907,11.139259,11.455516,11.771772,12.084125,12.400381,12.712734,13.025085,13.337439,13.64979,13.962143,12.369146,10.77615,9.183154,7.5940623,6.001066,5.3607445,4.7243266,4.087909,3.4514916,2.8111696,2.5886188,2.3621633,2.135708,1.9131571,1.6867018,1.6164225,1.5461433,1.475864,1.4055848,1.33921,1.5031948,1.6710842,1.8389735,2.0068626,2.174752,2.182561,2.1903696,2.1981785,2.2059872,2.2137961,2.1161861,2.018576,1.9209659,1.8233559,1.7257458,1.9443923,2.1591344,2.377781,2.5964274,2.8111696,2.9751544,3.1391394,3.2992198,3.4632049,3.6232853,3.5373883,3.4514916,3.3616903,3.2757936,3.1859922,2.9907722,2.7994564,2.6042364,2.4090161,2.2137961,2.1005683,1.9873407,1.8741131,1.7608855,1.6515622,1.7062237,1.7647898,1.8233559,1.8819219,1.9365835,1.8780174,1.8194515,1.756981,1.698415,1.6359446,2.4207294,3.2094188,3.9942036,4.7789884,5.563773,6.8756523,8.187531,9.499411,10.81129,12.123169,11.775677,11.428185,11.080693,10.733202,10.38571,10.526268,10.666827,10.807385,10.947944,11.088503,11.373524,11.66245,11.951375,12.236397,12.525322,11.240774,9.956225,8.671678,7.3832245,6.098676,5.3607445,4.618908,3.8809757,3.1391394,2.4012074,2.2489357,2.096664,1.9443923,1.7882162,1.6359446,1.3235924,1.0073358,0.6910792,0.37872702,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.3435874,0.39044023,0.43338865,0.48024148,0.5231899,0.44119745,0.3553006,0.26940376,0.1835069,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.13665408,0.26940376,0.40605783,0.5388075,0.6754616,1.3665408,2.0537157,2.7447948,3.435874,4.126953,5.6535745,7.180196,8.706817,10.2334385,11.763964,9.464272,7.168483,4.8687897,2.5730011,0.27330816,0.24207294,0.21083772,0.1756981,0.14446288,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.3357786,0.6754616,1.0112402,1.3509232,1.6867018,1.3509232,1.0112402,0.6754616,0.3357786,0.0,0.1717937,0.3435874,0.5192855,0.6910792,0.8628729,0.6910792,0.5192855,0.3435874,0.1717937,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.19522011,0.19131571,0.1835069,0.1796025,0.1756981,0.15227169,0.12884527,0.10932326,0.08589685,0.062470436,0.12884527,0.19912452,0.26549935,0.3318742,0.39824903,0.37872702,0.359205,0.339683,0.32016098,0.30063897,0.25378615,0.20693332,0.15617609,0.10932326,0.062470436,0.078088045,0.09761006,0.113227665,0.13274968,0.14836729,0.1639849,0.1796025,0.19522011,0.21083772,0.22645533,4.9546866,9.679013,14.407245,19.135475,23.863707,19.225277,14.590752,9.956225,5.3217,0.6871748,0.58175594,0.47633708,0.3709182,0.26940376,0.1639849,0.6559396,1.1478943,1.639849,2.1318035,2.6237583,2.1005683,1.5734742,1.0502841,0.5231899,0.0,0.6754616,1.3509232,2.0263848,2.7018464,3.3734035,3.1859922,2.9946766,2.803361,2.6159496,2.4246337,8.85128,15.277926,21.708477,28.135122,34.561768,29.931149,25.304432,20.67381,16.043188,11.412568,13.723974,16.039284,18.35069,20.662096,22.973503,28.912098,34.842884,40.781483,46.71617,52.650864,45.708836,38.770714,31.828688,24.890564,17.948538,18.823124,19.693806,20.568392,21.439074,22.31366,20.338032,18.362404,16.386776,14.411149,12.439425,11.642927,10.84643,10.053836,9.257338,8.460839,8.152391,7.843944,7.531592,7.223144,6.910792,7.6838636,8.456935,9.230007,10.003078,10.77615,10.4286585,10.085071,9.741484,9.393991,9.050405,9.116779,9.183154,9.253433,9.319808,9.386183,10.573121,11.763964,12.950902,14.13784,15.324779,13.263254,11.205634,9.14411,7.08649,5.024966,6.9537406,8.878611,10.807385,12.73616,14.661031,13.247637,11.834243,10.416945,9.0035515,7.5862536,6.2860875,4.9820175,3.6818514,2.377781,1.0737107,0.8589685,0.6442264,0.42948425,0.21474212,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.038571,2.0732377,3.1118085,4.1503797,5.1889505,4.2362766,3.2836022,2.330928,1.3782539,0.42557985,0.3513962,0.27330816,0.19912452,0.12494087,0.05075723,0.6442264,1.2415999,1.8350691,2.4285383,3.0259118,2.4207294,1.815547,1.2103647,0.60518235,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,1.4251068,2.7018464,3.9746814,5.251421,6.524256,6.703859,6.8795567,7.0591593,7.2348576,7.4105554,8.663869,9.913278,11.162686,12.412095,13.661504,12.806439,11.947471,11.088503,10.2334385,9.37447,8.792714,8.210958,7.629202,7.043542,6.461786,5.700427,4.939069,4.173806,3.4124475,2.6510892,2.1278992,1.6047094,1.0815194,0.5583295,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10932326,0.21864653,0.3318742,0.44119745,0.5505207,0.74964523,0.94876975,1.1517987,1.3509232,1.5500476,1.2845483,1.0190489,0.75354964,0.48805028,0.22645533,0.20693332,0.1835069,0.1639849,0.14446288,0.12494087,0.1835069,0.24597734,0.30454338,0.3631094,0.42557985,1.5266213,2.6237583,3.7247996,4.825841,5.9268827,5.196759,4.4705405,3.7443218,3.0141985,2.2879796,1.8311646,1.3743496,0.9136301,0.45681506,0.0,0.5544251,1.1088502,1.6632754,2.2216048,2.77603,2.6667068,2.5612879,2.4519646,2.3465457,2.2372224,3.4710135,4.7009,5.9346914,7.168483,8.398369,7.523783,6.6452928,5.7668023,4.8883114,4.0137253,4.6735697,5.3334136,5.9932575,6.6531014,7.3129454,6.746807,6.1767645,5.610626,5.040583,4.474445,4.084005,3.6935644,3.3031244,2.9165885,2.5261483,2.3738766,2.2216048,2.069333,1.9131571,1.7608855,1.8780174,1.9912452,2.1083772,2.2216048,2.338737,3.5100577,4.6813784,5.8566036,7.027924,8.1992445,7.5667315,6.930314,6.2938967,5.661383,5.024966,5.716045,6.4110284,7.1021075,7.793187,8.488171,8.823949,9.155824,9.491602,9.82738,10.163159,10.975275,11.787391,12.599506,13.411622,14.223738,12.431617,10.6355915,8.839567,7.043542,5.251421,4.650143,4.0488653,3.4514916,2.8502135,2.2489357,2.1005683,1.9482968,1.7999294,1.6515622,1.4992905,1.5578566,1.6164225,1.6710842,1.7296503,1.7882162,1.893635,2.0029583,2.1083772,2.2177005,2.3231194,2.2918842,2.260649,2.2294137,2.194274,2.1630387,2.0615244,1.9561055,1.8545911,1.7530766,1.6515622,1.756981,1.8663043,1.9717231,2.0810463,2.1864653,2.4012074,2.612045,2.8267872,3.0376248,3.2484627,3.2250361,3.2016098,3.174279,3.1508527,3.1235218,2.9322062,2.7408905,2.5456703,2.3543546,2.1630387,2.0732377,1.9873407,1.901444,1.8116426,1.7257458,1.717937,1.7101282,1.7023194,1.6945106,1.6867018,1.6593709,1.6320401,1.6047094,1.5773785,1.5500476,2.3270237,3.1039999,3.8809757,4.661856,5.4388323,7.098203,8.761478,10.424754,12.08803,13.751305,13.520945,13.29449,13.068034,12.841579,12.611219,12.634645,12.658072,12.681499,12.70102,12.724447,13.536563,14.348679,15.160794,15.976814,16.788929,14.723501,12.658072,10.592644,8.527214,6.461786,5.591104,4.716518,3.8458362,2.97125,2.1005683,2.0146716,1.9287747,1.8467822,1.7608855,1.6749885,1.3509232,1.0307622,0.7066968,0.38653582,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08980125,0.1796025,0.26940376,0.359205,0.44900626,0.5192855,0.58566034,0.6520352,0.71841,0.78868926,0.659844,0.5309987,0.40605783,0.27721256,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.08980125,0.1796025,0.26940376,0.359205,0.44900626,1.358732,2.2684577,3.1781836,4.0918136,5.001539,6.5867267,8.16801,9.753197,11.338385,12.923572,10.397423,7.871275,5.3412223,2.815074,0.28892577,0.24597734,0.20302892,0.16008049,0.11713207,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.22645533,0.44900626,0.6754616,0.9019169,1.1244678,0.9019169,0.6754616,0.44900626,0.22645533,0.0,0.113227665,0.23035973,0.3435874,0.46071947,0.57394713,0.46071947,0.3435874,0.23035973,0.113227665,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.1678893,0.16008049,0.15227169,0.14446288,0.13665408,0.12103647,0.10932326,0.093705654,0.078088045,0.062470436,0.10932326,0.15227169,0.19912452,0.24207294,0.28892577,0.28111696,0.27721256,0.27330816,0.26940376,0.26159495,0.22255093,0.1835069,0.14055848,0.10151446,0.062470436,0.08199245,0.10151446,0.12103647,0.14055848,0.1639849,0.1717937,0.1835069,0.19131571,0.20302892,0.21083772,4.4861584,8.757574,13.028991,17.30431,21.575727,17.370686,13.169549,8.968412,4.7633705,0.5622339,0.49195468,0.42167544,0.3513962,0.28111696,0.21083772,0.5192855,0.8277333,1.1361811,1.4407244,1.7491722,1.4016805,1.0502841,0.698888,0.3513962,0.0,0.6871748,1.3743496,2.0615244,2.7486992,3.435874,3.213323,2.9907722,2.7682211,2.5456703,2.3231194,10.2100115,18.093,25.979893,33.866787,41.749775,36.756042,31.758408,26.764677,21.770947,16.773312,16.94901,17.124708,17.300406,17.476105,17.651802,25.979893,34.304077,42.632168,50.96026,59.28835,50.612766,41.94109,33.269413,24.597734,15.926057,17.440966,18.955873,20.470781,21.98569,23.500597,21.036919,18.573242,16.113468,13.64979,11.186112,10.409137,9.628256,8.847376,8.066495,7.2856145,7.1099167,6.9342184,6.754616,6.578918,6.3993154,7.2270484,8.054782,8.882515,9.710248,10.537982,10.131924,9.725866,9.323712,8.917655,8.511597,8.546737,8.577971,8.609207,8.644346,8.675582,10.135828,11.599979,13.06413,14.524376,15.988527,13.68493,11.381332,9.081639,6.7780423,4.474445,6.1103897,7.746334,9.378374,11.014318,12.650263,12.365242,12.08022,11.795199,11.510178,11.225157,9.304191,7.37932,5.4583545,3.533484,1.6125181,1.2884527,0.96829176,0.6442264,0.3240654,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.698888,1.4016805,2.1005683,2.7994564,3.4983444,2.900971,2.3035975,1.7062237,1.1088502,0.5114767,0.42557985,0.3357786,0.24988174,0.1639849,0.07418364,0.49195468,0.9097257,1.3274968,1.7452679,2.1630387,1.7296503,1.2962615,0.8667773,0.43338865,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.9878138,1.8741131,2.7643168,3.6506162,4.5369153,5.083532,5.6340523,6.180669,6.727285,7.2739015,8.113348,8.94889,9.788337,10.6238785,11.4633255,10.42085,9.378374,8.335898,7.2934237,6.250948,6.4969254,6.7389984,6.984976,7.230953,7.47693,6.375889,5.2748475,4.173806,3.076669,1.9756275,1.5851873,1.1947471,0.80430686,0.41386664,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05466163,0.10932326,0.1639849,0.21864653,0.27330816,0.37482262,0.47633708,0.57394713,0.6754616,0.77307165,0.6442264,0.5114767,0.37872702,0.24597734,0.113227665,0.10151446,0.093705654,0.08199245,0.07418364,0.062470436,0.15617609,0.24597734,0.339683,0.43338865,0.5231899,1.999054,3.474918,4.950782,6.426646,7.898606,6.930314,5.958118,4.989826,4.0215344,3.049338,2.4402514,1.8311646,1.2181735,0.60908675,0.0,0.42557985,0.8550641,1.2806439,1.7101282,2.135708,2.3035975,2.4675822,2.631567,2.7994564,2.9634414,3.7208953,4.482254,5.2436123,6.001066,6.7624245,6.278279,5.7980375,5.3138914,4.83365,4.349504,5.181142,6.008875,6.8405128,7.6682463,8.499884,7.6721506,6.844417,6.016684,5.1889505,4.3612175,3.9044023,3.4475873,2.9907722,2.533957,2.0732377,1.9561055,1.8350691,1.7140326,1.5969005,1.475864,1.620327,1.7647898,1.9092526,2.0537157,2.1981785,3.892689,5.5832953,7.277806,8.968412,10.662923,9.280765,7.90251,6.524256,5.142098,3.7638438,4.240181,4.716518,5.196759,5.6730967,6.1494336,6.504734,6.860035,7.2153354,7.570636,7.9259367,9.237816,10.549695,11.861574,13.173453,14.489237,12.490183,10.491129,8.495979,6.4969254,4.5017757,3.9356375,3.3734035,2.8111696,2.2489357,1.6867018,1.6125181,1.5383345,1.4641509,1.3860629,1.3118792,1.4992905,1.6827974,1.8663043,2.0537157,2.2372224,2.2840753,2.330928,2.3816853,2.4285383,2.475391,2.4012074,2.330928,2.2567444,2.1864653,2.1122816,2.0068626,1.8975395,1.7882162,1.6827974,1.5734742,1.5734742,1.5695697,1.5656652,1.5656652,1.5617609,1.8233559,2.0888553,2.35045,2.612045,2.87364,2.912684,2.951728,2.9868677,3.0259118,3.0610514,2.87364,2.6823244,2.4910088,2.3035975,2.1122816,2.0498111,1.9873407,1.9248703,1.8623998,1.7999294,1.7257458,1.6554666,1.5812829,1.5110037,1.43682,1.4407244,1.4485333,1.4524376,1.456342,1.4641509,2.233318,3.0024853,3.7716527,4.5408196,5.3138914,7.3246584,9.339331,11.350098,13.360865,15.375536,15.266212,15.160794,15.051471,14.946052,14.836729,14.743023,14.649317,14.551707,14.458001,14.364296,15.699601,17.03881,18.374117,19.713327,21.048632,18.206228,15.359919,12.513609,9.671205,6.824895,5.8214636,4.814128,3.8106966,2.803361,1.7999294,1.7843118,1.7647898,1.7491722,1.7296503,1.7140326,1.3821584,1.0541886,0.7223144,0.39434463,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12103647,0.23816854,0.359205,0.48024148,0.60127795,0.6910792,0.78088045,0.8706817,0.96048295,1.0502841,0.8784905,0.7106012,0.5388075,0.3709182,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.08980125,0.13665408,0.1796025,0.22645533,1.3548276,2.4831998,3.6154766,4.743849,5.8761253,7.5159745,9.159728,10.803481,12.44333,14.087084,11.330575,8.574067,5.813655,3.057147,0.30063897,0.24597734,0.19522011,0.14055848,0.08980125,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.113227665,0.22645533,0.3357786,0.44900626,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.058566034,0.113227665,0.1717937,0.23035973,0.28892577,0.23035973,0.1717937,0.113227665,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.14055848,0.12884527,0.12103647,0.10932326,0.10151446,0.093705654,0.08589685,0.078088045,0.07027924,0.062470436,0.08589685,0.10932326,0.12884527,0.15227169,0.1756981,0.1835069,0.19522011,0.20693332,0.21474212,0.22645533,0.19131571,0.16008049,0.12884527,0.093705654,0.062470436,0.08589685,0.10932326,0.12884527,0.15227169,0.1756981,0.1796025,0.1835069,0.19131571,0.19522011,0.19912452,4.01763,7.8361354,11.650736,15.469242,19.287746,15.516094,11.748346,7.9766936,4.2089458,0.43729305,0.40215343,0.3670138,0.3318742,0.29673457,0.26159495,0.38653582,0.5075723,0.62860876,0.75354964,0.8745861,0.698888,0.5231899,0.3513962,0.1756981,0.0,0.698888,1.4016805,2.1005683,2.7994564,3.4983444,3.2445583,2.9907722,2.7330816,2.4792955,2.2255092,11.568744,20.908073,30.251308,39.594543,48.93778,43.577034,38.21629,32.855545,27.498705,22.13796,20.174046,18.214037,16.250122,14.286208,12.326198,23.043781,33.76527,44.48676,55.20434,65.925835,55.5206,45.115368,34.710136,24.304905,13.899672,16.058807,18.214037,20.37317,22.5284,24.687536,21.735807,18.787983,15.836256,12.888432,9.936704,9.171441,8.406178,7.6409154,6.8756523,6.114294,6.067441,6.0205884,5.9776397,5.930787,5.8878384,6.7702336,7.6526284,8.535024,9.4174185,10.299813,9.835189,9.370565,8.905942,8.441318,7.9766936,7.9727893,7.968885,7.968885,7.9649806,7.9610763,9.698535,11.435994,13.173453,14.9109125,16.64837,14.106606,11.560935,9.0152645,6.4695945,3.9239242,5.267039,6.610153,7.9532676,9.296382,10.6355915,11.482847,12.326198,13.173453,14.016804,14.864059,12.318389,9.776623,7.2348576,4.6930914,2.1513257,1.7218413,1.2884527,0.8589685,0.42948425,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3631094,0.7262188,1.0893283,1.4485333,1.8116426,1.5695697,1.3274968,1.0854238,0.8433509,0.60127795,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.339683,0.58175594,0.8199245,1.0580931,1.3001659,1.038571,0.78088045,0.5192855,0.26159495,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.5505207,1.0502841,1.5500476,2.0498111,2.5495746,3.4671092,4.3846436,5.3021784,6.2197127,7.137247,7.562827,7.988407,8.413987,8.835662,9.261242,8.03526,6.805373,5.579391,4.3534083,3.1235218,4.1972322,5.270943,6.3407493,7.4144597,8.488171,7.0513506,5.610626,4.173806,2.736986,1.3001659,1.0424755,0.78478485,0.5270943,0.26940376,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,2.475391,4.3260775,6.1767645,8.023546,9.874233,8.663869,7.4495993,6.239235,5.024966,3.8106966,3.049338,2.2879796,1.5266213,0.76135844,0.0,0.30063897,0.60127795,0.9019169,1.1986516,1.4992905,1.9365835,2.3738766,2.8111696,3.2484627,3.6857557,3.9746814,4.263607,4.548629,4.8375545,5.12648,5.036679,4.950782,4.860981,4.775084,4.689187,5.688714,6.688241,7.687768,8.687295,9.686822,8.601398,7.5120697,6.426646,5.337318,4.251894,3.7247996,3.2016098,2.6745155,2.1513257,1.6242313,1.5383345,1.4485333,1.3626363,1.2767396,1.1869383,1.3626363,1.5383345,1.7140326,1.8858263,2.0615244,4.2753205,6.4891167,8.699008,10.912805,13.1266,10.998701,8.874706,6.7507114,4.6267166,2.4988174,2.7643168,3.0259118,3.2875066,3.5491016,3.8106966,4.1894236,4.564246,4.939069,5.3138914,5.688714,7.5003567,9.311999,11.123642,12.939189,14.750832,12.548749,10.350571,8.148487,5.950309,3.7482262,3.2250361,2.7018464,2.174752,1.6515622,1.1244678,1.1244678,1.1244678,1.1244678,1.1244678,1.1244678,1.43682,1.7491722,2.0615244,2.3738766,2.6862288,2.6745155,2.6628022,2.6510892,2.639376,2.6237583,2.514435,2.4012074,2.2879796,2.174752,2.0615244,1.9482968,1.8389735,1.7257458,1.6125181,1.4992905,1.3860629,1.2767396,1.1635119,1.0502841,0.93705654,1.2494087,1.5617609,1.8741131,2.1864653,2.4988174,2.6003318,2.7018464,2.7994564,2.900971,2.998581,2.8111696,2.6237583,2.436347,2.2489357,2.0615244,2.0263848,1.9873407,1.9482968,1.9131571,1.8741131,1.737459,1.6008049,1.4641509,1.3235924,1.1869383,1.2259823,1.261122,1.3001659,1.33921,1.3743496,2.135708,2.900971,3.6623292,4.423688,5.1889505,7.551114,9.913278,12.27544,14.637604,16.999767,17.01148,17.023193,17.03881,17.050524,17.062239,16.8514,16.636658,16.42582,16.211079,16.00024,17.86264,5052.0,21.58744,23.44984,25.31224,21.688955,18.061766,14.438479,10.81129,7.1880045,6.0518236,4.911738,3.775557,2.639376,1.4992905,1.5500476,1.6008049,1.6515622,1.698415,1.7491722,1.4133936,1.0737107,0.737932,0.39824903,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14836729,0.30063897,0.44900626,0.60127795,0.74964523,0.8628729,0.97610056,1.0893283,1.1986516,1.3118792,1.1010414,0.8862993,0.6754616,0.46071947,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.3509232,2.7018464,4.0488653,5.3997884,6.7507114,8.449126,10.151445,11.849861,13.548276,15.250595,12.263727,9.276859,6.2860875,3.2992198,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,3.5491016,6.910792,10.276386,13.638077,16.999767,13.661504,10.323239,6.98888,3.6506162,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.0,0.0,0.0,0.0,0.0,0.7106012,1.4251068,2.135708,2.8502135,3.5608149,3.2757936,2.9868677,2.7018464,2.4129205,2.1239948,12.927476,23.723148,34.52663,45.326206,56.125782,50.398026,44.67417,38.950317,33.226463,27.498705,23.399082,19.29946,15.199838,11.100216,7.000593,20.111576,33.226463,46.337444,59.44843,72.56332,60.42453,48.289646,36.15086,24.012074,11.873287,14.676648,17.476105,20.27556,23.075018,25.874474,22.4386,18.998821,15.562947,12.123169,8.687295,7.9376497,7.1880045,6.4383593,5.688714,4.939069,5.024966,5.1108627,5.2006636,5.2865605,5.376362,6.3134184,7.250475,8.187531,9.124588,10.061645,9.538455,9.01136,8.488171,7.9610763,7.437886,7.3988423,7.363703,7.3246584,7.2856145,7.250475,9.261242,11.275913,13.286681,15.3013525,17.31212,14.524376,11.736633,8.94889,6.1611466,3.3734035,4.423688,5.473972,6.524256,7.57454,8.624825,10.600452,12.576079,14.551707,16.52343,18.499058,15.336493,12.173926,9.01136,5.8487945,2.6862288,2.1513257,1.6125181,1.0737107,0.5388075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.23816854,0.3513962,0.46071947,0.57394713,0.6871748,0.57394713,0.46071947,0.3513962,0.23816854,0.12494087,0.18741131,0.24988174,0.31235218,0.37482262,0.43729305,0.3513962,0.26159495,0.1756981,0.08589685,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.113227665,0.22645533,0.3357786,0.44900626,0.5622339,1.8506867,3.1391394,4.423688,5.7121406,7.000593,7.012306,7.0240197,7.0357327,7.0513506,7.0630636,5.64967,4.2362766,2.8267872,1.4133936,0.0,1.901444,3.7989833,5.700427,7.5979667,9.499411,7.726812,5.950309,4.173806,2.4012074,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,1.9834363,3.4710135,4.9546866,6.4383593,7.9259367,6.9810715,6.036206,5.0913405,4.1464753,3.2016098,2.8463092,2.4910088,2.135708,1.7804074,1.4251068,1.3782539,1.3353056,1.2884527,1.2455044,1.1986516,1.6008049,1.999054,2.4012074,2.7994564,3.2016098,3.4007344,3.6037633,3.8067923,4.009821,4.21285,4.1191444,4.029343,3.9356375,3.8419318,3.7482262,4.5564375,5.3607445,6.165051,6.969358,7.773665,7.191909,6.610153,6.028397,5.446641,4.860981,4.2284675,3.59205,2.9556324,2.3231194,1.6867018,1.5812829,1.4719596,1.3665408,1.2572175,1.1517987,1.2533131,1.358732,1.4641509,1.5695697,1.6749885,3.4436827,5.2162814,6.984976,8.75367,10.526268,8.831758,7.1333427,5.4388323,3.7443218,2.0498111,2.3231194,2.5964274,2.8658314,3.1391394,3.4124475,3.638903,3.8692627,4.095718,4.322173,4.548629,6.001066,7.4495993,8.898132,10.350571,11.799104,10.0382185,8.281238,6.520352,4.759466,2.998581,2.7643168,2.5261483,2.2879796,2.0498111,1.8116426,1.7452679,1.678893,1.6086137,1.542239,1.475864,1.7843118,2.096664,2.4051118,2.7135596,3.0259118,3.0883822,3.154757,3.2211318,3.2836022,3.349977,3.1039999,2.8619268,2.6159496,2.3699722,2.1239948,1.999054,1.8702087,1.7413634,1.6164225,1.4875772,1.3821584,1.2767396,1.1713207,1.0659018,0.96438736,1.2142692,1.4641509,1.7140326,1.9639144,2.2137961,2.3114061,2.4129205,2.514435,2.612045,2.7135596,2.6003318,2.4871042,2.3738766,2.260649,2.1513257,2.1903696,2.2294137,2.2684577,2.3114061,2.35045,2.1630387,1.9756275,1.7882162,1.6008049,1.4133936,1.4290112,1.4407244,1.456342,1.4719596,1.4875772,2.069333,2.6510892,3.2367494,3.8185053,4.4002614,6.446168,8.495979,10.541886,12.591698,14.637604,14.723501,14.813302,14.899199,14.989,15.074897,15.168603,15.258404,15.35211,15.445815,15.535617,17.124708,18.7138,20.298986,21.888079,23.473267,20.607435,17.741604,14.871868,12.006037,9.136301,7.914223,6.688241,5.462259,4.2362766,3.0141985,2.7526035,2.4910088,2.233318,1.9717231,1.7140326,1.4055848,1.097137,0.78868926,0.48414588,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12103647,0.23816854,0.359205,0.48024148,0.60127795,0.6910792,0.78088045,0.8706817,0.96048295,1.0502841,0.8784905,0.7106012,0.5388075,0.3709182,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0815194,2.1591344,3.240654,4.318269,5.3997884,6.75852,8.121157,9.479889,10.838621,12.201257,9.811763,7.426173,5.036679,2.6510892,0.26159495,0.21083772,0.15617609,0.10541886,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.07027924,0.08980125,0.10932326,0.12884527,0.14836729,0.12884527,0.10932326,0.08980125,0.07027924,0.05075723,0.07418364,0.093705654,0.11713207,0.14055848,0.1639849,0.19912452,0.23816854,0.27330816,0.31235218,0.3513962,3.2914112,6.2314262,9.171441,12.111456,15.051471,12.166118,9.280765,6.395411,3.5100577,0.62470436,0.57394713,0.5192855,0.46852827,0.41386664,0.3631094,0.28892577,0.21864653,0.14446288,0.07418364,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.58956474,1.1557031,1.7218413,2.2840753,2.8502135,2.6667068,2.4831998,2.3035975,2.1200905,1.9365835,11.951375,21.962263,31.977055,41.98794,51.99883,46.470196,40.945465,35.416832,29.888199,24.36347,21.415646,18.467823,15.519999,12.572175,9.6243515,19.748466,29.868677,39.992794,50.113003,60.237118,51.99102,43.74883,35.50273,27.256632,19.014439,20.025679,21.036919,22.048159,23.063305,24.074545,21.466404,18.858263,16.254026,13.645885,11.037745,10.733202,10.4286585,10.124115,9.815667,9.511124,8.628729,7.746334,6.8639393,5.9815445,5.099149,5.8683167,6.6335793,7.4027467,8.171914,8.937177,8.870802,8.804427,8.734148,8.667773,8.601398,8.675582,8.749765,8.823949,8.898132,8.976221,10.311526,11.650736,12.986042,14.325252,15.660558,13.302299,10.944039,8.581876,6.223617,3.8614538,4.6969957,5.532538,6.36808,7.2036223,8.039165,9.936704,11.834243,13.731783,15.629322,17.526861,14.848442,12.173926,9.499411,6.824895,4.1503797,3.4241607,2.6940374,1.9678187,1.2415999,0.5114767,0.41386664,0.31235218,0.21083772,0.113227665,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.10151446,0.093705654,0.08199245,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.19131571,0.28111696,0.3709182,0.46071947,0.5505207,0.46071947,0.3709182,0.28111696,0.19131571,0.10151446,0.14836729,0.19912452,0.24988174,0.30063897,0.3513962,0.28111696,0.21083772,0.14055848,0.07027924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08980125,0.1796025,0.26940376,0.359205,0.44900626,1.4797685,2.5105307,3.541293,4.5681505,5.5989127,5.9776397,6.356367,6.7311897,7.1099167,7.4886436,5.989353,4.493967,2.9946766,1.4992905,0.0,1.8389735,3.6818514,5.520825,7.3597984,9.198771,7.473026,5.743376,4.01763,2.2918842,0.5622339,0.5192855,0.47243267,0.42557985,0.38263142,0.3357786,0.26940376,0.20302892,0.13665408,0.06637484,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,1.4953861,2.6159496,3.736513,4.853172,5.9737353,5.298274,4.618908,3.9434462,3.2640803,2.5886188,2.639376,2.6940374,2.7447948,2.7994564,2.8502135,2.4597735,2.069333,1.678893,1.2884527,0.9019169,1.261122,1.6242313,1.9873407,2.35045,2.7135596,2.8306916,2.9478238,3.0649557,3.182088,3.2992198,3.2016098,3.1039999,3.0063896,2.9087796,2.8111696,3.4241607,4.0332475,4.6423345,5.251421,5.8644123,5.786324,5.708236,5.630148,5.55206,5.473972,4.728231,3.9863946,3.240654,2.494913,1.7491722,1.6242313,1.4953861,1.3665408,1.2415999,1.1127546,1.1478943,1.183034,1.2181735,1.2533131,1.2884527,2.6159496,3.9434462,5.270943,6.5984397,7.9259367,6.66091,5.395884,4.1308575,2.8658314,1.6008049,1.8819219,2.1630387,2.4480603,2.7291772,3.0141985,3.0922866,3.174279,3.252367,3.3343596,3.4124475,4.5017757,5.5871997,6.676528,7.7619514,8.85128,7.531592,6.211904,4.8883114,3.5686235,2.2489357,2.2996929,2.35045,2.4012074,2.4480603,2.4988174,2.366068,2.2294137,2.096664,1.9600099,1.8233559,2.1318035,2.4402514,2.7486992,3.0532427,3.3616903,3.506153,3.6467118,3.7911747,3.9317331,4.0761957,3.697469,3.3187418,2.9439192,2.5651922,2.1864653,2.0459068,1.901444,1.7608855,1.6164225,1.475864,1.3782539,1.2806439,1.183034,1.0854238,0.9878138,1.175225,1.3626363,1.5500476,1.737459,1.9248703,2.0263848,2.1239948,2.2255092,2.3231194,2.4246337,2.3855898,2.35045,2.3114061,2.2762666,2.2372224,2.3543546,2.4714866,2.5886188,2.7057507,2.8267872,2.5886188,2.35045,2.1122816,1.8741131,1.6359446,1.6281357,1.6242313,1.6164225,1.6086137,1.6008049,2.0029583,2.4051118,2.8072653,3.2094188,3.611572,5.3451266,7.0786815,8.8083315,10.541886,12.27544,12.439425,12.599506,12.763491,12.923572,13.087557,13.4858055,13.884054,14.278399,14.676648,15.074897,16.386776,17.698656,19.014439,20.326319,21.638197,19.525915,17.417538,15.309161,13.196879,11.088503,9.776623,8.460839,7.1489606,5.8370814,4.5252023,3.9551594,3.3851168,2.815074,2.2450314,1.6749885,1.397776,1.1205635,0.8433509,0.5661383,0.28892577,0.23035973,0.1717937,0.113227665,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08980125,0.1796025,0.26940376,0.359205,0.44900626,0.5192855,0.58566034,0.6520352,0.71841,0.78868926,0.659844,0.5309987,0.40605783,0.27721256,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.80821127,1.620327,2.4285383,3.240654,4.0488653,5.0718184,6.0908675,7.1099167,8.128965,9.151918,7.363703,5.575486,3.78727,1.999054,0.21083772,0.1717937,0.12884527,0.08589685,0.042948425,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.05075723,0.06637484,0.08199245,0.09761006,0.113227665,0.09761006,0.08199245,0.06637484,0.05075723,0.039044023,0.058566034,0.078088045,0.09761006,0.11713207,0.13665408,0.21083772,0.28892577,0.3631094,0.43729305,0.5114767,3.0298162,5.548156,8.066495,10.58093,13.09927,10.666827,8.234385,5.801942,3.3694992,0.93705654,0.8316377,0.7262188,0.62079996,0.5192855,0.41386664,0.3318742,0.24597734,0.1639849,0.08199245,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.46852827,0.8862993,1.3040704,1.7218413,2.135708,2.0615244,1.9834363,1.9053483,1.8272603,1.7491722,10.975275,20.201378,29.423576,38.649677,47.875782,42.546272,37.216763,31.883348,26.55384,21.22433,19.428307,17.636185,15.84016,14.044135,12.24811,19.381453,26.514795,33.64814,40.781483,47.91092,43.561417,39.208008,34.8546,30.50119,26.151686,25.37471,24.601639,23.824663,23.05159,22.274614,20.498112,18.72161,16.941202,15.164699,13.388195,13.528754,13.6693125,13.805966,13.946525,14.087084,12.236397,10.381805,8.531119,6.676528,4.825841,5.423215,6.0205884,6.617962,7.2153354,7.812709,8.203149,8.59359,8.98403,9.370565,9.761005,9.948417,10.135828,10.323239,10.510651,10.698062,11.361811,12.025558,12.689307,13.349152,14.012899,12.08022,10.147541,8.214863,6.282183,4.349504,4.970304,5.591104,6.211904,6.8287997,7.4495993,9.269051,11.088503,12.911859,14.73131,16.55076,14.364296,12.173926,9.987461,7.800996,5.610626,4.6930914,3.7794614,2.8619268,1.9443923,1.0268579,0.8238289,0.62470436,0.42557985,0.22645533,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.093705654,0.08589685,0.078088045,0.07027924,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.14055848,0.21083772,0.27721256,0.3435874,0.41386664,0.3435874,0.27721256,0.21083772,0.14055848,0.07418364,0.113227665,0.14836729,0.18741131,0.22645533,0.26159495,0.21083772,0.15617609,0.10541886,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06637484,0.13665408,0.20302892,0.26940376,0.3357786,1.1088502,1.8819219,2.6549935,3.4280653,4.2011366,4.942973,5.6848097,6.426646,7.168483,7.914223,6.329036,4.747753,3.1664703,1.5812829,0.0,1.7804074,3.5608149,5.3412223,7.1216297,8.898132,7.2192397,5.5403466,3.8614538,2.1786566,0.4997635,0.5349031,0.5700427,0.60518235,0.64032197,0.6754616,0.5388075,0.40605783,0.26940376,0.13665408,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,1.0034313,1.7608855,2.514435,3.2718892,4.025439,3.6154766,3.2055142,2.795552,2.3855898,1.9756275,2.436347,2.893162,3.3538816,3.814601,4.2753205,3.541293,2.803361,2.069333,1.3353056,0.60127795,0.92534333,1.2494087,1.5734742,1.901444,2.2255092,2.2567444,2.2918842,2.3231194,2.3543546,2.3855898,2.2840753,2.182561,2.0810463,1.9756275,1.8741131,2.2918842,2.7057507,3.1196175,3.533484,3.951255,4.376835,4.806319,5.2318993,5.661383,6.086963,5.2318993,4.376835,3.521771,2.6667068,1.8116426,1.6632754,1.5188124,1.3704453,1.2220778,1.0737107,1.038571,1.0034313,0.96829176,0.93315214,0.9019169,1.7843118,2.6706111,3.5569105,4.4393053,5.3256044,4.4900627,3.6545205,2.8189783,1.9834363,1.1517987,1.4407244,1.7335546,2.0263848,2.3192148,2.612045,2.5456703,2.4792955,2.4090161,2.3426414,2.2762666,2.998581,3.7247996,4.4510183,5.173333,5.899552,5.0210614,4.138666,3.260176,2.3816853,1.4992905,1.8389735,2.174752,2.514435,2.8502135,3.1859922,2.9868677,2.7838387,2.5808098,2.377781,2.174752,2.4792955,2.7838387,3.0883822,3.39683,3.7013733,3.9200199,4.138666,4.3612175,4.579864,4.7985106,4.290938,3.7794614,3.2718892,2.7604125,2.2489357,2.0927596,1.9365835,1.7765031,1.620327,1.4641509,1.3743496,1.2806439,1.1908426,1.1010414,1.0112402,1.1361811,1.261122,1.3860629,1.5110037,1.6359446,1.737459,1.8389735,1.9365835,2.0380979,2.135708,2.174752,2.2137961,2.2489357,2.2879796,2.3231194,2.5183394,2.7135596,2.9087796,3.1039999,3.2992198,3.0141985,2.7252727,2.436347,2.1513257,1.8623998,1.8311646,1.8038338,1.7725986,1.7413634,1.7140326,1.9365835,2.1591344,2.3816853,2.6042364,2.8267872,4.2440853,5.661383,7.0786815,8.495979,9.913278,10.151445,10.38571,10.6238785,10.862047,11.100216,11.803008,12.5058,13.208592,13.911386,14.614178,15.648844,16.687416,17.725986,18.760653,19.799223,18.448301,17.093473,15.74255,14.391626,13.036799,11.639023,10.237343,8.835662,7.437886,6.036206,5.1577153,4.279225,3.39683,2.5183394,1.6359446,1.3899672,1.1439898,0.8941081,0.6481308,0.39824903,0.32016098,0.23816854,0.16008049,0.078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.3435874,0.39044023,0.43338865,0.48024148,0.5231899,0.44119745,0.3553006,0.26940376,0.1835069,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5388075,1.0815194,1.620327,2.1591344,2.7018464,3.3812122,4.0605783,4.7399445,5.4193106,6.098676,4.911738,3.7247996,2.5378613,1.3509232,0.1639849,0.12884527,0.09761006,0.06637484,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.046852827,0.039044023,0.03513962,0.031235218,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.03513962,0.046852827,0.05466163,0.06637484,0.07418364,0.06637484,0.05466163,0.046852827,0.03513962,0.023426414,0.042948425,0.058566034,0.078088045,0.093705654,0.113227665,0.22645533,0.3357786,0.44900626,0.5622339,0.6754616,2.7682211,4.8648853,6.9615493,9.054309,11.150972,9.171441,7.191909,5.2084727,3.2289407,1.2494087,1.0932326,0.93315214,0.77697605,0.62079996,0.46071947,0.3709182,0.27721256,0.1835069,0.093705654,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.3435874,0.61689556,0.8862993,1.1557031,1.4251068,1.4524376,1.4797685,1.5070993,1.53443,1.5617609,9.999174,18.436588,26.874,35.311413,43.74883,38.618443,33.484154,28.35377,23.21948,18.089096,17.44487,16.800642,16.16032,15.516094,14.875772,19.018343,23.160913,27.303486,31.446056,35.588627,35.127907,34.667187,34.206467,33.74575,33.288933,30.723742,28.162453,25.601166,23.035973,20.474686,19.525915,18.58105,17.63228,16.683512,15.738646,16.324306,16.906061,17.491722,18.077383,18.663042,15.84016,13.017277,10.194394,7.3715115,4.548629,4.9781127,5.4036927,5.833177,6.2587566,6.688241,7.535496,8.382751,9.230007,10.077262,10.924518,11.225157,11.525795,11.826434,12.123169,12.423808,12.412095,12.400381,12.388668,12.376955,12.361338,10.858143,9.351044,7.8478484,6.3407493,4.8375545,5.2436123,5.645766,6.0518236,6.4578815,6.8639393,8.605303,10.346666,12.091934,13.833297,15.57466,13.8762455,12.173926,10.475512,8.773191,7.0747766,5.9659266,4.860981,3.7521305,2.6432803,1.5383345,1.2376955,0.93705654,0.63641757,0.3357786,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.08199245,0.078088045,0.07418364,0.06637484,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.093705654,0.14055848,0.1835069,0.23035973,0.27330816,0.23035973,0.1835069,0.14055848,0.093705654,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.08980125,0.13665408,0.1796025,0.22645533,0.7418364,1.2533131,1.7686942,2.2840753,2.7994564,3.9083066,5.0132523,6.1221027,7.230953,8.335898,6.6687193,5.001539,3.3343596,1.6671798,0.0,1.7218413,3.4397783,5.1616197,6.8795567,8.601398,6.9654536,5.3334136,3.7013733,2.069333,0.43729305,0.5544251,0.6676528,0.78088045,0.8980125,1.0112402,0.80821127,0.60908675,0.40605783,0.20302892,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.5153811,0.9058213,1.2962615,1.6867018,2.0732377,1.9326792,1.7882162,1.6476578,1.5031948,1.3626363,2.2294137,3.096191,3.9668727,4.83365,5.700427,4.618908,3.541293,2.4597735,1.3782539,0.30063897,0.58566034,0.8745861,1.1635119,1.4485333,1.737459,1.6867018,1.6320401,1.5812829,1.5266213,1.475864,1.3665408,1.261122,1.1517987,1.0463798,0.93705654,1.1557031,1.3782539,1.5969005,1.815547,2.0380979,2.97125,3.9044023,4.83365,5.7668023,6.699954,5.735567,4.7711797,3.8067923,2.8385005,1.8741131,1.7062237,1.5383345,1.3743496,1.2064602,1.038571,0.93315214,0.8277333,0.7223144,0.61689556,0.5114767,0.95657855,1.397776,1.8389735,2.2840753,2.7252727,2.3192148,1.9131571,1.5110037,1.1049459,0.698888,1.0034313,1.3040704,1.6086137,1.9092526,2.2137961,1.999054,1.7843118,1.5656652,1.3509232,1.1361811,1.4992905,1.8623998,2.2255092,2.5886188,2.951728,2.5105307,2.069333,1.6281357,1.1908426,0.74964523,1.3743496,1.999054,2.6237583,3.2484627,3.873167,3.6037633,3.3343596,3.0649557,2.795552,2.5261483,2.8267872,3.1313305,3.4319696,3.736513,4.037152,4.3338866,4.630621,4.93126,5.2279944,5.5247293,4.884407,4.240181,3.5959544,2.9556324,2.3114061,2.1396124,1.9678187,1.796025,1.6242313,1.4485333,1.3665408,1.2845483,1.2025559,1.1205635,1.038571,1.1010414,1.1635119,1.2259823,1.2884527,1.3509232,1.4485333,1.5500476,1.6515622,1.7491722,1.8506867,1.9639144,2.0732377,2.1864653,2.2996929,2.4129205,2.6862288,2.9556324,3.2289407,3.5022488,3.775557,3.435874,3.1000953,2.7643168,2.4246337,2.0888553,2.0341935,1.9834363,1.9287747,1.8780174,1.8233559,1.8663043,1.9092526,1.9522011,1.9951496,2.0380979,3.1391394,4.2440853,5.3451266,6.446168,7.551114,7.8634663,8.175818,8.488171,8.800523,9.112875,10.120211,11.127546,12.134882,13.142218,14.149553,14.9109125,15.676175,16.437534,17.198893,17.964155,17.366781,16.773312,16.175938,15.582469,14.989,13.501423,12.013845,10.526268,9.0386915,7.551114,6.3602715,5.169429,3.978586,2.7916477,1.6008049,1.3821584,1.1635119,0.94876975,0.7301232,0.5114767,0.40996224,0.30844778,0.20693332,0.10151446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.1717937,0.19522011,0.21864653,0.23816854,0.26159495,0.21864653,0.1756981,0.13665408,0.093705654,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26940376,0.5388075,0.80821127,1.0815194,1.3509232,1.6906061,2.0302892,2.3699722,2.7096553,3.049338,2.463678,1.8741131,1.2884527,0.698888,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.019522011,0.015617609,0.015617609,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.015617609,0.023426414,0.027330816,0.031235218,0.039044023,0.031235218,0.027330816,0.023426414,0.015617609,0.011713207,0.027330816,0.042948425,0.058566034,0.07418364,0.08589685,0.23816854,0.38653582,0.5388075,0.6871748,0.8394465,2.5105307,4.181615,5.8566036,7.5276875,9.198771,7.6721506,6.1455293,4.618908,3.0883822,1.5617609,1.3509232,1.1439898,0.93315214,0.7223144,0.5114767,0.40996224,0.30844778,0.20693332,0.10151446,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.22255093,0.3435874,0.46852827,0.58956474,0.7106012,0.8433509,0.97610056,1.1088502,1.2415999,1.3743496,9.026978,16.675701,24.324427,31.97315,39.62578,34.690613,29.75545,24.820286,19.88512,14.949956,15.461433,15.969006,16.480482,16.991959,17.49953,18.651329,19.803127,20.958832,22.11063,23.262428,26.694399,30.126368,33.55834,36.994213,40.42618,36.076675,31.723269,27.373764,23.02426,18.674755,18.557625,18.440493,18.32336,18.206228,18.089096,19.115953,20.146715,21.177479,22.20824,23.239002,19.443924,15.652749,11.861574,8.066495,4.2753205,4.533011,4.7907014,5.0483923,5.3060827,5.563773,6.8678436,8.171914,9.475985,10.783959,12.08803,12.501896,12.911859,13.325725,13.735687,14.149553,13.462379,12.775204,12.08803,11.400854,10.71368,9.636065,8.55845,7.480835,6.4032197,5.3256044,5.5169206,5.704332,5.8956475,6.083059,6.2743745,7.941554,9.60483,11.268105,12.935285,14.59856,13.388195,12.173926,10.963562,9.749292,8.538928,7.238762,5.9425,4.646239,3.3460727,2.0498111,1.6515622,1.2494087,0.8511597,0.44900626,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.07418364,0.07027924,0.06637484,0.06637484,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.046852827,0.07027924,0.093705654,0.113227665,0.13665408,0.113227665,0.093705654,0.07027924,0.046852827,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.3709182,0.62860876,0.8862993,1.1439898,1.4016805,2.87364,4.3455997,5.8175592,7.289519,8.761478,7.008402,5.2592297,3.506153,1.7530766,0.0,1.6593709,3.3187418,4.9781127,6.6413884,8.300759,6.715572,5.1303844,3.5451972,1.9600099,0.37482262,0.5700427,0.76526284,0.96048295,1.1557031,1.3509232,1.0815194,0.80821127,0.5388075,0.26940376,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,0.74964523,2.0263848,3.2992198,4.575959,5.8487945,7.125534,5.700427,4.2753205,2.8502135,1.4251068,0.0,0.24988174,0.4997635,0.74964523,0.999527,1.2494087,1.1127546,0.97610056,0.8394465,0.698888,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,1.5617609,2.998581,4.4393053,5.8761253,7.3129454,6.239235,5.1616197,4.087909,3.0141985,1.9365835,1.7491722,1.5617609,1.3743496,1.1869383,0.999527,0.8238289,0.6481308,0.47633708,0.30063897,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.14836729,0.1756981,0.19912452,0.22645533,0.24988174,0.5622339,0.8745861,1.1869383,1.4992905,1.8116426,1.4485333,1.0893283,0.7262188,0.3631094,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.9136301,1.8233559,2.736986,3.6506162,4.564246,4.224563,3.8887846,3.5491016,3.213323,2.87364,3.174279,3.474918,3.775557,4.0761957,4.376835,4.7516575,5.12648,5.5013027,5.8761253,6.250948,5.473972,4.7009,3.9239242,3.1508527,2.3738766,2.1864653,1.999054,1.8116426,1.6242313,1.43682,1.3626363,1.2884527,1.2142692,1.1361811,1.0619974,1.0619974,1.0619974,1.0619974,1.0619974,1.0619974,1.1635119,1.261122,1.3626363,1.4641509,1.5617609,1.7491722,1.9365835,2.1239948,2.3114061,2.4988174,2.8502135,3.2016098,3.5491016,3.900498,4.251894,3.8614538,3.474918,3.0883822,2.7018464,2.3114061,2.2372224,2.1630387,2.0888553,2.0107672,1.9365835,1.7999294,1.6632754,1.5266213,1.3860629,1.2494087,2.0380979,2.8267872,3.611572,4.4002614,5.1889505,5.575486,5.9620223,6.348558,6.7389984,7.125534,8.437413,9.749292,11.061172,12.376955,13.688834,14.176885,14.661031,15.14908,15.637131,16.125181,16.289165,16.449247,16.613232,16.773312,16.937298,15.363823,13.786445,12.212971,10.6355915,9.062118,7.562827,6.0635366,4.564246,3.0610514,1.5617609,1.3743496,1.1869383,0.999527,0.81211567,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.24988174,0.43729305,0.62470436,0.81211567,0.999527,2.2489357,3.4983444,4.7516575,6.001066,7.250475,6.1767645,5.099149,4.025439,2.951728,1.8741131,1.6125181,1.3509232,1.0893283,0.8238289,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.23816854,0.47633708,0.7106012,0.94876975,1.1869383,8.050878,14.9109125,21.77485,28.63879,35.498825,30.762785,26.026745,21.2868,16.55076,11.810817,13.4740925,15.137367,16.800642,18.463919,20.12329,18.28822,16.449247,14.614178,12.775204,10.936231,18.264793,25.585548,32.914112,40.23877,47.563427,41.42571,35.287987,29.150267,23.012547,16.874826,17.589333,18.299932,19.014439,5052.0,20.435642,21.911505,23.38737,24.863234,26.339098,27.811058,23.05159,18.28822,13.524849,8.761478,3.998108,4.087909,4.173806,4.263607,4.349504,4.4393053,6.2001905,7.9610763,9.725866,11.486752,13.251541,13.774731,14.301826,14.825015,15.348206,15.875299,14.512663,13.150026,11.787391,10.424754,9.062118,8.413987,7.7619514,7.113821,6.461786,5.813655,5.786324,5.7628975,5.735567,5.7121406,5.688714,7.2739015,8.862993,10.44818,12.037272,13.626364,12.900145,12.173926,11.4516115,10.725393,9.999174,8.511597,7.0240197,5.5364423,4.0488653,2.5612879,2.0615244,1.5617609,1.0619974,0.5622339,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.8389735,3.6740425,5.5130157,7.348085,9.187058,7.348085,5.5130157,3.6740425,1.8389735,0.0,1.6008049,3.2016098,4.7985106,6.3993154,8.00012,6.461786,4.9234514,3.3890212,1.8506867,0.31235218,0.58566034,0.8628729,1.1361811,1.4133936,1.6867018,1.3509232,1.0112402,0.6754616,0.3357786,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.60127795,1.6671798,2.7330816,3.802888,4.8687897,5.938596,5.087436,4.2362766,3.3890212,2.5378613,1.6867018,1.6437533,1.6008049,1.5617609,1.5188124,1.475864,1.3353056,1.1947471,1.0541886,0.9136301,0.77307165,0.6637484,0.5505207,0.43729305,0.3240654,0.21083772,0.19131571,0.1717937,0.15227169,0.13274968,0.113227665,1.261122,2.4090161,3.5569105,4.7009,5.8487945,4.9937305,4.138666,3.2836022,2.4285383,1.5734742,1.4212024,1.2650263,1.1088502,0.95657855,0.80040246,0.6637484,0.5309987,0.39434463,0.26159495,0.12494087,0.12103647,0.113227665,0.10932326,0.10541886,0.10151446,0.12103647,0.14055848,0.16008049,0.1796025,0.19912452,0.44900626,0.698888,0.94876975,1.1986516,1.4485333,1.1596074,0.8706817,0.58175594,0.28892577,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7301232,1.4602464,2.1903696,2.920493,3.6506162,3.3812122,3.1118085,2.8385005,2.5690966,2.2996929,2.5495746,2.7994564,3.049338,3.2992198,3.5491016,3.873167,4.2011366,4.5252023,4.8492675,5.173333,4.5837684,3.9942036,3.4046388,2.815074,2.2255092,2.2762666,2.3231194,2.3738766,2.4246337,2.475391,2.233318,1.9951496,1.7530766,1.5149081,1.2767396,1.2494087,1.2259823,1.1986516,1.175225,1.1517987,1.2298868,1.3118792,1.3899672,1.4680552,1.5500476,1.6593709,1.7686942,1.8819219,1.9912452,2.1005683,2.4012074,2.7018464,2.998581,3.2992198,3.5998588,3.377308,3.154757,2.9322062,2.7096553,2.4871042,2.3348327,2.182561,2.0302892,1.8780174,1.7257458,1.5929961,1.4602464,1.3274968,1.1947471,1.0619974,1.7101282,2.358259,3.0063896,3.6506162,4.298747,4.6657605,5.02887,5.395884,5.758993,6.126007,7.309041,8.495979,9.679013,10.865952,12.0489855,12.513609,12.974329,13.438952,13.899672,14.364296,14.446288,14.532186,14.618082,14.703979,14.785972,13.536563,12.28325,11.029937,9.776623,8.52331,7.4417906,6.356367,5.270943,4.185519,3.1000953,2.9946766,2.8892577,2.7838387,2.67842,2.5769055,2.2372224,1.901444,1.5617609,1.2259823,0.8862993,0.7262188,0.5622339,0.39824903,0.23816854,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.21083772,0.359205,0.5036679,0.6520352,0.80040246,1.8194515,2.8345962,3.853645,4.8687897,5.8878384,5.0132523,4.142571,3.2718892,2.397303,1.5266213,1.3235924,1.1205635,0.91753453,0.7145056,0.5114767,0.40996224,0.30844778,0.20693332,0.10151446,0.0,0.042948425,0.08589685,0.12884527,0.1717937,0.21083772,0.1835069,0.15227169,0.12103647,0.093705654,0.062470436,0.23816854,0.41777104,0.59346914,0.77307165,0.94876975,6.871748,12.790822,18.709896,24.62897,30.548042,27.10436,23.660677,20.21309,16.769407,13.325725,13.950429,14.575133,15.199838,15.824542,16.449247,15.629322,14.809398,13.989473,13.169549,12.349625,18.116426,23.879324,29.646126,35.409023,41.175827,36.76385,32.35578,27.943808,23.535736,19.123762,19.326792,19.525915,5052.0,19.924164,20.12329,21.083773,22.04035,22.99693,23.953508,24.91399,21.013493,17.1169,13.220306,9.323712,5.423215,5.1030536,4.786797,4.466636,4.1464753,3.8263142,5.181142,6.5359693,7.890797,9.245625,10.600452,11.018223,11.4398985,11.861574,12.2793455,12.70102,11.62731,10.553599,9.483793,8.410083,7.336372,6.98888,6.6413884,6.2938967,5.9464045,5.5989127,5.6848097,5.7707067,5.8566036,5.938596,6.0244927,7.152865,8.281238,9.405705,10.534078,11.66245,13.068034,14.473619,15.879204,17.280884,18.68647,15.793307,12.90405,10.010887,7.1177254,4.224563,3.9434462,3.6662338,3.3851168,3.1039999,2.8267872,2.3114061,1.7999294,1.2884527,0.77307165,0.26159495,0.21474212,0.1678893,0.12103647,0.07418364,0.023426414,0.023426414,0.019522011,0.015617609,0.015617609,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.03513962,0.046852827,0.05466163,0.06637484,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.4719596,2.9400148,4.40807,5.8800297,7.348085,5.8800297,4.40807,2.9400148,1.4719596,0.0,1.2806439,2.5612879,3.8419318,5.1186714,6.3993154,5.185046,3.970777,2.7565079,1.5383345,0.3240654,0.76916724,1.2103647,1.6515622,2.096664,2.5378613,2.0888553,1.6359446,1.1869383,0.737932,0.28892577,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.44900626,1.3118792,2.1708477,3.0298162,3.8887846,4.7516575,4.474445,4.2011366,3.9239242,3.6506162,3.3734035,3.0415294,2.7057507,2.3699722,2.0341935,1.698415,1.5578566,1.4133936,1.2728351,1.1283722,0.9878138,0.8745861,0.76135844,0.6481308,0.5388075,0.42557985,0.359205,0.29673457,0.23035973,0.1639849,0.10151446,0.95657855,1.815547,2.6706111,3.5295796,4.388548,3.7521305,3.1157131,2.4831998,1.8467822,1.2142692,1.0893283,0.96829176,0.8433509,0.7223144,0.60127795,0.5036679,0.40996224,0.31625658,0.21864653,0.12494087,0.113227665,0.10541886,0.093705654,0.08589685,0.07418364,0.08980125,0.10541886,0.12103647,0.13665408,0.14836729,0.3357786,0.5231899,0.7106012,0.9019169,1.0893283,0.8706817,0.6520352,0.43338865,0.21864653,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5466163,1.0932326,1.6437533,2.1903696,2.736986,2.533957,2.330928,2.1318035,1.9287747,1.7257458,1.9248703,2.1239948,2.3231194,2.5261483,2.7252727,2.998581,3.2757936,3.5491016,3.8263142,4.0996222,3.6935644,3.2914112,2.8853533,2.4792955,2.0732377,2.3621633,2.6510892,2.9361105,3.2250361,3.513962,3.1079042,2.7018464,2.2957885,1.893635,1.4875772,1.43682,1.3860629,1.33921,1.2884527,1.2376955,1.2962615,1.358732,1.4172981,1.475864,1.5383345,1.5695697,1.6008049,1.6359446,1.6671798,1.698415,1.9482968,2.1981785,2.4480603,2.7018464,2.951728,2.893162,2.8345962,2.77603,2.7213683,2.6628022,2.4324427,2.2020829,1.9717231,1.7413634,1.5110037,1.3860629,1.2572175,1.1283722,1.0034313,0.8745861,1.3821584,1.8897307,2.397303,2.9048753,3.4124475,3.7560349,4.095718,4.4393053,4.7828927,5.12648,6.180669,7.238762,8.296855,9.354948,10.413041,10.850334,11.287627,11.72492,12.162213,12.599506,12.607315,12.615124,12.622932,12.630741,12.63855,11.709302,10.77615,9.846903,8.917655,7.988407,7.3168497,6.649197,5.9776397,5.3060827,4.6384296,4.6150036,4.591577,4.5681505,4.548629,4.5252023,3.9746814,3.4241607,2.87364,2.3231194,1.7765031,1.4485333,1.1244678,0.80040246,0.47633708,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.1717937,0.27721256,0.38653582,0.49195468,0.60127795,1.3860629,2.1708477,2.9556324,3.7404175,4.5252023,3.853645,3.1859922,2.514435,1.8467822,1.175225,1.0307622,0.8902037,0.74574083,0.60518235,0.46071947,0.3709182,0.27721256,0.1835069,0.093705654,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.26549935,0.23035973,0.19522011,0.16008049,0.12494087,0.24207294,0.359205,0.47633708,0.59346914,0.7106012,5.688714,10.666827,15.644939,20.623053,25.601166,23.445936,21.29461,19.143284,16.988054,14.836729,14.426766,14.012899,13.599033,13.189071,12.775204,12.974329,13.169549,13.368673,13.563893,13.763018,17.96806,22.1731,26.378141,30.583183,34.788223,32.1059,29.423576,26.741251,24.058928,21.376602,21.06425,20.751898,20.435642,20.12329,19.810938,20.252134,20.693333,21.130625,21.571823,22.01302,18.9793,15.949483,12.915763,9.882042,6.8483214,6.1221027,5.395884,4.6657605,3.9395418,3.213323,4.1581883,5.1069584,6.055728,7.000593,7.9493628,8.265619,8.581876,8.894228,9.2104845,9.526741,8.741957,7.9610763,7.1762915,6.395411,5.610626,5.5676775,5.520825,5.477876,5.4310236,5.388075,5.5832953,5.7785153,5.9737353,6.168956,6.364176,7.0318284,7.6955767,8.36323,9.030883,9.698535,13.235924,16.769407,20.306797,23.84028,27.373764,23.078922,18.780174,14.481428,10.186585,5.8878384,5.8292727,5.7668023,5.708236,5.645766,5.5871997,4.575959,3.5608149,2.5495746,1.5383345,0.5231899,0.42948425,0.3357786,0.23816854,0.14446288,0.05075723,0.046852827,0.039044023,0.03513962,0.031235218,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.058566034,0.06637484,0.07418364,0.078088045,0.08589685,0.08589685,0.08589685,0.08589685,0.08589685,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1010414,2.2059872,3.3070288,4.40807,5.5130157,4.40807,3.3070288,2.2059872,1.1010414,0.0,0.96048295,1.9209659,2.8814487,3.8380275,4.7985106,3.9083066,3.0141985,2.1239948,1.2298868,0.3357786,0.94876975,1.5578566,2.1669433,2.77603,3.3890212,2.8267872,2.260649,1.698415,1.1361811,0.57394713,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.30063897,0.95267415,1.6047094,2.2567444,2.9087796,3.5608149,3.8614538,4.1620927,4.462732,4.7633705,5.0640097,4.435401,3.8067923,3.1781836,2.5534792,1.9248703,1.7804074,1.6359446,1.4914817,1.3431144,1.1986516,1.0893283,0.97610056,0.8628729,0.74964523,0.63641757,0.5270943,0.41777104,0.30844778,0.19912452,0.08589685,0.6559396,1.2220778,1.7882162,2.358259,2.9243972,2.5105307,2.096664,1.678893,1.2650263,0.8511597,0.76135844,0.6715572,0.58175594,0.48805028,0.39824903,0.3435874,0.28892577,0.23426414,0.1796025,0.12494087,0.10932326,0.093705654,0.078088045,0.06637484,0.05075723,0.058566034,0.07027924,0.078088045,0.08980125,0.10151446,0.22645533,0.3513962,0.47633708,0.60127795,0.7262188,0.58175594,0.43338865,0.28892577,0.14446288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3631094,0.7301232,1.0932326,1.4602464,1.8233559,1.6906061,1.5539521,1.4212024,1.2845483,1.1517987,1.3001659,1.4485333,1.6008049,1.7491722,1.901444,2.1239948,2.35045,2.5769055,2.7994564,3.0259118,2.803361,2.5847144,2.366068,2.1435168,1.9248703,2.4480603,2.9751544,3.4983444,4.025439,4.548629,3.978586,3.408543,2.8385005,2.2684577,1.698415,1.6242313,1.5500476,1.475864,1.4016805,1.3235924,1.3665408,1.4055848,1.4446288,1.4836729,1.5266213,1.4797685,1.43682,1.3899672,1.3431144,1.3001659,1.4992905,1.698415,1.901444,2.1005683,2.2996929,2.4090161,2.514435,2.6237583,2.7291772,2.8385005,2.5300527,2.2216048,1.9131571,1.6086137,1.3001659,1.1791295,1.0541886,0.93315214,0.80821127,0.6871748,1.0541886,1.4212024,1.7882162,2.1591344,2.5261483,2.8463092,3.1664703,3.4866312,3.8067923,4.126953,5.056201,5.985449,6.914696,7.843944,8.773191,9.187058,9.600925,10.010887,10.424754,10.838621,10.768341,10.698062,10.627783,10.557504,10.487225,9.878138,9.272955,8.663869,8.058686,7.4495993,7.195813,6.9381227,6.6843367,6.4305506,6.1767645,6.2353306,6.2938967,6.356367,6.4149327,6.473499,5.7121406,4.950782,4.185519,3.4241607,2.6628022,2.174752,1.6867018,1.1986516,0.7106012,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.12884527,0.19912452,0.26549935,0.3318742,0.39824903,0.95267415,1.5031948,2.05762,2.6081407,3.1625657,2.6940374,2.2294137,1.7608855,1.2923572,0.8238289,0.7418364,0.659844,0.57785153,0.4958591,0.41386664,0.3318742,0.24597734,0.1639849,0.08199245,0.0,0.078088045,0.15617609,0.23426414,0.30844778,0.38653582,0.3474918,0.30844778,0.26940376,0.22645533,0.18741131,0.24597734,0.30063897,0.359205,0.41777104,0.47633708,4.5095844,8.546737,12.579984,16.613232,20.650383,19.791414,18.928543,18.069574,17.210606,16.351637,14.899199,13.450665,11.998228,10.549695,9.101162,10.315431,11.5297,12.743969,13.958238,15.176412,17.819693,20.466877,23.110157,25.753437,28.400621,27.444044,26.49137,25.53479,24.578213,23.625538,22.801708,21.973976,21.150146,20.326319,19.498585,19.4244,19.346313,19.268225,19.190138,19.11205,16.945107,14.778163,12.611219,10.444276,8.273428,7.141152,6.0049706,4.8687897,3.736513,2.6003318,3.1391394,3.6818514,4.220659,4.759466,5.298274,5.5091114,5.7199492,5.930787,6.141625,6.348558,5.8566036,5.364649,4.872694,4.380739,3.8887846,4.1464753,4.4041657,4.661856,4.9156423,5.173333,5.481781,5.786324,6.0908675,6.395411,6.699954,6.9068875,7.113821,7.320754,7.531592,7.7385254,13.403813,19.069101,24.734388,30.395771,36.061058,30.360632,24.6563,18.955873,13.251541,7.551114,7.7111945,7.871275,8.031356,8.191436,8.351517,6.8366084,5.3256044,3.8106966,2.2996929,0.78868926,0.6442264,0.5036679,0.359205,0.21864653,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.078088045,0.08589685,0.08980125,0.093705654,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7340276,1.4719596,2.2059872,2.9400148,3.6740425,2.9400148,2.2059872,1.4680552,0.7340276,0.0,0.64032197,1.2806439,1.9209659,2.5612879,3.2016098,2.631567,2.0615244,1.4914817,0.92143893,0.3513962,1.1283722,1.9053483,2.6823244,3.4593005,4.2362766,3.5608149,2.8892577,2.2137961,1.5383345,0.8628729,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.59346914,1.038571,1.4836729,1.9287747,2.3738766,3.2484627,4.123049,5.001539,5.8761253,6.7507114,5.8292727,4.911738,3.9902992,3.06886,2.1513257,2.0029583,1.8545911,1.7062237,1.5617609,1.4133936,1.3001659,1.1869383,1.0737107,0.96438736,0.8511597,0.6949836,0.5388075,0.38653582,0.23035973,0.07418364,0.3513962,0.62860876,0.9058213,1.1869383,1.4641509,1.2689307,1.0737107,0.8784905,0.6832704,0.48805028,0.42948425,0.3709182,0.31625658,0.25769055,0.19912452,0.1835069,0.1717937,0.15617609,0.14055848,0.12494087,0.10541886,0.08589685,0.06637484,0.046852827,0.023426414,0.031235218,0.03513962,0.039044023,0.046852827,0.05075723,0.113227665,0.1756981,0.23816854,0.30063897,0.3631094,0.28892577,0.21864653,0.14446288,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1835069,0.3631094,0.5466163,0.7301232,0.9136301,0.8433509,0.77697605,0.7106012,0.6442264,0.57394713,0.6754616,0.77307165,0.8745861,0.97610056,1.0737107,1.2494087,1.4251068,1.6008049,1.7765031,1.9482968,1.9131571,1.8819219,1.8467822,1.8116426,1.7765031,2.5378613,3.2992198,4.0644827,4.825841,5.5871997,4.853172,4.1191444,3.3812122,2.6471848,1.9131571,1.8116426,1.7140326,1.6125181,1.5110037,1.4133936,1.4329157,1.4524376,1.4719596,1.4914817,1.5110037,1.3899672,1.2689307,1.1439898,1.0229534,0.9019169,1.0502841,1.1986516,1.3509232,1.4992905,1.6515622,1.9209659,2.194274,2.4675822,2.7408905,3.0141985,2.6276627,2.241127,1.8584955,1.4719596,1.0893283,0.96829176,0.8511597,0.7340276,0.61689556,0.4997635,0.7262188,0.95657855,1.183034,1.4094892,1.6359446,1.9365835,2.233318,2.5300527,2.8267872,3.1235218,3.9278288,4.728231,5.532538,6.336845,7.137247,7.523783,7.914223,8.300759,8.687295,9.073831,8.929368,8.781001,8.632633,8.484266,8.335898,8.050878,7.7658563,7.480835,7.195813,6.910792,7.0708723,7.230953,7.3910336,7.551114,7.7111945,7.8556576,7.996216,8.140678,8.281238,8.4257,7.4495993,6.473499,5.5013027,4.5252023,3.5491016,2.900971,2.2489357,1.6008049,0.94876975,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.08980125,0.11713207,0.14446288,0.1717937,0.19912452,0.5192855,0.8394465,1.1596074,1.4797685,1.7999294,1.53443,1.2689307,1.0034313,0.7418364,0.47633708,0.45291066,0.42948425,0.40605783,0.38653582,0.3631094,0.28892577,0.21864653,0.14446288,0.07418364,0.0,0.093705654,0.19131571,0.28502136,0.37872702,0.47633708,0.42948425,0.38653582,0.339683,0.29673457,0.24988174,0.24597734,0.24597734,0.24207294,0.23816854,0.23816854,3.330455,6.422742,9.515028,12.607315,15.699601,16.13299,16.56638,16.995863,17.429253,17.86264,15.375536,12.888432,10.401327,7.914223,5.423215,7.656533,9.889851,12.123169,14.356487,16.585901,17.671324,18.756748,19.842173,20.927597,22.01302,22.78609,23.559164,24.328331,25.101402,25.874474,24.539167,23.199959,21.860748,20.525442,19.186234,18.592764,17.999294,17.40192,16.808453,16.211079,14.9109125,13.606842,12.306676,11.002605,9.698535,8.156297,6.6140575,5.0718184,3.5295796,1.9873407,2.1200905,2.25284,2.3855898,2.5183394,2.6510892,2.7565079,2.8580225,2.9634414,3.06886,3.174279,2.97125,2.7682211,2.5690966,2.366068,2.1630387,2.7213683,3.2836022,3.8419318,4.4041657,4.9624953,5.376362,5.794133,6.2079997,6.621866,7.0357327,6.785851,6.532065,6.278279,6.028397,5.774611,13.571702,21.36489,29.16198,36.955166,44.748356,37.64234,30.53633,23.426414,16.320402,9.21439,9.593117,9.971844,10.354475,10.733202,11.111929,9.101162,7.08649,5.0757227,3.0610514,1.0502841,0.8589685,0.6715572,0.48024148,0.28892577,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.10151446,0.10541886,0.10932326,0.10932326,0.113227665,0.113227665,0.113227665,0.113227665,0.113227665,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3670138,0.7340276,1.1010414,1.4680552,1.8389735,1.4680552,1.1010414,0.7340276,0.3670138,0.0,0.32016098,0.64032197,0.96048295,1.2806439,1.6008049,1.3509232,1.1049459,0.8589685,0.60908675,0.3631094,1.3079748,2.25284,3.1977055,4.142571,5.087436,4.298747,3.513962,2.7252727,1.9365835,1.1517987,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23816854,0.47633708,0.7106012,0.94876975,1.1869383,2.639376,4.087909,5.5364423,6.98888,8.437413,7.223144,6.012779,4.7985106,3.5881457,2.3738766,2.2255092,2.0732377,1.9248703,1.7765031,1.6242313,1.5110037,1.4016805,1.2884527,1.175225,1.0619974,0.8628729,0.6637484,0.46071947,0.26159495,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.37482262,0.4997635,0.62470436,0.74964523,0.8745861,1.0268579,1.175225,1.3235924,1.475864,1.6242313,2.6237583,3.6232853,4.6267166,5.6262436,6.6257706,5.7238536,4.825841,3.9239242,3.0259118,2.1239948,1.999054,1.8741131,1.7491722,1.6242313,1.4992905,1.4992905,1.4992905,1.4992905,1.4992905,1.4992905,1.3001659,1.1010414,0.9019169,0.698888,0.4997635,0.60127795,0.698888,0.80040246,0.9019169,0.999527,1.43682,1.8741131,2.3114061,2.7486992,3.1859922,2.7252727,2.260649,1.7999294,1.33921,0.8745861,0.76135844,0.6481308,0.5388075,0.42557985,0.31235218,0.39824903,0.48805028,0.57394713,0.6637484,0.74964523,1.0268579,1.3001659,1.5734742,1.8506867,2.1239948,2.7994564,3.474918,4.1503797,4.825841,5.5013027,5.8644123,6.223617,6.5867267,6.949836,7.3129454,7.08649,6.8639393,6.6374836,6.4110284,6.1884775,6.223617,6.262661,6.3017054,6.336845,6.375889,6.949836,7.523783,8.101635,8.675582,9.249529,9.475985,9.698535,9.924991,10.151445,10.373997,9.187058,8.00012,6.813182,5.6262436,4.4393053,3.6232853,2.8111696,1.999054,1.1869383,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.37482262,0.31235218,0.24988174,0.18741131,0.12494087,0.1639849,0.19912452,0.23816854,0.27330816,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.113227665,0.22645533,0.3357786,0.44900626,0.5622339,0.5114767,0.46071947,0.41386664,0.3631094,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,2.1513257,4.298747,6.4500723,8.601398,10.748819,12.4745655,14.200311,15.926057,17.651802,19.373644,15.847969,12.326198,8.800523,5.2748475,1.7491722,5.001539,8.250002,11.498465,14.750832,17.999294,17.526861,17.050524,16.574188,16.101755,15.625418,18.124235,20.623053,23.125774,25.624592,28.12341,26.276627,24.425941,22.575254,20.724567,18.87388,17.761126,16.64837,15.535617,14.426766,13.314012,12.8767185,12.439425,11.998228,11.560935,11.123642,9.175345,7.223144,5.2748475,3.3265507,1.3743496,1.1010414,0.8238289,0.5505207,0.27330816,0.0,0.0,0.0,0.0,0.0,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,1.3001659,2.1630387,3.0259118,3.8887846,4.7516575,5.2748475,5.7980375,6.3251314,6.8483214,7.375416,6.66091,5.950309,5.2358036,4.5252023,3.8106966,13.739592,23.660677,33.589573,43.514565,53.43565,44.924053,36.412457,27.900858,19.389261,10.87376,11.475039,12.076316,12.67369,13.274967,13.8762455,11.361811,8.85128,6.336845,3.8263142,1.3118792,1.0737107,0.8394465,0.60127795,0.3631094,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,1.4875772,2.6003318,3.7130866,4.825841,5.938596,5.036679,4.138666,3.2367494,2.338737,1.43682,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19131571,0.37872702,0.5700427,0.76135844,0.94876975,2.194274,3.4397783,4.6852827,5.930787,7.1762915,6.168956,5.165524,4.1581883,3.154757,2.1513257,2.1903696,2.2294137,2.2684577,2.3114061,2.35045,2.2137961,2.0732377,1.9365835,1.7999294,1.6632754,1.3782539,1.097137,0.8160201,0.5309987,0.24988174,0.20302892,0.15617609,0.10932326,0.058566034,0.011713207,0.031235218,0.046852827,0.06637484,0.08199245,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.30063897,0.39824903,0.4997635,0.60127795,0.698888,0.8199245,0.94096094,1.0580931,1.1791295,1.3001659,2.1005683,2.900971,3.7013733,4.5017757,5.298274,4.579864,3.8614538,3.1391394,2.4207294,1.698415,1.6008049,1.5031948,1.4055848,1.3118792,1.2142692,1.2337911,1.2572175,1.2806439,1.3040704,1.3235924,1.1986516,1.0698062,0.94096094,0.8160201,0.6871748,0.79259366,0.8980125,1.0034313,1.1088502,1.2142692,1.7882162,2.3621633,2.9361105,3.513962,4.087909,3.5998588,3.1118085,2.6237583,2.135708,1.6515622,1.3782539,1.1049459,0.8316377,0.5583295,0.28892577,0.3513962,0.41777104,0.48414588,0.5466163,0.61299115,0.8902037,1.1674163,1.4446288,1.7218413,1.999054,2.6003318,3.2016098,3.7989833,4.4002614,5.001539,5.3724575,5.743376,6.1181984,6.4891167,6.8639393,6.754616,6.649197,6.5398736,6.4305506,6.3251314,6.1767645,6.0244927,5.8761253,5.7238536,5.575486,6.0635366,6.5554914,7.043542,7.535496,8.023546,8.226576,8.4257,8.624825,8.823949,9.023073,8.086017,7.1489606,6.211904,5.2748475,4.337791,3.5451972,2.7526035,1.9600099,1.1674163,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.12103647,0.093705654,0.06637484,0.039044023,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.019522011,0.015617609,0.015617609,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.10151446,0.1756981,0.24988174,0.3240654,0.39824903,0.3240654,0.24988174,0.1756981,0.10151446,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.3240654,0.26940376,0.21864653,0.1639849,0.113227665,0.14055848,0.1678893,0.19522011,0.22255093,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.10151446,0.20693332,0.30844778,0.40996224,0.5114767,0.46071947,0.40605783,0.3553006,0.30063897,0.24988174,0.23816854,0.23035973,0.21864653,0.21083772,0.19912452,2.1435168,4.084005,6.028397,7.968885,9.913278,11.04165,12.173926,13.302299,14.430671,15.562947,13.688834,11.810817,9.936704,8.062591,6.1884775,9.089449,11.986515,14.8874855,17.788456,20.689428,20.958832,21.228235,21.497639,21.767042,22.036446,23.188246,24.33614,25.487938,26.635832,27.78763,26.549934,25.31224,24.074545,22.83685,21.599154,19.838268,18.081287,16.320402,14.559516,12.798631,12.517513,12.236397,11.951375,11.6702585,11.389141,9.331521,7.277806,5.22409,3.1664703,1.1127546,0.8941081,0.679366,0.46071947,0.24207294,0.023426414,0.03513962,0.046852827,0.05466163,0.06637484,0.07418364,0.22255093,0.3709182,0.5192855,0.6637484,0.81211567,1.43682,2.0615244,2.6862288,3.310933,3.9356375,4.369026,4.7985106,5.2279944,5.657479,6.086963,5.481781,4.872694,4.263607,3.6584249,3.049338,10.990892,18.928543,26.870096,34.81165,42.749302,37.185528,31.625658,26.061886,20.498112,14.938243,14.789876,14.641508,14.493141,14.348679,14.200311,11.916236,9.636065,7.3519893,5.0718184,2.787743,2.366068,1.9482968,1.5266213,1.1088502,0.6871748,0.5583295,0.43338865,0.30454338,0.1756981,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.13665408,0.13274968,0.12884527,0.12884527,0.12494087,0.12884527,0.12884527,0.13274968,0.13665408,0.13665408,0.113227665,0.08589685,0.062470436,0.039044023,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06637484,0.12884527,0.19522011,0.26159495,0.3240654,1.2806439,2.241127,3.1977055,4.154284,5.1108627,4.3260775,3.5373883,2.7486992,1.9639144,1.175225,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14055848,0.28502136,0.42557985,0.5700427,0.7106012,1.7530766,2.7916477,3.8341231,4.872694,5.911265,5.114767,4.318269,3.521771,2.7213683,1.9248703,2.15523,2.3855898,2.6159496,2.8463092,3.076669,2.912684,2.7486992,2.5886188,2.4246337,2.260649,1.8975395,1.53443,1.1674163,0.80430686,0.43729305,0.3553006,0.27330816,0.19131571,0.10932326,0.023426414,0.03513962,0.046852827,0.05466163,0.06637484,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.22645533,0.30063897,0.37482262,0.44900626,0.5231899,0.61689556,0.7066968,0.79649806,0.8862993,0.97610056,1.5734742,2.174752,2.77603,3.3734035,3.9746814,3.435874,2.893162,2.3543546,1.815547,1.2767396,1.2064602,1.1361811,1.0659018,0.9956226,0.92534333,0.96829176,1.0151446,1.0580931,1.1049459,1.1517987,1.0932326,1.038571,0.98390937,0.92924774,0.8745861,0.98390937,1.0932326,1.2064602,1.3157835,1.4251068,2.135708,2.8502135,3.5608149,4.2753205,4.985922,4.474445,3.9629683,3.4514916,2.9361105,2.4246337,1.9912452,1.5617609,1.1283722,0.6949836,0.26159495,0.30454338,0.3474918,0.39044023,0.43338865,0.47633708,0.75354964,1.0346665,1.3157835,1.5969005,1.8741131,2.4012074,2.9243972,3.4514916,3.9746814,4.5017757,4.884407,5.263134,5.645766,6.028397,6.4110284,6.422742,6.4305506,6.4422636,6.453977,6.461786,6.126007,5.786324,5.4505453,5.1108627,4.775084,5.181142,5.5832953,5.989353,6.395411,6.801469,6.9732623,7.1489606,7.3246584,7.5003567,7.676055,6.98888,6.3017054,5.610626,4.9234514,4.2362766,3.4632049,2.6940374,1.9209659,1.1478943,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.14446288,0.113227665,0.08589685,0.05466163,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.046852827,0.039044023,0.03513962,0.031235218,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.19912452,0.3513962,0.4997635,0.6481308,0.80040246,0.6481308,0.4997635,0.3513962,0.19912452,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.26940376,0.22645533,0.1835069,0.14055848,0.10151446,0.11713207,0.13665408,0.15227169,0.1717937,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.093705654,0.1835069,0.27721256,0.3709182,0.46071947,0.40605783,0.3513962,0.29673457,0.24207294,0.18741131,0.23035973,0.27330816,0.31625658,0.359205,0.39824903,2.135708,3.8692627,5.606722,7.3402762,9.073831,9.608734,10.143637,10.67854,11.213444,11.748346,11.525795,11.29934,11.076789,10.850334,10.6238785,13.173453,15.723028,18.276506,20.826082,23.375656,24.3908,25.405945,26.42109,27.436235,28.45138,28.24835,28.049225,27.850101,27.650976,27.451853,26.823244,26.19854,25.573835,24.949131,24.324427,21.919313,19.510298,17.101282,14.69617,12.287154,12.158309,12.033368,11.904523,11.775677,11.650736,9.491602,7.328563,5.169429,3.0102942,0.8511597,0.6910792,0.5309987,0.3709182,0.21083772,0.05075723,0.07027924,0.08980125,0.10932326,0.12884527,0.14836729,0.359205,0.5661383,0.77307165,0.98000497,1.1869383,1.5734742,1.9639144,2.35045,2.736986,3.1235218,3.4593005,3.795079,4.1308575,4.466636,4.7985106,4.298747,3.795079,3.2914112,2.7916477,2.2879796,8.242193,14.196406,20.154524,26.108738,32.06295,29.450907,26.838861,24.226816,21.610867,18.998821,18.104713,17.210606,16.316498,15.418485,14.524376,12.470661,10.42085,8.367134,6.3134184,4.263607,3.6584249,3.057147,2.455869,1.8506867,1.2494087,1.0073358,0.76526284,0.5231899,0.28111696,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.14446288,0.14055848,0.13665408,0.12884527,0.12494087,0.12884527,0.13665408,0.14055848,0.14446288,0.14836729,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05466163,0.10932326,0.1639849,0.21864653,0.27330816,1.077615,1.8819219,2.6823244,3.4866312,4.2870336,3.611572,2.9361105,2.260649,1.5890918,0.9136301,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.093705654,0.19131571,0.28502136,0.37872702,0.47633708,1.3118792,2.1435168,2.979059,3.814601,4.650143,4.0605783,3.4710135,2.8814487,2.2918842,1.698415,2.1200905,2.541766,2.959537,3.3812122,3.7989833,3.611572,3.4241607,3.2367494,3.049338,2.8619268,2.416825,1.9678187,1.5188124,1.0737107,0.62470436,0.5075723,0.39044023,0.27330816,0.15617609,0.039044023,0.039044023,0.042948425,0.046852827,0.046852827,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.14836729,0.19912452,0.24988174,0.30063897,0.3513962,0.40996224,0.46852827,0.5309987,0.58956474,0.6481308,1.0502841,1.4485333,1.8506867,2.2489357,2.6510892,2.2918842,1.9287747,1.5695697,1.2103647,0.8511597,0.80821127,0.76526284,0.7223144,0.679366,0.63641757,0.7066968,0.77307165,0.8394465,0.9058213,0.97610056,0.9917182,1.0112402,1.0268579,1.0463798,1.0619974,1.1791295,1.2923572,1.4055848,1.5227169,1.6359446,2.4871042,3.338264,4.1894236,5.036679,5.8878384,5.349031,4.814128,4.2753205,3.736513,3.2016098,2.6081407,2.0146716,1.4212024,0.8316377,0.23816854,0.25769055,0.27721256,0.29673457,0.31625658,0.3357786,0.62079996,0.9019169,1.1869383,1.4680552,1.7491722,2.1981785,2.6510892,3.1000953,3.5491016,3.998108,4.3924527,4.786797,5.1772375,5.571582,5.9620223,6.0908675,6.2158084,6.3446536,6.473499,6.5984397,6.0752497,5.548156,5.024966,4.5017757,3.9746814,4.2948427,4.6150036,4.9351645,5.2553253,5.575486,5.7238536,5.8761253,6.0244927,6.1767645,6.3251314,5.8878384,5.4505453,5.0132523,4.575959,4.138666,3.3851168,2.631567,1.8819219,1.1283722,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.1678893,0.13665408,0.10151446,0.07027924,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.30063897,0.5231899,0.74964523,0.97610056,1.1986516,0.97610056,0.74964523,0.5231899,0.30063897,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.21864653,0.1835069,0.15227169,0.12103647,0.08589685,0.093705654,0.10151446,0.10932326,0.11713207,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.08199245,0.1639849,0.24597734,0.3318742,0.41386664,0.3553006,0.29673457,0.23816854,0.1835069,0.12494087,0.21864653,0.31625658,0.40996224,0.5036679,0.60127795,2.1278992,3.6545205,5.181142,6.7116675,8.238289,8.175818,8.117252,8.058686,7.996216,7.9376497,9.362757,10.787864,12.212971,13.638077,15.063184,17.261362,19.463446,21.661623,23.863707,26.061886,27.822771,29.583656,31.340637,33.10152,34.862408,33.31236,31.762312,30.212265,28.662216,27.11217,27.100456,27.088743,27.073126,27.061413,27.049698,23.996456,20.93931,17.886066,14.828919,11.775677,11.803008,11.8303385,11.85767,11.885,11.912332,9.647778,7.3832245,5.1186714,2.854118,0.58566034,0.48414588,0.38263142,0.28111696,0.1756981,0.07418364,0.10541886,0.13665408,0.1639849,0.19522011,0.22645533,0.49195468,0.76135844,1.0268579,1.2962615,1.5617609,1.7140326,1.8623998,2.0107672,2.1630387,2.3114061,2.5534792,2.7916477,3.0337205,3.2718892,3.513962,3.1157131,2.717464,2.3192148,1.9209659,1.5266213,5.493494,9.464272,13.435048,17.405825,21.376602,21.712381,22.048159,22.387842,22.723621,23.063305,21.41955,19.775797,18.135948,16.492195,14.848442,13.028991,11.205634,9.382278,7.558923,5.735567,4.950782,4.165997,3.3812122,2.5964274,1.8116426,1.456342,1.097137,0.7418364,0.38263142,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.031235218,0.06637484,0.09761006,0.12884527,0.1639849,0.15617609,0.14836729,0.14055848,0.13274968,0.12494087,0.13274968,0.14055848,0.14836729,0.15617609,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.08980125,0.13665408,0.1796025,0.22645533,0.8706817,1.5188124,2.1669433,2.815074,3.4632049,2.900971,2.338737,1.7765031,1.2142692,0.6481308,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.093705654,0.14055848,0.19131571,0.23816854,0.8667773,1.4992905,2.1278992,2.7565079,3.3890212,3.0063896,2.6237583,2.241127,1.8584955,1.475864,2.084951,2.6940374,3.3031244,3.9161155,4.5252023,4.3143644,4.0996222,3.8887846,3.6740425,3.4632049,2.9322062,2.4012074,1.8741131,1.3431144,0.81211567,0.659844,0.5075723,0.3553006,0.20302892,0.05075723,0.046852827,0.039044023,0.03513962,0.031235218,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.1756981,0.20693332,0.23426414,0.26549935,0.29673457,0.3240654,0.5231899,0.7262188,0.92534333,1.1244678,1.3235924,1.1439898,0.96438736,0.78478485,0.60518235,0.42557985,0.40996224,0.39434463,0.37872702,0.3631094,0.3513962,0.44119745,0.5309987,0.62079996,0.7106012,0.80040246,0.8902037,0.98000497,1.0698062,1.1596074,1.2494087,1.3704453,1.4914817,1.6086137,1.7296503,1.8506867,2.8385005,3.8263142,4.814128,5.801942,6.785851,6.223617,5.661383,5.099149,4.5369153,3.9746814,3.2211318,2.4714866,1.717937,0.96438736,0.21083772,0.21083772,0.20693332,0.20693332,0.20302892,0.19912452,0.48414588,0.76916724,1.0541886,1.33921,1.6242313,1.999054,2.3738766,2.7486992,3.1235218,3.4983444,3.9044023,4.3065557,4.7087092,5.1108627,5.5130157,5.758993,6.001066,6.2470436,6.493021,6.7389984,6.0244927,5.3138914,4.5993857,3.8887846,3.174279,3.408543,3.6467118,3.8809757,4.11524,4.349504,4.474445,4.5993857,4.7243266,4.8492675,4.9742084,4.786797,4.5993857,4.4119744,4.224563,4.037152,3.3031244,2.5730011,1.8389735,1.1088502,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.046852827,0.08980125,0.13665408,0.1796025,0.22645533,0.19131571,0.15617609,0.12103647,0.08589685,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.39824903,0.698888,0.999527,1.3001659,1.6008049,1.3001659,0.999527,0.698888,0.39824903,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.1639849,0.14055848,0.12103647,0.09761006,0.07418364,0.07418364,0.07027924,0.06637484,0.06637484,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.07418364,0.14446288,0.21864653,0.28892577,0.3631094,0.30063897,0.24207294,0.1835069,0.12103647,0.062470436,0.21083772,0.359205,0.5036679,0.6520352,0.80040246,2.1200905,3.4397783,4.759466,6.0791545,7.3988423,6.746807,6.0908675,5.434928,4.7789884,4.123049,7.1997175,10.276386,13.349152,16.42582,19.498585,21.349272,23.199959,25.050644,26.90133,28.748114,31.25474,33.761368,36.264088,38.770714,41.273438,38.37637,35.4754,32.57443,29.673458,26.77639,27.373764,27.975042,28.57632,29.173695,29.774971,26.073599,22.36832,18.666946,14.965574,11.2642,11.443803,11.62731,11.810817,11.994324,12.173926,9.803954,7.433982,5.0640097,2.6940374,0.3240654,0.28111696,0.23426414,0.19131571,0.14446288,0.10151446,0.14055848,0.1796025,0.21864653,0.26159495,0.30063897,0.62860876,0.95657855,1.2806439,1.6086137,1.9365835,1.8506867,1.7608855,1.6749885,1.5890918,1.4992905,1.6437533,1.7882162,1.9365835,2.0810463,2.2255092,1.9326792,1.639849,1.3470187,1.0541886,0.76135844,2.7486992,4.732136,6.715572,8.702912,10.686349,13.973856,17.261362,20.548868,23.836376,27.123882,24.734388,22.344894,19.9554,17.565907,15.176412,13.583415,11.990419,10.397423,8.804427,7.211431,6.2431393,5.278752,4.31046,3.3421683,2.3738766,1.901444,1.4290112,0.95657855,0.48414588,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.1639849,0.15617609,0.14446288,0.13665408,0.12494087,0.13665408,0.14446288,0.15617609,0.1639849,0.1756981,0.14836729,0.12494087,0.10151446,0.07418364,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.6676528,1.1596074,1.6515622,2.1435168,2.639376,2.1864653,1.737459,1.2884527,0.8394465,0.38653582,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.42557985,0.8511597,1.2767396,1.698415,2.1239948,1.9482968,1.7765031,1.6008049,1.4251068,1.2494087,2.0498111,2.8502135,3.6506162,4.4510183,5.251421,5.0132523,4.775084,4.5369153,4.298747,4.0605783,3.4514916,2.8385005,2.2255092,1.6125181,0.999527,0.81211567,0.62470436,0.43729305,0.24988174,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.1756981,0.28892577,0.39824903,0.5114767,0.62470436,0.78868926,0.94876975,1.1127546,1.2767396,1.43682,1.5617609,1.6867018,1.8116426,1.9365835,2.0615244,3.1859922,4.3143644,5.4388323,6.5633,7.687768,7.098203,6.5125427,5.9268827,5.337318,4.7516575,3.8380275,2.9243972,2.0107672,1.1010414,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.3513962,0.63641757,0.92534333,1.2142692,1.4992905,1.7999294,2.1005683,2.4012074,2.7018464,2.998581,3.4124475,3.8263142,4.2362766,4.650143,5.0640097,5.423215,5.786324,6.1494336,6.5125427,6.8756523,5.9737353,5.0757227,4.173806,3.2757936,2.3738766,2.5261483,2.6745155,2.8267872,2.9751544,3.1235218,3.2250361,3.3265507,3.4241607,3.5256753,3.6232853,3.6857557,3.7482262,3.8106966,3.873167,3.9356375,3.2250361,2.514435,1.7999294,1.0893283,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.4997635,0.8745861,1.2494087,1.6242313,1.999054,1.6242313,1.2494087,0.8745861,0.4997635,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.19912452,0.39824903,0.60127795,0.80040246,0.999527,2.1122816,3.2250361,4.337791,5.4505453,6.5633,5.3138914,4.0644827,2.8111696,1.5617609,0.31235218,5.036679,9.761005,14.489237,19.213564,23.937891,25.437181,26.936472,28.435762,29.938957,31.438248,34.68671,37.939075,41.18754,44.436,47.68837,43.436474,39.188484,34.936592,30.688602,26.436708,27.650976,28.861341,30.075611,31.285975,32.500244,28.15074,23.801235,19.451733,15.098324,10.748819,11.088503,11.424281,11.763964,12.099743,12.439425,9.964035,7.4886436,5.0132523,2.5378613,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.1756981,0.22645533,0.27330816,0.3240654,0.37482262,0.76135844,1.1517987,1.5383345,1.9248703,2.3114061,1.9873407,1.6632754,1.33921,1.0112402,0.6871748,0.737932,0.78868926,0.8394465,0.8862993,0.93705654,0.74964523,0.5622339,0.37482262,0.18741131,0.0,0.0,0.0,0.0,0.0,0.0,6.239235,12.4745655,18.7138,24.949131,31.188366,28.049225,24.91399,21.77485,18.635712,15.500477,14.13784,12.775204,11.412568,10.049932,8.687295,7.535496,6.387602,5.2358036,4.087909,2.9361105,2.35045,1.7608855,1.175225,0.58566034,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.46071947,0.80040246,1.1361811,1.475864,1.8116426,1.475864,1.1361811,0.80040246,0.46071947,0.12494087,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.339683,0.679366,1.0190489,1.358732,1.698415,1.5734742,1.4446288,1.3157835,1.1908426,1.0619974,1.6906061,2.3192148,2.9439192,3.5725281,4.2011366,4.009821,3.8185053,3.631094,3.4397783,3.2484627,2.7604125,2.2684577,1.7804074,1.2884527,0.80040246,0.6481308,0.4997635,0.3513962,0.19912452,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.14055848,0.23035973,0.32016098,0.40996224,0.4997635,0.64032197,0.78088045,0.92143893,1.0580931,1.1986516,1.397776,1.5969005,1.7921207,1.9912452,2.1864653,3.076669,3.9668727,4.8570766,5.74728,6.6374836,6.1455293,5.6535745,5.1616197,4.6657605,4.173806,3.408543,2.639376,1.8741131,1.1049459,0.3357786,0.28892577,0.23816854,0.18741131,0.13665408,0.08589685,0.3240654,0.5622339,0.80040246,1.038571,1.2767396,1.5305257,1.7843118,2.0380979,2.2957885,2.5495746,2.8619268,3.174279,3.4866312,3.7989833,4.1113358,4.6540475,5.196759,5.7394714,6.282183,6.824895,6.114294,5.3997884,4.689187,3.9746814,3.2640803,3.279698,3.2992198,3.3148375,3.3343596,3.349977,3.3616903,3.3734035,3.3890212,3.4007344,3.4124475,3.435874,3.4632049,3.4866312,3.513962,3.5373883,2.900971,2.2684577,1.6320401,0.9956226,0.3631094,0.28892577,0.21864653,0.14446288,0.07418364,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.29673457,0.39044023,0.48414588,0.58175594,0.6754616,0.5466163,0.41386664,0.28502136,0.15617609,0.023426414,0.031235218,0.039044023,0.046852827,0.05466163,0.062470436,0.07027924,0.078088045,0.08589685,0.093705654,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.113227665,0.12494087,0.13665408,0.14836729,0.1639849,0.18741131,0.21083772,0.23816854,0.26159495,0.28892577,0.30844778,0.3318742,0.3553006,0.37872702,0.39824903,0.3709182,0.339683,0.30844778,0.28111696,0.24988174,0.22255093,0.19522011,0.1678893,0.14055848,0.113227665,0.40996224,0.7066968,1.0034313,1.3040704,1.6008049,1.3001659,0.999527,0.698888,0.39824903,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.10151446,0.14055848,0.1835069,0.22255093,0.26159495,0.21083772,0.15617609,0.10541886,0.05075723,0.0,0.58175594,1.1635119,1.7491722,2.330928,2.912684,3.416352,3.9239242,4.4275923,4.93126,5.4388323,4.40807,3.3812122,2.3543546,1.3274968,0.30063897,4.9546866,9.60483,14.258877,18.90902,23.563068,24.504028,25.448895,26.389854,27.330816,28.27568,31.426535,34.58129,37.732143,40.8869,44.037754,40.051357,36.061058,32.074665,28.08827,24.101875,27.881336,31.660797,35.440258,39.21972,42.999184,40.363712,37.724335,35.088863,32.449486,29.814016,27.088743,24.367374,21.646006,18.920732,16.199366,13.228115,10.260769,7.289519,4.318269,1.3509232,1.2142692,1.0815194,0.94486535,0.80821127,0.6754616,0.60518235,0.5349031,0.46462387,0.39434463,0.3240654,0.7262188,1.1283722,1.53443,1.9365835,2.338737,2.0537157,1.7725986,1.4914817,1.2064602,0.92534333,0.94876975,0.97610056,0.999527,1.0268579,1.0502841,0.9917182,0.92924774,0.8706817,0.80821127,0.74964523,0.6871748,0.62470436,0.5622339,0.4997635,0.43729305,5.3412223,10.241247,15.145176,20.049105,24.949131,22.4386,19.92807,17.421442,14.9109125,12.400381,11.311053,10.221725,9.128492,8.039165,6.949836,6.028397,5.1108627,4.1894236,3.2718892,2.35045,1.8780174,1.4094892,0.94096094,0.46852827,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.05466163,0.09761006,0.14055848,0.1835069,0.22645533,0.20693332,0.19131571,0.1717937,0.15617609,0.13665408,0.14055848,0.14836729,0.15227169,0.15617609,0.1639849,0.14055848,0.12103647,0.10151446,0.08199245,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.44900626,0.74574083,1.0424755,1.33921,1.6359446,1.3314011,1.0229534,0.7145056,0.40605783,0.10151446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25378615,0.5114767,0.76526284,1.0190489,1.2767396,1.1947471,1.116659,1.0346665,0.95657855,0.8745861,1.3314011,1.7843118,2.241127,2.6940374,3.1508527,3.0063896,2.8658314,2.7213683,2.5808098,2.436347,2.069333,1.7023194,1.3353056,0.96829176,0.60127795,0.48805028,0.37482262,0.26159495,0.14836729,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.10541886,0.1717937,0.23816854,0.30844778,0.37482262,0.49195468,0.60908675,0.7262188,0.8433509,0.96438736,1.2337911,1.5031948,1.7725986,2.0420024,2.3114061,2.9673457,3.6232853,4.279225,4.93126,5.5871997,5.1889505,4.7907014,4.396357,3.998108,3.5998588,2.979059,2.3543546,1.7335546,1.1088502,0.48805028,0.41386664,0.3357786,0.26159495,0.18741131,0.113227665,0.30063897,0.48805028,0.6754616,0.8628729,1.0502841,1.261122,1.4680552,1.678893,1.8897307,2.1005683,2.3114061,2.5261483,2.736986,2.951728,3.1625657,3.8848803,4.607195,5.3295093,6.0518236,6.774138,6.250948,5.7238536,5.2006636,4.6735697,4.1503797,4.0332475,3.9200199,3.8067923,3.68966,3.5764325,3.4983444,3.4241607,3.349977,3.2757936,3.2016098,3.1859922,3.174279,3.1625657,3.1508527,3.1391394,2.5808098,2.0224805,1.4641509,0.9058213,0.3513962,0.28111696,0.21083772,0.14055848,0.07027924,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.37872702,0.60518235,0.8316377,1.0580931,1.2884527,1.038571,0.79259366,0.5466163,0.29673457,0.05075723,0.06637484,0.078088045,0.093705654,0.10932326,0.12494087,0.113227665,0.10541886,0.093705654,0.08589685,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.13665408,0.1639849,0.18741131,0.21083772,0.23816854,0.26159495,0.3240654,0.38653582,0.44900626,0.5114767,0.57394713,0.62079996,0.6637484,0.7106012,0.75354964,0.80040246,0.7418364,0.679366,0.62079996,0.5583295,0.4997635,0.42167544,0.339683,0.26159495,0.1796025,0.10151446,0.32016098,0.5388075,0.76135844,0.98000497,1.1986516,0.97610056,0.74964523,0.5231899,0.30063897,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.14055848,0.16008049,0.1756981,0.19522011,0.21083772,0.1717937,0.12884527,0.08589685,0.042948425,0.0,0.96438736,1.9287747,2.893162,3.8614538,4.825841,4.7243266,4.618908,4.5173936,4.415879,4.3143644,3.506153,2.7018464,1.8975395,1.0932326,0.28892577,4.8687897,9.448653,14.028518,18.608381,23.188246,23.570877,23.957413,24.343948,24.72658,25.113115,28.166357,31.223505,34.27675,37.333893,40.38714,36.66234,32.93754,29.212738,25.487938,21.763138,28.111696,34.45635,40.80491,47.153465,53.502026,52.57668,51.651337,50.725994,49.80065,48.87531,43.092888,37.310467,31.528048,25.745628,19.96321,16.4961,13.032895,9.565785,6.1025805,2.639376,2.3543546,2.0732377,1.7882162,1.5070993,1.2259823,1.0346665,0.8433509,0.6559396,0.46462387,0.27330816,0.6910792,1.1088502,1.5266213,1.9443923,2.3621633,2.1239948,1.8819219,1.6437533,1.4016805,1.1635119,1.1635119,1.1635119,1.1635119,1.1635119,1.1635119,1.2298868,1.2962615,1.3665408,1.4329157,1.4992905,1.3743496,1.2494087,1.1244678,0.999527,0.8745861,4.4432096,8.007929,11.576552,15.145176,18.7138,16.827974,14.946052,13.06413,11.182208,9.300286,8.484266,7.6643414,6.8483214,6.028397,5.212377,4.521298,3.8341231,3.1430438,2.4519646,1.7608855,1.4094892,1.0580931,0.7066968,0.3513962,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.07418364,0.12103647,0.1678893,0.21474212,0.26159495,0.23816854,0.21864653,0.19522011,0.1717937,0.14836729,0.14836729,0.14446288,0.14055848,0.14055848,0.13665408,0.12103647,0.10932326,0.093705654,0.078088045,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.43338865,0.6910792,0.94876975,1.2064602,1.4641509,1.183034,0.9058213,0.62860876,0.3513962,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1717937,0.339683,0.5114767,0.679366,0.8511597,0.8160201,0.78478485,0.75354964,0.71841,0.6871748,0.96829176,1.2533131,1.53443,1.8194515,2.1005683,2.0068626,1.9092526,1.815547,1.7218413,1.6242313,1.3782539,1.1361811,0.8902037,0.6442264,0.39824903,0.3240654,0.24988174,0.1756981,0.10151446,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.07027924,0.113227665,0.16008049,0.20693332,0.24988174,0.3435874,0.44119745,0.5349031,0.62860876,0.7262188,1.0659018,1.4094892,1.7530766,2.096664,2.436347,2.8580225,3.2757936,3.697469,4.1191444,4.5369153,4.2362766,3.9317331,3.631094,3.3265507,3.0259118,2.5456703,2.069333,1.5929961,1.116659,0.63641757,0.5388075,0.43729305,0.3357786,0.23816854,0.13665408,0.27330816,0.41386664,0.5505207,0.6871748,0.8238289,0.9917182,1.1557031,1.319688,1.4836729,1.6515622,1.7608855,1.8741131,1.9873407,2.1005683,2.2137961,3.1157131,4.01763,4.919547,5.8214636,6.7233806,6.387602,6.0518236,5.7121406,5.376362,5.036679,4.7907014,4.5408196,4.2948427,4.0488653,3.7989833,3.638903,3.474918,3.310933,3.1508527,2.9868677,2.9361105,2.8892577,2.8385005,2.787743,2.736986,2.2567444,1.7765031,1.2962615,0.8160201,0.3357786,0.26940376,0.20302892,0.13665408,0.06637484,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.46071947,0.8199245,1.1791295,1.5383345,1.901444,1.53443,1.1713207,0.80430686,0.44119745,0.07418364,0.09761006,0.12103647,0.14055848,0.1639849,0.18741131,0.16008049,0.13274968,0.10541886,0.078088045,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.1756981,0.21083772,0.24988174,0.28892577,0.3240654,0.3631094,0.46071947,0.5622339,0.6637484,0.76135844,0.8628729,0.92924774,0.9956226,1.0659018,1.1322767,1.1986516,1.1088502,1.0190489,0.92924774,0.8394465,0.74964523,0.61689556,0.48414588,0.3513962,0.21864653,0.08589685,0.23035973,0.3709182,0.5153811,0.6559396,0.80040246,0.6481308,0.4997635,0.3513962,0.19912452,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.046852827,0.039044023,0.03513962,0.031235218,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.1835069,0.1756981,0.1717937,0.1678893,0.1639849,0.12884527,0.09761006,0.06637484,0.031235218,0.0,1.3470187,2.6940374,4.041056,5.388075,6.7389984,6.028397,5.3177958,4.607195,3.8965936,3.1859922,2.6042364,2.0224805,1.4407244,0.8589685,0.27330816,4.7828927,9.288573,13.798158,18.303837,22.813423,22.641628,22.46593,22.294136,22.122343,21.95055,24.906181,27.865719,30.821352,33.780888,36.736523,33.273315,29.814016,26.350811,22.887606,19.4244,28.342056,37.255806,46.169556,55.083305,64.00096,64.78574,65.57443,66.36313,67.15182,67.9366,59.09313,50.253563,41.41009,32.56662,23.723148,19.764084,15.80502,11.845957,7.882988,3.9239242,3.49444,3.0649557,2.6354716,2.2059872,1.7765031,1.4641509,1.1557031,0.8433509,0.5349031,0.22645533,0.6559396,1.0893283,1.5227169,1.9561055,2.3855898,2.1903696,1.9912452,1.796025,1.5969005,1.4016805,1.3743496,1.3509232,1.3235924,1.3001659,1.2767396,1.4719596,1.6632754,1.8584955,2.0537157,2.2489357,2.0615244,1.8741131,1.6867018,1.4992905,1.3118792,3.5451972,5.7785153,8.011833,10.241247,12.4745655,11.221252,9.964035,8.710721,7.453504,6.2001905,5.6535745,5.1108627,4.564246,4.0215344,3.474918,3.0141985,2.5534792,2.096664,1.6359446,1.175225,0.94096094,0.7066968,0.46852827,0.23426414,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.08980125,0.14055848,0.19522011,0.24597734,0.30063897,0.27330816,0.24597734,0.21864653,0.19131571,0.1639849,0.15227169,0.14055848,0.13274968,0.12103647,0.113227665,0.10151446,0.093705654,0.08199245,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.41777104,0.63641757,0.8511597,1.0698062,1.2884527,1.038571,0.79259366,0.5466163,0.29673457,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08589685,0.1717937,0.25378615,0.339683,0.42557985,0.44119745,0.45681506,0.46852827,0.48414588,0.4997635,0.60908675,0.71841,0.8316377,0.94096094,1.0502841,1.0034313,0.95657855,0.9058213,0.8589685,0.81211567,0.6910792,0.5661383,0.44510186,0.3240654,0.19912452,0.1639849,0.12494087,0.08589685,0.05075723,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.03513962,0.058566034,0.078088045,0.10151446,0.12494087,0.19912452,0.26940376,0.3435874,0.41386664,0.48805028,0.9019169,1.3157835,1.7335546,2.1474214,2.5612879,2.7486992,2.9322062,3.1157131,3.3031244,3.4866312,3.279698,3.0727646,2.8658314,2.6588979,2.4480603,2.1161861,1.7843118,1.4524376,1.1205635,0.78868926,0.6637484,0.5388075,0.41386664,0.28892577,0.1639849,0.24988174,0.3357786,0.42557985,0.5114767,0.60127795,0.71841,0.8394465,0.96048295,1.0815194,1.1986516,1.2142692,1.2259823,1.2376955,1.2494087,1.261122,2.3465457,3.4280653,4.5095844,5.591104,6.676528,6.524256,6.375889,6.223617,6.0752497,5.9268827,5.5442514,5.165524,4.786797,4.4041657,4.025439,3.775557,3.5256753,3.2757936,3.0259118,2.77603,2.6862288,2.6003318,2.514435,2.4246337,2.338737,1.9365835,1.53443,1.1283722,0.7262188,0.3240654,0.26159495,0.19522011,0.12884527,0.06637484,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.5427119,1.0346665,1.5266213,2.018576,2.514435,2.0302892,1.5461433,1.0659018,0.58175594,0.10151446,0.12884527,0.16008049,0.19131571,0.21864653,0.24988174,0.20693332,0.16008049,0.113227665,0.07027924,0.023426414,0.062470436,0.10151446,0.13665408,0.1756981,0.21083772,0.26159495,0.31235218,0.3631094,0.41386664,0.46071947,0.60127795,0.737932,0.8745861,1.0112402,1.1517987,1.2415999,1.3314011,1.4212024,1.5110037,1.6008049,1.4797685,1.358732,1.2415999,1.1205635,0.999527,0.8160201,0.62860876,0.44510186,0.26159495,0.07418364,0.14055848,0.20693332,0.26940376,0.3357786,0.39824903,0.3240654,0.24988174,0.1756981,0.10151446,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.019522011,0.015617609,0.015617609,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.22255093,0.19522011,0.1678893,0.14055848,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,1.7296503,3.4593005,5.1889505,6.918601,8.648251,7.3324676,6.016684,4.6969957,3.3812122,2.0615244,1.7023194,1.3431144,0.98390937,0.62079996,0.26159495,4.6969957,9.132397,13.567798,18.003199,22.4386,21.708477,20.978354,20.24823,19.518106,18.787983,21.646006,24.507933,27.365955,30.227882,33.085903,29.888199,26.68659,23.488884,20.287273,17.085665,28.572416,40.051357,51.534206,63.01705,74.4999,76.99872,79.50144,82.00026,84.49908,87.00179,75.097275,63.196655,51.292133,39.391514,27.486992,23.032068,18.577147,14.122223,9.6673,5.212377,4.6345253,4.056674,3.4788225,2.900971,2.3231194,1.893635,1.4641509,1.0346665,0.60518235,0.1756981,0.62079996,1.0698062,1.5188124,1.9639144,2.4129205,2.2567444,2.1005683,1.9482968,1.7921207,1.6359446,1.5890918,1.5383345,1.4875772,1.43682,1.3860629,1.7101282,2.0341935,2.3543546,2.67842,2.998581,2.7486992,2.4988174,2.2489357,1.999054,1.7491722,2.6471848,3.5451972,4.4432096,5.3412223,6.239235,5.610626,4.9820175,4.3534083,3.7287042,3.1000953,2.8267872,2.5534792,2.2840753,2.0107672,1.737459,1.5070993,1.2767396,1.0463798,0.8160201,0.58566034,0.46852827,0.3513962,0.23426414,0.11713207,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.10932326,0.1639849,0.22255093,0.28111696,0.3357786,0.30454338,0.27330816,0.23816854,0.20693332,0.1756981,0.15617609,0.14055848,0.12103647,0.10541886,0.08589685,0.08199245,0.078088045,0.07418364,0.06637484,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.08980125,0.13665408,0.1796025,0.22645533,0.40215343,0.58175594,0.75745404,0.93315214,1.1127546,0.8941081,0.679366,0.46071947,0.24207294,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.737932,1.2259823,1.7140326,2.1981785,2.6862288,2.639376,2.5886188,2.5378613,2.4871042,2.436347,2.3231194,2.2137961,2.1005683,1.9873407,1.8741131,1.6867018,1.4992905,1.3118792,1.1244678,0.93705654,0.78868926,0.63641757,0.48805028,0.3357786,0.18741131,0.22645533,0.26159495,0.30063897,0.3357786,0.37482262,0.44900626,0.5231899,0.60127795,0.6754616,0.74964523,0.6637484,0.57394713,0.48805028,0.39824903,0.31235218,1.5734742,2.8385005,4.0996222,5.3607445,6.6257706,6.66091,6.699954,6.7389984,6.774138,6.813182,6.3017054,5.786324,5.2748475,4.7633705,4.251894,3.912211,3.5764325,3.2367494,2.900971,2.5612879,2.436347,2.3114061,2.1864653,2.0615244,1.9365835,1.6125181,1.2884527,0.96438736,0.63641757,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.0,0.0,0.0,0.0,0.0,0.62470436,1.2494087,1.8741131,2.4988174,3.1235218,2.5261483,1.9248703,1.3235924,0.7262188,0.12494087,0.1639849,0.19912452,0.23816854,0.27330816,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.31235218,0.37482262,0.43729305,0.4997635,0.5622339,0.737932,0.9136301,1.0893283,1.261122,1.43682,1.5500476,1.6632754,1.7765031,1.8858263,1.999054,1.8506867,1.698415,1.5500476,1.4016805,1.2494087,1.0112402,0.77307165,0.5388075,0.30063897,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,2.1122816,4.224563,6.336845,8.449126,10.561408,8.636538,6.7116675,4.786797,2.8619268,0.93705654,0.80040246,0.6637484,0.5231899,0.38653582,0.24988174,4.6110992,8.976221,13.337439,17.698656,22.063778,20.775324,19.486872,18.19842,16.91387,15.625418,18.38583,21.150146,23.914463,26.674877,29.439194,26.499178,23.563068,20.623053,17.686943,14.750832,28.802776,42.850815,56.898853,70.9508,84.99884,89.211685,93.42454,97.63739,101.850235,106.06309,91.09751,76.13975,61.174175,46.212505,31.250835,26.300053,21.349272,16.398489,11.4516115,6.5008297,5.774611,5.0483923,4.3260775,3.5998588,2.87364,2.3231194,1.7765031,1.2259823,0.6754616,0.12494087,0.58566034,1.0502841,1.5110037,1.9756275,2.436347,2.3231194,2.2137961,2.1005683,1.9873407,1.8741131,1.7999294,1.7257458,1.6515622,1.5734742,1.4992905,1.9482968,2.4012074,2.8502135,3.2992198,3.7482262,3.435874,3.1235218,2.8111696,2.4988174,2.1864653,1.7491722,1.3118792,0.8745861,0.43729305,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.37482262,0.3357786,0.30063897,0.26159495,0.22645533,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.38653582,0.5231899,0.6637484,0.80040246,0.93705654,0.74964523,0.5622339,0.37482262,0.18741131,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.093705654,0.08980125,0.08589685,0.078088045,0.07418364,0.19912452,0.32016098,0.44119745,0.5661383,0.6871748,0.59346914,0.5036679,0.40996224,0.31625658,0.22645533,0.1835069,0.14446288,0.10541886,0.06637484,0.023426414,0.3357786,0.6481308,0.96438736,1.2767396,1.5890918,1.3509232,1.116659,0.8823949,0.6481308,0.41386664,0.3318742,0.24597734,0.1639849,0.08199245,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.58956474,0.98000497,1.3704453,1.7608855,2.1513257,2.1083772,2.069333,2.0302892,1.9912452,1.9482968,1.8584955,1.7686942,1.678893,1.5890918,1.4992905,1.3548276,1.2103647,1.0659018,0.92143893,0.77307165,0.6676528,0.5583295,0.45291066,0.3435874,0.23816854,0.25769055,0.27721256,0.29673457,0.31625658,0.3357786,0.7066968,1.077615,1.4485333,1.8194515,2.1864653,1.8741131,1.5617609,1.2494087,0.93705654,0.62470436,1.5656652,2.5066261,3.4436827,4.3846436,5.3256044,5.446641,5.563773,5.6848097,5.805846,5.9268827,5.6809053,5.434928,5.1889505,4.9468775,4.7009,4.482254,4.263607,4.0488653,3.8302186,3.611572,3.39683,3.1781836,2.959537,2.7408905,2.5261483,2.2450314,1.9639144,1.6867018,1.4055848,1.1244678,1.0073358,0.8902037,0.77307165,0.6559396,0.5388075,0.71841,0.8980125,1.077615,1.2572175,1.43682,1.7257458,2.018576,2.3075018,2.5964274,2.8892577,2.3543546,1.8194515,1.2806439,0.74574083,0.21083772,0.28502136,0.359205,0.42948425,0.5036679,0.57394713,0.46071947,0.3513962,0.23816854,0.12494087,0.011713207,0.06637484,0.12103647,0.1756981,0.23426414,0.28892577,0.5192855,0.75354964,0.98390937,1.2181735,1.4485333,1.53443,1.6164225,1.698415,1.7804074,1.8623998,1.8467822,1.8272603,1.8116426,1.7921207,1.7765031,1.620327,1.4641509,1.3118792,1.1557031,0.999527,0.80821127,0.62079996,0.42948425,0.23816854,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.078088045,0.06637484,0.058566034,0.046852827,0.039044023,0.031235218,0.027330816,0.023426414,0.015617609,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.30844778,0.24597734,0.1796025,0.113227665,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,1.815547,3.631094,5.446641,7.2582836,9.073831,7.4183645,5.7668023,4.1113358,2.455869,0.80040246,0.679366,0.5583295,0.44119745,0.32016098,0.19912452,3.7091823,7.2153354,10.721489,14.231546,17.7377,16.921679,16.10566,15.293544,14.477524,13.661504,16.175938,18.694279,21.208714,23.723148,26.237583,24.820286,23.402987,21.98569,20.568392,19.151093,30.325493,41.499893,52.67429,63.84869,75.02309,77.88892,80.75475,83.62058,86.48641,89.34834,77.272026,65.199615,53.1233,41.050884,28.97457,24.601639,20.228708,15.855778,11.486752,7.113821,6.6257706,6.13772,5.64967,5.1616197,4.6735697,3.9473507,3.2211318,2.4910088,1.7647898,1.038571,1.2572175,1.475864,1.698415,1.9170616,2.135708,2.0107672,1.8858263,1.7608855,1.6359446,1.5110037,1.4485333,1.3860629,1.3235924,1.261122,1.1986516,1.5617609,1.9209659,2.280171,2.639376,2.998581,2.7486992,2.4988174,2.2489357,1.999054,1.7491722,1.4016805,1.0502841,0.698888,0.3513962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.027330816,0.042948425,0.058566034,0.07418364,0.08589685,0.14055848,0.19131571,0.24597734,0.29673457,0.3513962,0.31235218,0.27330816,0.23816854,0.19912452,0.1639849,0.14055848,0.12103647,0.10151446,0.08199245,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.30844778,0.42167544,0.5309987,0.64032197,0.74964523,0.62079996,0.48805028,0.359205,0.23035973,0.10151446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.08980125,0.10541886,0.12103647,0.13665408,0.14836729,0.39434463,0.64032197,0.8862993,1.1283722,1.3743496,1.1908426,1.0034313,0.8199245,0.63641757,0.44900626,0.3709182,0.28892577,0.21083772,0.12884527,0.05075723,0.61299115,1.175225,1.737459,2.2996929,2.8619268,2.455869,2.0459068,1.639849,1.2337911,0.8238289,0.659844,0.4958591,0.3318742,0.1639849,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.44119745,0.7340276,1.0268579,1.319688,1.6125181,1.5812829,1.5539521,1.5227169,1.4914817,1.4641509,1.3938715,1.3274968,1.261122,1.1908426,1.1244678,1.0229534,0.92143893,0.8160201,0.7145056,0.61299115,0.5466163,0.48414588,0.41777104,0.3513962,0.28892577,0.28892577,0.29283017,0.29673457,0.29673457,0.30063897,0.96438736,1.6281357,2.2957885,2.959537,3.6232853,3.0883822,2.5495746,2.0107672,1.475864,0.93705654,1.5539521,2.1708477,2.7916477,3.408543,4.025439,4.2284675,4.4314966,4.630621,4.83365,5.036679,5.0601053,5.083532,5.1030536,5.12648,5.1499066,5.0522966,4.9546866,4.8570766,4.759466,4.661856,4.3534083,4.041056,3.7326086,3.4241607,3.1118085,2.8775444,2.6432803,2.4090161,2.1708477,1.9365835,1.7647898,1.5929961,1.4212024,1.2494087,1.0737107,1.43682,1.796025,2.15523,2.514435,2.87364,2.8306916,2.7838387,2.7408905,2.6940374,2.6510892,2.1786566,1.7101282,1.2415999,0.76916724,0.30063897,0.40605783,0.5153811,0.62079996,0.7301232,0.8394465,0.6754616,0.5114767,0.3513962,0.18741131,0.023426414,0.08589685,0.14446288,0.20693332,0.26549935,0.3240654,0.7262188,1.1283722,1.53443,1.9365835,2.338737,2.3270237,2.3192148,2.3075018,2.2957885,2.2879796,2.1396124,1.9912452,1.8467822,1.698415,1.5500476,1.3899672,1.2298868,1.0698062,0.9097257,0.74964523,0.60908675,0.46462387,0.3240654,0.1796025,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.15617609,0.13665408,0.113227665,0.093705654,0.07418364,0.06637484,0.05466163,0.046852827,0.03513962,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.359205,0.27721256,0.19912452,0.11713207,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,1.5188124,3.0337205,4.552533,6.0713453,7.5862536,6.2040954,4.8180323,3.4319696,2.0459068,0.6637484,0.5583295,0.45681506,0.3553006,0.25378615,0.14836729,2.803361,5.45445,8.109444,10.760532,13.411622,13.068034,12.728352,12.384764,12.041177,11.701493,13.966047,16.234505,18.502962,20.77142,23.035973,23.141392,23.242907,23.344421,23.445936,23.551353,31.852114,40.148968,48.449726,56.75049,65.05125,66.566154,68.08497,69.60378,71.11869,72.6375,63.45044,54.263382,45.076324,35.889267,26.698303,22.903223,19.11205,15.313066,11.521891,7.726812,7.47693,7.223144,6.9732623,6.7233806,6.473499,5.571582,4.6657605,3.7599394,2.854118,1.9482968,1.9287747,1.9053483,1.8819219,1.8584955,1.8389735,1.698415,1.5617609,1.4251068,1.2884527,1.1517987,1.1010414,1.0502841,0.999527,0.94876975,0.9019169,1.1713207,1.4407244,1.7101282,1.979532,2.2489357,2.0615244,1.8741131,1.6867018,1.4992905,1.3118792,1.0502841,0.78868926,0.5231899,0.26159495,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.042948425,0.058566034,0.078088045,0.093705654,0.113227665,0.15617609,0.19912452,0.23816854,0.28111696,0.3240654,0.28892577,0.24988174,0.21083772,0.1756981,0.13665408,0.12103647,0.10932326,0.093705654,0.078088045,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.23426414,0.31625658,0.39824903,0.48024148,0.5622339,0.48805028,0.41777104,0.3435874,0.27330816,0.19912452,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.08589685,0.12103647,0.15617609,0.19131571,0.22645533,0.59346914,0.96048295,1.3274968,1.6945106,2.0615244,1.7843118,1.5070993,1.2298868,0.95267415,0.6754616,0.5544251,0.43338865,0.31625658,0.19522011,0.07418364,0.8862993,1.698415,2.514435,3.3265507,4.138666,3.5569105,2.979059,2.397303,1.815547,1.2376955,0.9917182,0.7418364,0.4958591,0.24597734,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.29673457,0.48805028,0.6832704,0.8784905,1.0737107,1.0541886,1.0346665,1.0151446,0.9956226,0.97610056,0.92924774,0.8862993,0.8394465,0.79649806,0.74964523,0.6910792,0.62860876,0.5700427,0.5114767,0.44900626,0.42557985,0.40605783,0.38263142,0.359205,0.3357786,0.3240654,0.30844778,0.29283017,0.27721256,0.26159495,1.2220778,2.182561,3.1430438,4.1035266,5.0640097,4.298747,3.5373883,2.77603,2.0107672,1.2494087,1.5461433,1.8389735,2.135708,2.4285383,2.7252727,3.0102942,3.2953155,3.5803368,3.8653584,4.1503797,4.4393053,4.728231,5.0210614,5.309987,5.5989127,5.6223392,5.645766,5.6691923,5.688714,5.7121406,5.309987,4.9078336,4.50568,4.1035266,3.7013733,3.5100577,3.3187418,3.1313305,2.9400148,2.7486992,2.522244,2.2957885,2.069333,1.8389735,1.6125181,2.1513257,2.6940374,3.232845,3.7716527,4.3143644,3.9317331,3.5530062,3.174279,2.7916477,2.4129205,2.0068626,1.6008049,1.1986516,0.79259366,0.38653582,0.5309987,0.6715572,0.8160201,0.95657855,1.1010414,0.8862993,0.6754616,0.46071947,0.24988174,0.039044023,0.10151446,0.1678893,0.23426414,0.29673457,0.3631094,0.93315214,1.5070993,2.0810463,2.6510892,3.2250361,3.1235218,3.018103,2.9165885,2.815074,2.7135596,2.436347,2.1591344,1.8819219,1.6008049,1.3235924,1.1596074,0.9956226,0.8316377,0.6637484,0.4997635,0.40605783,0.30844778,0.21474212,0.12103647,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10541886,0.15617609,0.21083772,0.26159495,0.23426414,0.20302892,0.1717937,0.14055848,0.113227665,0.09761006,0.08199245,0.06637484,0.05075723,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.40605783,0.30844778,0.21474212,0.12103647,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,1.2181735,2.4402514,3.6584249,4.8805027,6.098676,4.985922,3.8692627,2.7565079,1.639849,0.5231899,0.44119745,0.3553006,0.26940376,0.1835069,0.10151446,1.8975395,3.6935644,5.493494,7.289519,9.089449,9.218294,9.347139,9.475985,9.608734,9.737579,11.756155,13.778636,15.797212,17.815788,19.838268,21.458595,23.082827,24.703154,26.327385,27.951616,33.374832,38.798046,44.225163,49.64838,55.075497,55.24339,55.41518,55.586975,55.754864,55.92666,49.624954,43.327152,37.025448,30.723742,24.425941,21.208714,17.991486,14.774258,11.553126,8.335898,8.324185,8.312472,8.300759,8.289046,8.273428,7.191909,6.1103897,5.02887,3.9434462,2.8619268,2.5964274,2.330928,2.069333,1.8038338,1.5383345,1.3860629,1.2376955,1.0893283,0.93705654,0.78868926,0.74964523,0.7106012,0.6754616,0.63641757,0.60127795,0.78088045,0.96048295,1.1400855,1.319688,1.4992905,1.3743496,1.2494087,1.1244678,0.999527,0.8745861,0.698888,0.5231899,0.3513962,0.1756981,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.058566034,0.078088045,0.09761006,0.11713207,0.13665408,0.1717937,0.20302892,0.23426414,0.26940376,0.30063897,0.26159495,0.22645533,0.18741131,0.14836729,0.113227665,0.10151446,0.093705654,0.08199245,0.07418364,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.15617609,0.21083772,0.26549935,0.32016098,0.37482262,0.359205,0.3435874,0.3318742,0.31625658,0.30063897,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.078088045,0.13665408,0.19131571,0.24597734,0.30063897,0.78868926,1.2806439,1.7686942,2.260649,2.7486992,2.3816853,2.0107672,1.639849,1.2689307,0.9019169,0.7418364,0.58175594,0.42167544,0.26159495,0.10151446,1.1635119,2.2255092,3.2875066,4.349504,5.4115014,4.661856,3.9083066,3.154757,2.4012074,1.6515622,1.319688,0.9917182,0.659844,0.3318742,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.14836729,0.24597734,0.3435874,0.44119745,0.5388075,0.5270943,0.5192855,0.5075723,0.4958591,0.48805028,0.46462387,0.44119745,0.42167544,0.39824903,0.37482262,0.359205,0.339683,0.3240654,0.30454338,0.28892577,0.30844778,0.3279698,0.3474918,0.3670138,0.38653582,0.3553006,0.3240654,0.28892577,0.25769055,0.22645533,1.4797685,2.7330816,3.9902992,5.2436123,6.5008297,5.5130157,4.5252023,3.5373883,2.5495746,1.5617609,1.53443,1.5070993,1.4797685,1.4524376,1.4251068,1.7921207,2.1591344,2.5261483,2.893162,3.2640803,3.8185053,4.376835,4.9351645,5.493494,6.0518236,6.192382,6.336845,6.477403,6.621866,6.7624245,6.266566,5.7707067,5.278752,4.7828927,4.2870336,4.142571,3.998108,3.853645,3.7091823,3.5608149,3.279698,2.998581,2.7135596,2.4324427,2.1513257,2.8697357,3.5881457,4.31046,5.02887,5.7511845,5.036679,4.318269,3.6037633,2.8892577,2.174752,1.8350691,1.4953861,1.1557031,0.8160201,0.47633708,0.6520352,0.8316377,1.0073358,1.1869383,1.3626363,1.1010414,0.8394465,0.57394713,0.31235218,0.05075723,0.12103647,0.19131571,0.26159495,0.3318742,0.39824903,1.1439898,1.8858263,2.6276627,3.3694992,4.1113358,3.9161155,3.7208953,3.5256753,3.3343596,3.1391394,2.7291772,2.3231194,1.9131571,1.5070993,1.1010414,0.92924774,0.76135844,0.58956474,0.42167544,0.24988174,0.20302892,0.15617609,0.10932326,0.058566034,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07027924,0.14055848,0.21083772,0.28111696,0.3513962,0.30844778,0.26940376,0.23035973,0.19131571,0.14836729,0.12884527,0.10932326,0.08980125,0.07027924,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.113227665,0.22645533,0.3357786,0.44900626,0.5622339,0.45291066,0.3435874,0.23426414,0.12103647,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.92143893,1.8467822,2.7682211,3.68966,4.6110992,3.767748,2.9243972,2.077142,1.2337911,0.38653582,0.32016098,0.25378615,0.1835069,0.11713207,0.05075723,0.9917182,1.9365835,2.8775444,3.8185053,4.7633705,5.364649,5.9659266,6.571109,7.172387,7.773665,9.546264,11.318862,13.091461,14.864059,16.636658,19.779701,22.922745,26.06579,29.208834,32.351875,34.90145,37.451027,40.000603,42.550175,45.09975,43.92062,42.745396,41.566265,40.39104,39.21191,35.799465,32.387016,28.97457,25.562122,22.149673,19.510298,16.870922,14.231546,11.588266,8.94889,9.175345,9.4018,9.6243515,9.850807,10.073358,8.81614,7.5550184,6.2938967,5.036679,3.775557,3.2679846,2.7604125,2.25284,1.7452679,1.2376955,1.0737107,0.9136301,0.74964523,0.58566034,0.42557985,0.39824903,0.37482262,0.3513962,0.3240654,0.30063897,0.39044023,0.48024148,0.5700427,0.659844,0.74964523,0.6871748,0.62470436,0.5622339,0.4997635,0.43729305,0.3513962,0.26159495,0.1756981,0.08589685,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.07418364,0.093705654,0.11713207,0.14055848,0.1639849,0.1835069,0.20693332,0.23035973,0.25378615,0.27330816,0.23816854,0.19912452,0.1639849,0.12494087,0.08589685,0.08199245,0.078088045,0.07418364,0.06637484,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.078088045,0.10541886,0.13274968,0.16008049,0.18741131,0.23035973,0.27330816,0.31625658,0.359205,0.39824903,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.9878138,1.6008049,2.2137961,2.8267872,3.435874,2.9751544,2.514435,2.0498111,1.5890918,1.1244678,0.92534333,0.7262188,0.5231899,0.3240654,0.12494087,1.43682,2.7486992,4.0644827,5.376362,6.688241,5.7628975,4.8375545,3.912211,2.9868677,2.0615244,1.6515622,1.2376955,0.8238289,0.41386664,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.18741131,0.24988174,0.31235218,0.37482262,0.43729305,0.38653582,0.3357786,0.28892577,0.23816854,0.18741131,1.737459,3.2875066,4.8375545,6.387602,7.9376497,6.7233806,5.5130157,4.298747,3.0883822,1.8741131,1.5266213,1.175225,0.8238289,0.47633708,0.12494087,0.57394713,1.0268579,1.475864,1.9248703,2.3738766,3.2016098,4.025439,4.8492675,5.6730967,6.5008297,6.7624245,7.0240197,7.2856145,7.551114,7.812709,7.223144,6.6374836,6.0518236,5.462259,4.8765984,4.775084,4.6735697,4.575959,4.474445,4.376835,4.037152,3.7013733,3.3616903,3.0259118,2.6862288,3.5881457,4.4861584,5.388075,6.2860875,7.1880045,6.13772,5.087436,4.037152,2.9868677,1.9365835,1.6632754,1.3860629,1.1127546,0.8394465,0.5622339,0.77307165,0.9878138,1.1986516,1.4133936,1.6242313,1.3118792,0.999527,0.6871748,0.37482262,0.062470436,0.13665408,0.21083772,0.28892577,0.3631094,0.43729305,1.3509232,2.260649,3.174279,4.087909,5.001539,4.7126136,4.423688,4.138666,3.8497405,3.5608149,3.0259118,2.4871042,1.9482968,1.4133936,0.8745861,0.698888,0.5231899,0.3513962,0.1756981,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.38653582,0.3357786,0.28892577,0.23816854,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.0,0.0,0.0,0.0,0.0,0.0,0.62470436,1.2494087,1.8741131,2.4988174,3.1235218,2.5495746,1.9756275,1.4016805,0.8238289,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,1.5110037,2.5886188,3.6623292,4.73604,5.813655,7.336372,8.862993,10.38571,11.912332,13.438952,18.10081,22.762665,27.424522,32.086376,36.748234,36.424168,36.1001,35.77604,35.448067,35.124004,32.601757,30.075611,27.549461,25.023314,22.50107,21.973976,21.450787,20.92369,20.400501,19.873407,17.811884,15.750359,13.688834,11.623405,9.561881,10.0265045,10.487225,10.951848,11.412568,11.873287,10.436467,8.999647,7.562827,6.126007,4.689187,3.9356375,3.1859922,2.436347,1.6867018,0.93705654,0.76135844,0.58566034,0.41386664,0.23816854,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.10932326,0.21864653,0.3318742,0.44119745,0.5505207,0.4997635,0.44900626,0.39824903,0.3513962,0.30063897,0.98390937,1.6710842,2.3543546,3.0415294,3.7247996,3.1977055,2.6706111,2.1435168,1.6164225,1.0893283,1.2064602,1.3274968,1.4485333,1.5656652,1.6867018,2.4441557,3.1977055,3.951255,4.7087092,5.462259,4.7126136,3.9629683,3.213323,2.463678,1.7140326,1.3743496,1.038571,0.698888,0.3631094,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.14836729,0.19912452,0.24988174,0.30063897,0.3513962,0.31625658,0.28502136,0.25378615,0.21864653,0.18741131,1.4485333,2.7057507,3.9668727,5.2279944,6.4891167,5.571582,4.657952,3.7443218,2.8267872,1.9131571,1.6281357,1.3431144,1.0580931,0.77307165,0.48805028,0.8238289,1.1557031,1.4914817,1.8272603,2.1630387,2.8385005,3.5178664,4.193328,4.872694,5.548156,5.8292727,6.1103897,6.3915067,6.6687193,6.949836,6.5672045,6.184573,5.801942,5.4193106,5.036679,4.8883114,4.73604,4.5876727,4.4393053,4.2870336,3.8887846,3.49444,3.096191,2.697942,2.2996929,3.0337205,3.7716527,4.50568,5.239708,5.9737353,5.376362,4.7789884,4.181615,3.5842414,2.9868677,2.5027218,2.018576,1.53443,1.0463798,0.5622339,0.7301232,0.8980125,1.0659018,1.2337911,1.4016805,1.1400855,0.8784905,0.62079996,0.359205,0.10151446,0.15617609,0.21083772,0.26549935,0.32016098,0.37482262,1.1010414,1.8233559,2.5495746,3.2757936,3.998108,3.802888,3.6037633,3.408543,3.2094188,3.0141985,2.7565079,2.5027218,2.2489357,1.9912452,1.737459,1.397776,1.0580931,0.71841,0.37872702,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08589685,0.1717937,0.25378615,0.339683,0.42557985,0.37482262,0.3240654,0.27330816,0.22645533,0.1756981,0.19131571,0.20693332,0.21864653,0.23426414,0.24988174,0.20302892,0.15617609,0.10932326,0.058566034,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.031235218,0.046852827,0.06637484,0.08199245,0.10151446,0.19131571,0.28502136,0.37872702,0.46852827,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.0,0.0,0.0,0.0,0.0,0.4997635,0.999527,1.4992905,1.999054,2.4988174,2.3192148,2.1396124,1.9600099,1.7804074,1.6008049,1.358732,1.1205635,0.8784905,0.64032197,0.39824903,0.42167544,0.44119745,0.46071947,0.48024148,0.4997635,2.533957,4.5681505,6.606249,8.640442,10.674636,10.729298,10.780055,10.8308115,10.885473,10.936231,15.484859,20.033487,24.578213,29.12684,33.67547,33.13666,32.59395,32.05514,31.516335,30.973623,29.255686,27.533844,25.815908,24.094067,22.37613,21.610867,20.845604,20.080341,19.315079,18.549814,16.597614,14.645412,12.693212,10.741011,8.78881,9.023073,9.261242,9.499411,9.737579,9.975748,8.761478,7.5433054,6.329036,5.114767,3.900498,3.3226464,2.7447948,2.1669433,1.5890918,1.0112402,0.8472553,0.6832704,0.5192855,0.3513962,0.18741131,0.16008049,0.13274968,0.10541886,0.078088045,0.05075723,0.14836729,0.24988174,0.3513962,0.44900626,0.5505207,0.4997635,0.44900626,0.39824903,0.3513962,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.07027924,0.08980125,0.10932326,0.12884527,0.14836729,0.16008049,0.1717937,0.1796025,0.19131571,0.19912452,0.1717937,0.14055848,0.10932326,0.078088045,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.12884527,0.10932326,0.08980125,0.07027924,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.1756981,0.14055848,0.10932326,0.078088045,0.046852827,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.093705654,0.14055848,0.19131571,0.23816854,0.19131571,0.14055848,0.093705654,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.21864653,0.44119745,0.659844,0.8784905,1.1010414,0.92534333,0.74964523,0.57394713,0.39824903,0.22645533,0.98390937,1.7413634,2.4988174,3.2562714,4.0137253,3.4202564,2.8267872,2.233318,1.6437533,1.0502841,1.4914817,1.9287747,2.3699722,2.8111696,3.2484627,3.4475873,3.6467118,3.8419318,4.041056,4.2362766,3.6623292,3.0883822,2.5105307,1.9365835,1.3626363,1.1010414,0.8394465,0.57394713,0.31235218,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.113227665,0.14836729,0.18741131,0.22645533,0.26159495,0.24597734,0.23426414,0.21864653,0.20302892,0.18741131,1.1557031,2.1278992,3.096191,4.068387,5.036679,4.4197836,3.802888,3.1859922,2.5690966,1.9482968,1.7296503,1.5110037,1.2884527,1.0698062,0.8511597,1.0698062,1.2884527,1.5110037,1.7296503,1.9482968,2.4792955,3.0102942,3.541293,4.068387,4.5993857,4.8961205,5.196759,5.493494,5.7902284,6.086963,5.911265,5.7316628,5.5559645,5.376362,5.2006636,5.001539,4.7985106,4.5993857,4.4002614,4.2011366,3.7443218,3.2836022,2.8267872,2.3699722,1.9131571,2.4831998,3.0532427,3.6232853,4.193328,4.7633705,4.618908,4.474445,4.3260775,4.181615,4.037152,3.3421683,2.6471848,1.9522011,1.2572175,0.5622339,0.6832704,0.80821127,0.92924774,1.0541886,1.175225,0.96829176,0.76135844,0.5544251,0.3435874,0.13665408,0.1717937,0.20693332,0.24207294,0.27721256,0.31235218,0.8511597,1.3860629,1.9248703,2.463678,2.998581,2.893162,2.7838387,2.67842,2.5690966,2.463678,2.4910088,2.5183394,2.5456703,2.5730011,2.6003318,2.096664,1.5890918,1.0854238,0.58175594,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08199245,0.1639849,0.24597734,0.3318742,0.41386664,0.3631094,0.31235218,0.26159495,0.21083772,0.1639849,0.21864653,0.27330816,0.3279698,0.38263142,0.43729305,0.3553006,0.27330816,0.19131571,0.10932326,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.058566034,0.093705654,0.12884527,0.1639849,0.19912452,0.26159495,0.32016098,0.37872702,0.44119745,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.0,0.0,0.0,0.0,0.0,0.37482262,0.74964523,1.1244678,1.4992905,1.8741131,2.0888553,2.3035975,2.5183394,2.7330816,2.951728,2.5183394,2.0888553,1.6593709,1.2298868,0.80040246,0.75354964,0.7066968,0.6559396,0.60908675,0.5622339,3.5569105,6.551587,9.546264,12.54094,15.535617,14.118319,12.697116,11.275913,9.858616,8.437413,12.86891,17.300406,21.735807,26.167303,30.5988,29.845251,29.091702,28.334248,27.580698,26.823244,25.909613,24.995983,24.07845,23.164818,22.251188,21.243853,20.240421,19.233086,18.229654,17.226223,15.383345,13.540467,11.697589,9.854712,8.011833,8.023546,8.039165,8.050878,8.062591,8.074304,7.082586,6.0908675,5.099149,4.1035266,3.1118085,2.7057507,2.3035975,1.8975395,1.4914817,1.0893283,0.93315214,0.77697605,0.62079996,0.46852827,0.31235218,0.26940376,0.22645533,0.1835069,0.14055848,0.10151446,0.30063897,0.4997635,0.698888,0.9019169,1.1010414,0.999527,0.9019169,0.80040246,0.698888,0.60127795,0.48024148,0.359205,0.23816854,0.12103647,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.05075723,0.06637484,0.08199245,0.09761006,0.113227665,0.12103647,0.12884527,0.13665408,0.14055848,0.14836729,0.12884527,0.10541886,0.08199245,0.058566034,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.10932326,0.10932326,0.10541886,0.10151446,0.10151446,0.14836729,0.19912452,0.24988174,0.30063897,0.3513962,0.28502136,0.21864653,0.15617609,0.08980125,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.093705654,0.19131571,0.28502136,0.37872702,0.47633708,0.37872702,0.28502136,0.19131571,0.093705654,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.3318742,0.659844,0.9917182,1.319688,1.6515622,1.3509232,1.0502841,0.74964523,0.44900626,0.14836729,0.98000497,1.8116426,2.639376,3.4710135,4.298747,3.6428072,2.9868677,2.3270237,1.6710842,1.0112402,1.7725986,2.533957,3.2914112,4.0527697,4.814128,4.4510183,4.0918136,3.7326086,3.3734035,3.0141985,2.612045,2.2137961,1.8116426,1.4133936,1.0112402,0.8238289,0.63641757,0.44900626,0.26159495,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.1756981,0.1756981,0.1796025,0.1835069,0.1835069,0.18741131,0.8667773,1.5461433,2.2294137,2.9087796,3.5881457,3.2679846,2.9478238,2.6276627,2.3075018,1.9873407,1.8311646,1.678893,1.5227169,1.3665408,1.2142692,1.3157835,1.4212024,1.5266213,1.6320401,1.737459,2.1200905,2.5027218,2.8853533,3.2679846,3.6506162,3.9668727,4.279225,4.5954814,4.911738,5.22409,5.251421,5.278752,5.3060827,5.3334136,5.3607445,5.1108627,4.860981,4.6110992,4.3612175,4.1113358,3.5959544,3.076669,2.5612879,2.0420024,1.5266213,1.9287747,2.3348327,2.7408905,3.1469483,3.5491016,3.8575494,4.165997,4.474445,4.7789884,5.087436,4.181615,3.2757936,2.3738766,1.4680552,0.5622339,0.64032197,0.71841,0.79649806,0.8706817,0.94876975,0.79649806,0.64032197,0.48414588,0.3318742,0.1756981,0.19131571,0.20693332,0.21864653,0.23426414,0.24988174,0.60127795,0.94876975,1.3001659,1.6515622,1.999054,1.9834363,1.9639144,1.9482968,1.9287747,1.9131571,2.2216048,2.533957,2.8424048,3.1508527,3.4632049,2.7916477,2.1239948,1.4524376,0.78088045,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,0.3513962,0.30063897,0.24988174,0.19912452,0.14836729,0.24597734,0.339683,0.43338865,0.5309987,0.62470436,0.5075723,0.39044023,0.27330816,0.15617609,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.08980125,0.14055848,0.19522011,0.24597734,0.30063897,0.3279698,0.3553006,0.38263142,0.40996224,0.43729305,0.3513962,0.26159495,0.1756981,0.08589685,0.0,0.0,0.0,0.0,0.0,0.0,0.24988174,0.4997635,0.74964523,0.999527,1.2494087,1.8584955,2.4714866,3.0805733,3.68966,4.298747,3.6818514,3.0610514,2.4402514,1.8194515,1.1986516,1.0854238,0.96829176,0.8550641,0.7418364,0.62470436,4.579864,8.535024,12.490183,16.445343,20.400501,17.50734,14.614178,11.721016,8.831758,5.938596,10.256865,14.571229,18.889498,23.207767,27.526035,26.55384,25.585548,24.613352,23.64506,22.67677,22.563541,22.454218,22.344894,22.23557,22.126247,20.880743,19.635239,18.389734,17.14423,15.8987255,14.169076,12.435521,10.701966,8.968412,7.238762,7.0240197,6.813182,6.5984397,6.387602,6.1767645,5.4036927,4.6345253,3.8653584,3.096191,2.3231194,2.0927596,1.8584955,1.6281357,1.3938715,1.1635119,1.0190489,0.8706817,0.7262188,0.58175594,0.43729305,0.37872702,0.3240654,0.26549935,0.20693332,0.14836729,0.44900626,0.74964523,1.0502841,1.3509232,1.6515622,1.4992905,1.3509232,1.1986516,1.0502841,0.9019169,0.71841,0.5388075,0.359205,0.1796025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.03513962,0.046852827,0.05466163,0.06637484,0.07418364,0.078088045,0.08589685,0.08980125,0.093705654,0.10151446,0.08589685,0.07027924,0.05466163,0.039044023,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.08980125,0.10541886,0.12103647,0.13665408,0.14836729,0.22645533,0.30063897,0.37482262,0.44900626,0.5231899,0.42557985,0.3318742,0.23426414,0.13665408,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.14055848,0.28502136,0.42557985,0.5700427,0.7106012,0.5700427,0.42557985,0.28502136,0.14055848,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,0.32016098,0.23816854,0.16008049,0.078088045,0.0,0.44119745,0.8784905,1.319688,1.7608855,2.1981785,1.7765031,1.3509232,0.92534333,0.4997635,0.07418364,0.97610056,1.8819219,2.7838387,3.6857557,4.5876727,3.8653584,3.1430438,2.4207294,1.698415,0.97610056,2.0537157,3.135235,4.2167544,5.2943697,6.375889,5.4583545,4.5408196,3.6232853,2.7057507,1.7882162,1.5617609,1.33921,1.1127546,0.8862993,0.6637484,0.5505207,0.43729305,0.3240654,0.21083772,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.10932326,0.12884527,0.14836729,0.1678893,0.18741131,0.57785153,0.96829176,1.358732,1.7491722,2.135708,2.1161861,2.0927596,2.069333,2.0459068,2.0263848,1.9365835,1.8467822,1.7530766,1.6632754,1.5734742,1.5656652,1.5539521,1.5461433,1.53443,1.5266213,1.7608855,1.9951496,2.2294137,2.463678,2.7018464,3.0337205,3.3655949,3.697469,4.029343,4.3612175,4.5954814,4.825841,5.0601053,5.2943697,5.5247293,5.22409,4.9234514,4.6267166,4.3260775,4.025439,3.4475873,2.8697357,2.2918842,1.7140326,1.1361811,1.3782539,1.6164225,1.8584955,2.096664,2.338737,3.096191,3.8575494,4.618908,5.376362,6.13772,5.0210614,3.9083066,2.7916477,1.678893,0.5622339,0.59346914,0.62860876,0.659844,0.6910792,0.7262188,0.62079996,0.5192855,0.41777104,0.31625658,0.21083772,0.20693332,0.20302892,0.19912452,0.19131571,0.18741131,0.3513962,0.5114767,0.6754616,0.8355421,0.999527,1.0737107,1.1439898,1.2181735,1.2884527,1.3626363,1.9561055,2.5456703,3.1391394,3.7326086,4.3260775,3.4905357,2.6549935,1.8194515,0.98390937,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.078088045,0.15617609,0.23426414,0.30844778,0.38653582,0.3357786,0.28892577,0.23816854,0.18741131,0.13665408,0.27330816,0.40605783,0.5427119,0.679366,0.81211567,0.659844,0.5075723,0.3553006,0.20302892,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.12103647,0.19131571,0.26159495,0.3318742,0.39824903,0.39434463,0.39044023,0.38653582,0.37872702,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,1.6281357,2.6354716,3.638903,4.646239,5.64967,4.841459,4.029343,3.2211318,2.4090161,1.6008049,1.4172981,1.2337911,1.0541886,0.8706817,0.6871748,5.602817,10.518459,15.434102,20.34584,25.261482,20.89636,16.531239,12.166118,7.800996,3.435874,7.6409154,11.842052,16.043188,20.24823,24.449368,23.266333,22.079395,20.89636,19.709423,18.526388,19.221373,19.916355,20.61134,21.306324,22.001307,20.51373,19.030056,17.546383,16.058807,14.575133,12.950902,11.330575,9.706344,8.086017,6.461786,6.0244927,5.5871997,5.1499066,4.7126136,4.2753205,3.7287042,3.1781836,2.631567,2.084951,1.5383345,1.475864,1.4172981,1.358732,1.2962615,1.2376955,1.1010414,0.96829176,0.8316377,0.698888,0.5622339,0.48805028,0.41777104,0.3435874,0.27330816,0.19912452,0.60127795,0.999527,1.4016805,1.7999294,2.1981785,1.999054,1.7999294,1.6008049,1.4016805,1.1986516,0.96048295,0.71841,0.48024148,0.23816854,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.015617609,0.023426414,0.027330816,0.031235218,0.039044023,0.039044023,0.042948425,0.046852827,0.046852827,0.05075723,0.042948425,0.03513962,0.027330816,0.019522011,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.07027924,0.10151446,0.13665408,0.1678893,0.19912452,0.30063897,0.39824903,0.4997635,0.60127795,0.698888,0.5700427,0.44119745,0.30844778,0.1796025,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.19131571,0.37872702,0.5700427,0.76135844,0.94876975,0.76135844,0.5700427,0.37872702,0.19131571,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.5505207,1.1010414,1.6515622,2.1981785,2.7486992,2.1981785,1.6515622,1.1010414,0.5505207,0.0,0.97610056,1.9482968,2.9243972,3.900498,4.8765984,4.087909,3.2992198,2.5105307,1.7257458,0.93705654,2.338737,3.736513,5.138193,6.5359693,7.9376497,6.461786,4.985922,3.513962,2.0380979,0.5622339,0.5114767,0.46071947,0.41386664,0.3631094,0.31235218,0.27330816,0.23816854,0.19912452,0.1639849,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.28892577,0.38653582,0.48805028,0.58566034,0.6871748,0.96438736,1.2376955,1.5110037,1.7882162,2.0615244,2.0380979,2.0107672,1.9873407,1.9639144,1.9365835,1.8116426,1.6867018,1.5617609,1.43682,1.3118792,1.4016805,1.4875772,1.5734742,1.6632754,1.7491722,2.1005683,2.4480603,2.7994564,3.1508527,3.4983444,3.9356375,4.376835,4.814128,5.251421,5.688714,5.337318,4.985922,4.6384296,4.2870336,3.9356375,3.2992198,2.6628022,2.0263848,1.3860629,0.74964523,0.8238289,0.9019169,0.97610056,1.0502841,1.1244678,2.338737,3.5491016,4.7633705,5.9737353,7.1880045,5.8644123,4.5369153,3.213323,1.8858263,0.5622339,0.5505207,0.5388075,0.5231899,0.5114767,0.4997635,0.44900626,0.39824903,0.3513962,0.30063897,0.24988174,0.22645533,0.19912452,0.1756981,0.14836729,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.1639849,0.3240654,0.48805028,0.6481308,0.81211567,1.6867018,2.5612879,3.435874,4.3143644,5.1889505,4.1894236,3.1859922,2.1864653,1.1869383,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.3240654,0.27330816,0.22645533,0.1756981,0.12494087,0.30063897,0.47633708,0.6481308,0.8238289,0.999527,0.81211567,0.62470436,0.43729305,0.24988174,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.14836729,0.23816854,0.3240654,0.41386664,0.4997635,0.46071947,0.42557985,0.38653582,0.3513962,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.4016805,2.7994564,4.2011366,5.5989127,7.000593,6.001066,5.001539,3.998108,2.998581,1.999054,1.7491722,1.4992905,1.2494087,0.999527,0.74964523,6.6257706,12.497992,18.374117,24.250242,30.126368,24.285381,18.448301,12.611219,6.774138,0.93705654,5.024966,9.112875,13.200784,17.288692,21.376602,19.974922,18.573242,17.175465,15.773785,14.376009,15.875299,17.37459,18.87388,20.37317,21.876366,20.15062,18.424873,16.69913,14.973383,13.251541,11.736633,10.22563,8.710721,7.1997175,5.688714,5.024966,4.3612175,3.7013733,3.0376248,2.3738766,2.0498111,1.7257458,1.4016805,1.0737107,0.74964523,0.8628729,0.97610056,1.0893283,1.1986516,1.3118792,1.1869383,1.0619974,0.93705654,0.81211567,0.6871748,0.60127795,0.5114767,0.42557985,0.3357786,0.24988174,0.74964523,1.2494087,1.7491722,2.2489357,2.7486992,2.4988174,2.2489357,1.999054,1.7491722,1.4992905,1.1986516,0.9019169,0.60127795,0.30063897,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.37482262,0.4997635,0.62470436,0.74964523,0.8745861,0.7106012,0.5505207,0.38653582,0.22645533,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.23816854,0.47633708,0.7106012,0.94876975,1.1869383,0.94876975,0.7106012,0.47633708,0.23816854,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.1717937,0.24597734,0.31625658,0.39044023,0.46071947,0.3709182,0.27721256,0.1835069,0.093705654,0.0,0.0,0.0,0.0,0.0,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,0.32016098,0.23816854,0.16008049,0.078088045,0.0,0.45681506,0.9136301,1.3743496,1.8311646,2.2879796,1.9209659,1.5578566,1.1908426,0.8277333,0.46071947,1.3274968,2.194274,3.057147,3.9239242,4.786797,4.029343,3.2679846,2.5066261,1.7491722,0.9878138,2.0615244,3.1313305,4.2050414,5.278752,6.348558,5.1889505,4.025439,2.8619268,1.698415,0.5388075,0.49195468,0.44900626,0.40215343,0.359205,0.31235218,0.26940376,0.22645533,0.1835069,0.14055848,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.23035973,0.30844778,0.39044023,0.46852827,0.5505207,0.76916724,0.9917182,1.2103647,1.4290112,1.6515622,1.6281357,1.6086137,1.5890918,1.5695697,1.5500476,1.4485333,1.3509232,1.2494087,1.1517987,1.0502841,1.1205635,1.1908426,1.261122,1.3314011,1.4016805,1.678893,1.9600099,2.241127,2.5183394,2.7994564,3.2172275,3.6349986,4.0527697,4.4705405,4.8883114,4.6696653,4.4510183,4.2362766,4.01763,3.7989833,3.5764325,3.349977,3.1235218,2.900971,2.6745155,2.4831998,2.2918842,2.096664,1.9053483,1.7140326,2.8814487,4.0488653,5.2162814,6.3836975,7.551114,6.250948,4.950782,3.6506162,2.35045,1.0502841,1.6047094,2.1591344,2.7135596,3.2718892,3.8263142,3.1079042,2.3894942,1.6710842,0.95657855,0.23816854,0.26159495,0.28111696,0.30454338,0.3279698,0.3513962,0.28892577,0.22645533,0.1639849,0.10151446,0.039044023,0.16008049,0.28111696,0.40605783,0.5270943,0.6481308,1.3509232,2.0498111,2.7486992,3.4514916,4.1503797,3.349977,2.5495746,1.7491722,0.94876975,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.26159495,0.21864653,0.1796025,0.14055848,0.10151446,0.24207294,0.38653582,0.5270943,0.6715572,0.81211567,0.659844,0.5075723,0.3553006,0.20302892,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.30063897,0.5114767,0.7262188,0.93705654,1.1517987,0.97610056,0.80430686,0.63251317,0.46071947,0.28892577,0.23426414,0.1835069,0.12884527,0.078088045,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,1.1283722,2.260649,3.3890212,4.521298,5.64967,4.841459,4.029343,3.2211318,2.4090161,1.6008049,1.4016805,1.1986516,0.999527,0.80040246,0.60127795,5.899552,11.20173,16.500004,21.798277,27.100456,22.251188,17.40192,12.548749,7.699481,2.8502135,5.8292727,8.8083315,11.791295,14.770353,17.749413,16.636658,15.519999,14.40334,13.2905855,12.173926,13.634172,15.090515,16.546856,18.003199,19.463446,17.761126,16.058807,14.356487,12.654168,10.951848,9.823476,8.695104,7.5667315,6.4383593,5.3138914,4.7985106,4.2870336,3.775557,3.2640803,2.7486992,2.6588979,2.5690966,2.4792955,2.3894942,2.2996929,2.2567444,2.2137961,2.1708477,2.1318035,2.0888553,2.0615244,2.0341935,2.0068626,1.9756275,1.9482968,1.8428779,1.7335546,1.6281357,1.5188124,1.4133936,1.6554666,1.8975395,2.1396124,2.3816853,2.6237583,2.4714866,2.3153105,2.1591344,2.0068626,1.8506867,1.4953861,1.1400855,0.78478485,0.42948425,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.24207294,0.47243267,0.7027924,0.93315214,1.1635119,1.0034313,0.8472553,0.6910792,0.5309987,0.37482262,0.30454338,0.23426414,0.1639849,0.093705654,0.023426414,0.023426414,0.019522011,0.015617609,0.015617609,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.10151446,0.18741131,0.27330816,0.3631094,0.44900626,0.42948425,0.40996224,0.39044023,0.3709182,0.3513962,0.80040246,1.2494087,1.698415,2.1513257,2.6003318,2.2255092,1.8506867,1.475864,1.1010414,0.7262188,0.71841,0.7145056,0.7106012,0.7066968,0.698888,0.57394713,0.44510186,0.31625658,0.19131571,0.062470436,0.23816854,0.41777104,0.59346914,0.77307165,0.94876975,0.76135844,0.5700427,0.37872702,0.19131571,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19912452,0.3435874,0.48805028,0.63641757,0.78088045,0.92534333,0.7418364,0.5544251,0.3709182,0.1835069,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.3631094,0.7301232,1.0932326,1.4602464,1.8233559,1.6437533,1.4641509,1.2845483,1.1049459,0.92534333,1.678893,2.436347,3.1898966,3.9434462,4.7009,3.9668727,3.2367494,2.5027218,1.7686942,1.038571,1.7843118,2.5261483,3.2718892,4.01763,4.7633705,3.912211,3.0610514,2.2137961,1.3626363,0.5114767,0.47243267,0.43338865,0.39434463,0.3513962,0.31235218,0.26549935,0.21864653,0.1717937,0.12103647,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.1717937,0.23426414,0.29283017,0.3513962,0.41386664,0.57785153,0.7418364,0.9058213,1.0737107,1.2376955,1.2220778,1.2064602,1.1908426,1.1791295,1.1635119,1.0893283,1.0112402,0.93705654,0.8628729,0.78868926,0.8394465,0.8941081,0.94486535,0.9956226,1.0502841,1.261122,1.4680552,1.678893,1.8897307,2.1005683,2.4988174,2.893162,3.2914112,3.68966,4.087909,4.0020123,3.9161155,3.8341231,3.7482262,3.6623292,3.8497405,4.037152,4.224563,4.4119744,4.5993857,4.138666,3.6818514,3.2211318,2.7604125,2.2996929,3.4241607,4.5447245,5.6691923,6.7897553,7.914223,6.6374836,5.3607445,4.087909,2.8111696,1.5383345,2.6588979,3.7833657,4.903929,6.028397,7.1489606,5.7668023,4.380739,2.9946766,1.6086137,0.22645533,0.29673457,0.3631094,0.43338865,0.5036679,0.57394713,0.47633708,0.37482262,0.27330816,0.1756981,0.07418364,0.15617609,0.23816854,0.3240654,0.40605783,0.48805028,1.0112402,1.5383345,2.0615244,2.5886188,3.1118085,2.514435,1.9131571,1.3118792,0.7106012,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.08980125,0.13665408,0.1796025,0.22645533,0.19522011,0.1639849,0.13665408,0.10541886,0.07418364,0.1835069,0.29673457,0.40605783,0.5153811,0.62470436,0.5075723,0.39044023,0.27330816,0.15617609,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.44900626,0.78868926,1.1244678,1.4641509,1.7999294,1.4914817,1.1869383,0.8784905,0.5700427,0.26159495,0.21864653,0.1756981,0.13665408,0.093705654,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.8589685,1.7218413,2.5808098,3.4397783,4.298747,3.6818514,3.0610514,2.4402514,1.8194515,1.1986516,1.0502841,0.9019169,0.74964523,0.60127795,0.44900626,5.173333,9.901564,14.625891,19.350218,24.074545,20.21309,16.351637,12.486279,8.624825,4.7633705,6.6335793,8.507692,10.381805,12.252014,14.126127,13.29449,12.466757,11.6351185,10.803481,9.975748,11.389141,12.806439,14.219833,15.633226,17.050524,15.371632,13.688834,12.009941,10.331048,8.648251,7.9064145,7.164578,6.422742,5.6809053,4.939069,4.575959,4.21285,3.8497405,3.4866312,3.1235218,3.2718892,3.416352,3.5608149,3.7052777,3.8497405,3.6506162,3.455396,3.2562714,3.0610514,2.8619268,2.9322062,3.0024853,3.0727646,3.1430438,3.213323,3.084478,2.9556324,2.8306916,2.7018464,2.5769055,2.5612879,2.5456703,2.5300527,2.514435,2.4988174,2.4402514,2.3816853,2.3192148,2.260649,2.1981785,1.7882162,1.3782539,0.96829176,0.5583295,0.14836729,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.48414588,0.94486535,1.4055848,1.8663043,2.3231194,2.0107672,1.6945106,1.3782539,1.0659018,0.74964523,0.60908675,0.46852827,0.3318742,0.19131571,0.05075723,0.046852827,0.039044023,0.03513962,0.031235218,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.19912452,0.37482262,0.5505207,0.7262188,0.9019169,0.80821127,0.71841,0.62860876,0.5388075,0.44900626,1.2259823,1.999054,2.77603,3.5491016,4.3260775,3.736513,3.1508527,2.5612879,1.9756275,1.3860629,1.3899672,1.3938715,1.3938715,1.397776,1.4016805,1.1439898,0.8902037,0.63641757,0.37872702,0.12494087,0.24207294,0.359205,0.47633708,0.59346914,0.7106012,0.5700427,0.42557985,0.28502136,0.14055848,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.30063897,0.5192855,0.7340276,0.95267415,1.1713207,1.3860629,1.1088502,0.8316377,0.5544251,0.27721256,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.27330816,0.5466163,0.8160201,1.0893283,1.3626363,1.3665408,1.3743496,1.3782539,1.3821584,1.3860629,2.0341935,2.67842,3.3226464,3.9668727,4.6110992,3.9083066,3.2016098,2.4988174,1.7921207,1.0893283,1.5031948,1.9209659,2.338737,2.7565079,3.174279,2.639376,2.1005683,1.5617609,1.0268579,0.48805028,0.45291066,0.41777104,0.38263142,0.3474918,0.31235218,0.26159495,0.20693332,0.15617609,0.10151446,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.113227665,0.15617609,0.19522011,0.23426414,0.27330816,0.38653582,0.4958591,0.60518235,0.7145056,0.8238289,0.8160201,0.80430686,0.79649806,0.78478485,0.77307165,0.7262188,0.6754616,0.62470436,0.57394713,0.5231899,0.5583295,0.59346914,0.62860876,0.6637484,0.698888,0.8394465,0.98000497,1.1205635,1.261122,1.4016805,1.7765031,2.15523,2.533957,2.9087796,3.2875066,3.3343596,3.3812122,3.4280653,3.4788225,3.5256753,4.123049,4.7243266,5.3256044,5.9268827,6.524256,5.7980375,5.0718184,4.3416953,3.6154766,2.8892577,3.9668727,5.040583,6.1181984,7.195813,8.273428,7.0240197,5.774611,4.5252023,3.2757936,2.0263848,3.7130866,5.4036927,7.094299,8.784905,10.475512,8.421796,6.3719845,4.318269,2.2645533,0.21083772,0.3318742,0.44900626,0.5661383,0.6832704,0.80040246,0.6637484,0.5231899,0.38653582,0.24988174,0.113227665,0.15617609,0.19912452,0.23816854,0.28111696,0.3240654,0.6754616,1.0268579,1.3743496,1.7257458,2.0732377,1.6749885,1.2767396,0.8745861,0.47633708,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.12884527,0.10932326,0.08980125,0.07027924,0.05075723,0.12884527,0.20693332,0.28111696,0.359205,0.43729305,0.3553006,0.27330816,0.19131571,0.10932326,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.60127795,1.0619974,1.5266213,1.9873407,2.4480603,2.0068626,1.5656652,1.1205635,0.679366,0.23816854,0.20693332,0.1717937,0.14055848,0.10932326,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.58956474,1.1791295,1.7686942,2.358259,2.951728,2.5183394,2.0888553,1.6593709,1.2298868,0.80040246,0.698888,0.60127795,0.4997635,0.39824903,0.30063897,4.4510183,8.601398,12.751778,16.898252,21.048632,18.174992,15.3013525,12.423808,9.550168,6.676528,7.4417906,8.203149,8.968412,9.733675,10.498938,9.956225,9.40961,8.866898,8.320281,7.773665,9.148014,10.518459,11.892809,13.263254,14.637604,12.978233,11.322766,9.663396,8.007929,6.348558,5.9932575,5.6340523,5.278752,4.919547,4.564246,4.349504,4.138666,3.9239242,3.7130866,3.4983444,3.8809757,4.2597027,4.6384296,5.0210614,5.3997884,5.0483923,4.6930914,4.3416953,3.9902992,3.638903,3.8067923,3.970777,4.138666,4.3065557,4.474445,4.3260775,4.181615,4.0332475,3.8848803,3.736513,3.4632049,3.193801,2.920493,2.6471848,2.3738766,2.4090161,2.4441557,2.4792955,2.514435,2.5495746,2.084951,1.620327,1.1557031,0.6910792,0.22645533,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.7262188,1.4172981,2.1083772,2.795552,3.4866312,3.0141985,2.541766,2.069333,1.5969005,1.1244678,0.9136301,0.7066968,0.4958591,0.28502136,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.30063897,0.5622339,0.8238289,1.0893283,1.3509232,1.1908426,1.0307622,0.8706817,0.7106012,0.5505207,1.6515622,2.7486992,3.8497405,4.950782,6.0518236,5.251421,4.4510183,3.6506162,2.8502135,2.0498111,2.0615244,2.069333,2.0810463,2.0888553,2.1005683,1.717937,1.3353056,0.95267415,0.5700427,0.18741131,0.24597734,0.30063897,0.359205,0.41777104,0.47633708,0.37872702,0.28502136,0.19131571,0.093705654,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.39824903,0.6910792,0.98000497,1.2689307,1.5617609,1.8506867,1.4797685,1.1088502,0.7418364,0.3709182,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.1796025,0.359205,0.5388075,0.71841,0.9019169,1.0893283,1.2806439,1.4680552,1.6593709,1.8506867,2.3855898,2.920493,3.455396,3.9902992,4.5252023,3.8458362,3.1703746,2.4910088,1.815547,1.1361811,1.2259823,1.3157835,1.4055848,1.4992905,1.5890918,1.3626363,1.1361811,0.9136301,0.6871748,0.46071947,0.43338865,0.40215343,0.3709182,0.3435874,0.31235218,0.25378615,0.19912452,0.14055848,0.08199245,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.058566034,0.078088045,0.09761006,0.11713207,0.13665408,0.19131571,0.24597734,0.30063897,0.359205,0.41386664,0.40605783,0.40215343,0.39824903,0.39434463,0.38653582,0.3631094,0.3357786,0.31235218,0.28892577,0.26159495,0.28111696,0.29673457,0.31625658,0.3318742,0.3513962,0.42167544,0.48805028,0.5583295,0.62860876,0.698888,1.0580931,1.4133936,1.7725986,2.1318035,2.4871042,2.6667068,2.8463092,3.0259118,3.2094188,3.3890212,4.4002614,5.4115014,6.426646,7.437886,8.449126,7.453504,6.461786,5.466163,4.4705405,3.474918,4.50568,5.5403466,6.571109,7.605776,8.636538,7.4144597,6.1884775,4.9624953,3.736513,2.514435,4.7711797,7.027924,9.284669,11.541413,13.798158,11.080693,8.359325,5.6418614,2.920493,0.19912452,0.3631094,0.5309987,0.6949836,0.8589685,1.0268579,0.8511597,0.6754616,0.4997635,0.3240654,0.14836729,0.15227169,0.15617609,0.15617609,0.16008049,0.1639849,0.3357786,0.5114767,0.6871748,0.8628729,1.038571,0.8355421,0.63641757,0.43729305,0.23816854,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.06637484,0.05466163,0.046852827,0.03513962,0.023426414,0.07027924,0.113227665,0.16008049,0.20693332,0.24988174,0.20302892,0.15617609,0.10932326,0.058566034,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.06637484,0.09761006,0.12884527,0.1639849,0.74964523,1.33921,1.9248703,2.514435,3.1000953,2.522244,1.9443923,1.3665408,0.78868926,0.21083772,0.19131571,0.1678893,0.14446288,0.12103647,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.32016098,0.64032197,0.96048295,1.2806439,1.6008049,1.358732,1.1205635,0.8784905,0.64032197,0.39824903,0.3513962,0.30063897,0.24988174,0.19912452,0.14836729,3.7247996,7.3012323,10.87376,14.450192,18.026625,16.136894,14.251068,12.361338,10.475512,8.58578,8.246098,7.90251,7.558923,7.2192397,6.8756523,6.6140575,6.356367,6.094772,5.833177,5.575486,6.9068875,8.234385,9.565785,10.893282,12.224684,10.588739,8.956698,7.320754,5.6848097,4.0488653,4.0761957,4.1035266,4.1308575,4.1581883,4.1894236,4.123049,4.0605783,3.998108,3.9356375,3.873167,4.4900627,5.1030536,5.7199492,6.336845,6.949836,6.4422636,5.9346914,5.4271193,4.919547,4.4119744,4.677474,4.942973,5.2084727,5.473972,5.7394714,5.571582,5.4036927,5.2358036,5.067914,4.900025,4.369026,3.8419318,3.310933,2.7799344,2.2489357,2.3816853,2.5105307,2.639376,2.7682211,2.900971,2.3816853,1.8584955,1.33921,0.8199245,0.30063897,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.96829176,1.8897307,2.8111696,3.7287042,4.650143,4.0215344,3.3890212,2.7604125,2.1318035,1.4992905,1.2181735,0.94096094,0.659844,0.37872702,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.39824903,0.74964523,1.1010414,1.4485333,1.7999294,1.5695697,1.33921,1.1088502,0.8784905,0.6481308,2.0732377,3.4983444,4.9234514,6.348558,7.773665,6.7624245,5.7511845,4.73604,3.7247996,2.7135596,2.7291772,2.7486992,2.7643168,2.7838387,2.7994564,2.2918842,1.7804074,1.2689307,0.76135844,0.24988174,0.24597734,0.24597734,0.24207294,0.23816854,0.23816854,0.19131571,0.14055848,0.093705654,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4997635,0.8628729,1.2259823,1.5890918,1.9482968,2.3114061,1.8506867,1.3860629,0.92534333,0.46071947,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.81211567,1.1869383,1.5617609,1.9365835,2.3114061,2.736986,3.1625657,3.5881457,4.0137253,4.4393053,3.78727,3.1391394,2.4871042,1.8389735,1.1869383,0.94876975,0.7106012,0.47633708,0.23816854,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.41386664,0.38653582,0.3631094,0.3357786,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3357786,0.6754616,1.0112402,1.3509232,1.6867018,1.999054,2.3114061,2.6237583,2.9361105,3.2484627,4.6735697,6.098676,7.523783,8.94889,10.373997,9.112875,7.8517528,6.5867267,5.3256044,4.0605783,5.0483923,6.036206,7.0240197,8.011833,8.999647,7.800996,6.5984397,5.3997884,4.2011366,2.998581,5.825368,8.648251,11.475039,14.301826,17.124708,13.735687,10.350571,6.9615493,3.5764325,0.18741131,0.39824903,0.61299115,0.8238289,1.038571,1.2494087,1.038571,0.8238289,0.61299115,0.39824903,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.9019169,1.6125181,2.3231194,3.0376248,3.7482262,3.0376248,2.3231194,1.6125181,0.9019169,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,2.998581,6.001066,8.999647,11.998228,15.000713,14.098797,13.200784,12.298867,11.400854,10.498938,9.050405,7.601871,6.1494336,4.7009,3.2484627,3.2757936,3.2992198,3.3265507,3.349977,3.3734035,4.661856,5.950309,7.238762,8.52331,9.811763,8.1992445,6.5867267,4.9742084,3.3616903,1.7491722,2.1630387,2.5769055,2.9868677,3.4007344,3.8106966,3.900498,3.9863946,4.0761957,4.1620927,4.251894,5.099149,5.950309,6.801469,7.648724,8.499884,7.8361354,7.1762915,6.5125427,5.8487945,5.1889505,5.548156,5.911265,6.2743745,6.6374836,7.000593,6.813182,6.6257706,6.4383593,6.250948,6.0635366,5.2748475,4.4861584,3.7013733,2.912684,2.1239948,2.35045,2.5769055,2.7994564,3.0259118,3.2484627,2.6745155,2.1005683,1.5266213,0.94876975,0.37482262,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,1.2142692,2.3621633,3.513962,4.661856,5.813655,5.024966,4.2362766,3.4514916,2.6628022,1.8741131,1.5266213,1.175225,0.8238289,0.47633708,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.4997635,0.93705654,1.3743496,1.8116426,2.2489357,1.9482968,1.6515622,1.3509232,1.0502841,0.74964523,2.4988174,4.251894,6.001066,7.7502384,9.499411,8.273428,7.0513506,5.825368,4.5993857,3.3734035,3.4007344,3.4241607,3.4514916,3.474918,3.4983444,2.8619268,2.2255092,1.5890918,0.94876975,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.39824903,0.6910792,0.98000497,1.2689307,1.5617609,1.8506867,1.4797685,1.1088502,0.7418364,0.3709182,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23426414,0.46852827,0.7066968,0.94096094,1.175225,1.1205635,1.0659018,1.0112402,0.95657855,0.9019169,1.0893283,1.2806439,1.4680552,1.6593709,1.8506867,2.4910088,3.135235,3.7794614,4.4197836,5.0640097,4.240181,3.416352,2.5964274,1.7725986,0.94876975,0.76916724,0.58956474,0.40996224,0.23035973,0.05075723,0.13274968,0.21474212,0.29673457,0.37872702,0.46071947,0.42167544,0.37872702,0.3357786,0.29283017,0.24988174,0.20693332,0.1639849,0.12103647,0.078088045,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26940376,0.5388075,0.80821127,1.0815194,1.3509232,1.6008049,1.8506867,2.1005683,2.35045,2.6003318,3.7443218,4.8883114,6.036206,7.180196,8.324185,7.3441806,6.364176,5.3841705,4.4041657,3.4241607,4.2167544,5.009348,5.801942,6.5945354,7.387129,6.4422636,5.4973984,4.552533,3.6076677,2.6628022,4.9937305,7.328563,9.659492,11.994324,14.325252,11.560935,8.796618,6.028397,3.2640803,0.4997635,0.61689556,0.7340276,0.8511597,0.96829176,1.0893283,0.95657855,0.8238289,0.6910792,0.5583295,0.42557985,0.339683,0.25378615,0.1717937,0.08589685,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.019522011,0.015617609,0.015617609,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.7340276,1.319688,1.9053483,2.4910088,3.076669,2.5261483,1.9756275,1.4251068,0.8745861,0.3240654,0.28502136,0.24597734,0.20693332,0.1639849,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,2.4597735,4.845363,7.230953,9.616543,11.998228,11.291532,10.584834,9.878138,9.171441,8.460839,7.289519,6.1181984,4.9468775,3.7716527,2.6003318,2.7565079,2.9165885,3.0727646,3.2289407,3.3890212,4.646239,5.9073606,7.168483,8.4257,9.686822,8.769287,7.8478484,6.9264097,6.008875,5.087436,4.845363,4.60329,4.3612175,4.1191444,3.873167,3.8419318,3.8067923,3.7716527,3.736513,3.7013733,4.3534083,5.009348,5.6652875,6.321227,6.9732623,6.5945354,6.2158084,5.833177,5.45445,5.0757227,5.5676775,6.0596323,6.551587,7.043542,7.5394006,7.012306,6.4891167,5.9620223,5.4388323,4.911738,4.279225,3.6428072,3.0063896,2.3738766,1.737459,1.9365835,2.135708,2.338737,2.5378613,2.736986,2.4988174,2.260649,2.0263848,1.7882162,1.5500476,1.4290112,1.3040704,1.183034,1.0580931,0.93705654,1.7140326,2.4871042,3.2640803,4.037152,4.814128,4.2284675,3.6428072,3.057147,2.4714866,1.8858263,1.8194515,1.7491722,1.678893,1.6086137,1.5383345,1.2767396,1.0190489,0.75745404,0.4958591,0.23816854,0.22645533,0.21864653,0.20693332,0.19912452,0.18741131,0.1717937,0.15227169,0.13665408,0.11713207,0.10151446,0.093705654,0.08980125,0.08589685,0.078088045,0.07418364,0.30063897,0.5309987,0.75745404,0.98390937,1.2142692,1.1517987,1.0893283,1.0268579,0.96438736,0.9019169,1.1713207,1.4446288,1.717937,1.9912452,2.260649,2.639376,3.0141985,3.3890212,3.7638438,4.138666,5.630148,7.1216297,8.617016,10.108498,11.599979,9.8195715,8.039165,6.2587566,4.478349,2.7018464,2.7252727,2.7486992,2.77603,2.7994564,2.8267872,2.3114061,1.7999294,1.2884527,0.77697605,0.26159495,0.22255093,0.1835069,0.14055848,0.10151446,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.30063897,0.5192855,0.7340276,0.95267415,1.1713207,1.3860629,1.1088502,0.8316377,0.5544251,0.27721256,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.46852827,0.94096094,1.4094892,1.8819219,2.35045,2.1513257,1.9561055,1.756981,1.5617609,1.3626363,1.3665408,1.3743496,1.3782539,1.3821584,1.3860629,2.2489357,3.1079042,3.9668727,4.825841,5.688714,4.6930914,3.697469,2.7018464,1.7062237,0.7106012,0.58956474,0.46852827,0.3435874,0.22255093,0.10151446,0.1756981,0.25378615,0.3318742,0.40996224,0.48805028,0.42557985,0.3670138,0.30844778,0.24597734,0.18741131,0.1639849,0.14055848,0.12103647,0.09761006,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.20302892,0.40605783,0.60908675,0.80821127,1.0112402,1.1986516,1.3860629,1.5734742,1.7608855,1.9482968,2.815074,3.6818514,4.5447245,5.4115014,6.2743745,5.579391,4.8805027,4.181615,3.4866312,2.787743,3.3851168,3.9824903,4.579864,5.1772375,5.774611,5.083532,4.396357,3.7052777,3.0141985,2.3231194,4.165997,6.0049706,7.843944,9.686822,11.525795,9.382278,7.238762,5.099149,2.9556324,0.81211567,0.8355421,0.8589685,0.8784905,0.9019169,0.92534333,0.8706817,0.8199245,0.76916724,0.7145056,0.6637484,0.5309987,0.39824903,0.26549935,0.13274968,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.046852827,0.039044023,0.03513962,0.031235218,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.5700427,1.0268579,1.4836729,1.9443923,2.4012074,2.0107672,1.6242313,1.2376955,0.8511597,0.46071947,0.39434463,0.3279698,0.26159495,0.19131571,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,1.9209659,3.68966,5.4583545,7.230953,8.999647,8.484266,7.968885,7.453504,6.9381227,6.426646,5.5286336,4.6345253,3.7404175,2.8463092,1.9482968,2.241127,2.5300527,2.8189783,3.1118085,3.4007344,4.6345253,5.8644123,7.098203,8.32809,9.561881,9.335425,9.108971,8.878611,8.652155,8.4257,7.5276875,6.629675,5.7316628,4.83365,3.9356375,3.7794614,3.6232853,3.4632049,3.3070288,3.1508527,3.611572,4.068387,4.5291066,4.989826,5.4505453,5.3529353,5.2553253,5.1577153,5.0601053,4.9624953,5.5832953,6.2079997,6.8287997,7.453504,8.074304,7.211431,6.348558,5.4856853,4.6267166,3.7638438,3.279698,2.7994564,2.3153105,1.8311646,1.3509232,1.5266213,1.698415,1.8741131,2.0498111,2.2255092,2.3231194,2.4246337,2.5261483,2.6237583,2.7252727,2.541766,2.358259,2.1786566,1.9951496,1.8116426,2.2137961,2.612045,3.0141985,3.4124475,3.8106966,3.4280653,3.049338,2.6667068,2.2840753,1.901444,2.1083772,2.3192148,2.5300527,2.7408905,2.951728,2.4441557,1.9365835,1.4290112,0.92143893,0.41386664,0.39434463,0.3709182,0.3513962,0.3318742,0.31235218,0.27721256,0.24207294,0.20693332,0.1717937,0.13665408,0.12884527,0.11713207,0.10932326,0.09761006,0.08589685,0.5544251,1.0229534,1.4914817,1.9561055,2.4246337,2.2879796,2.1513257,2.0107672,1.8741131,1.737459,1.8467822,1.9522011,2.0615244,2.1669433,2.2762666,3.3265507,4.376835,5.423215,6.473499,7.523783,8.761478,9.99527,11.229061,12.466757,13.700547,11.365715,9.030883,6.6960497,4.3612175,2.0263848,2.0498111,2.0732377,2.1005683,2.1239948,2.1513257,1.7608855,1.3743496,0.9878138,0.60127795,0.21083772,0.19522011,0.1756981,0.16008049,0.14055848,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19912452,0.3435874,0.48805028,0.63641757,0.78088045,0.92534333,0.7418364,0.5544251,0.3709182,0.1835069,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7066968,1.4094892,2.1161861,2.8189783,3.5256753,3.1859922,2.8463092,2.5066261,2.1630387,1.8233559,1.6437533,1.4641509,1.2845483,1.1049459,0.92534333,2.0029583,3.0805733,4.1581883,5.2358036,6.3134184,5.1460023,3.978586,2.8111696,1.6437533,0.47633708,0.40996224,0.3435874,0.28111696,0.21474212,0.14836729,0.22255093,0.29673457,0.3670138,0.44119745,0.5114767,0.43338865,0.359205,0.28111696,0.20302892,0.12494087,0.12103647,0.12103647,0.11713207,0.113227665,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13665408,0.26940376,0.40605783,0.5388075,0.6754616,0.80040246,0.92534333,1.0502841,1.175225,1.3001659,1.8858263,2.4714866,3.0532427,3.638903,4.224563,3.8106966,3.39683,2.979059,2.5651922,2.1513257,2.5534792,2.9556324,3.357786,3.7599394,4.1620927,3.7287042,3.2914112,2.8580225,2.4207294,1.9873407,3.3343596,4.6813784,6.028397,7.37932,8.726339,7.2036223,5.6848097,4.165997,2.6432803,1.1244678,1.0541886,0.98000497,0.9058213,0.8355421,0.76135844,0.78868926,0.8160201,0.8433509,0.8706817,0.9019169,0.71841,0.5388075,0.359205,0.1796025,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.40605783,0.7340276,1.0659018,1.3938715,1.7257458,1.4992905,1.2767396,1.0502841,0.8238289,0.60127795,0.5036679,0.40996224,0.31625658,0.21864653,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.046852827,0.08980125,0.13665408,0.1796025,0.22645533,1.3782539,2.533957,3.68966,4.845363,6.001066,5.677001,5.35684,5.0327744,4.7087092,4.388548,3.7716527,3.1508527,2.533957,1.9170616,1.3001659,1.7218413,2.1435168,2.5690966,2.9907722,3.4124475,4.618908,5.8214636,7.027924,8.234385,9.43694,9.901564,10.366188,10.8308115,11.29934,11.763964,10.2100115,8.65606,7.1060123,5.55206,3.998108,3.7208953,3.4397783,3.1586614,2.8814487,2.6003318,2.8658314,3.1313305,3.39683,3.6584249,3.9239242,4.1113358,4.2948427,4.478349,4.6657605,4.8492675,5.602817,6.356367,7.1060123,7.859562,8.6131115,7.4105554,6.211904,5.0132523,3.8106966,2.612045,2.2840753,1.9522011,1.6242313,1.2923572,0.96438736,1.1127546,1.261122,1.4133936,1.5617609,1.7140326,2.1513257,2.5886188,3.0259118,3.4632049,3.900498,3.6584249,3.416352,3.174279,2.9283018,2.6862288,2.7135596,2.736986,2.7643168,2.787743,2.8111696,2.631567,2.4519646,2.2723622,2.0927596,1.9131571,2.4012074,2.893162,3.3812122,3.873167,4.3612175,3.6076677,2.854118,2.096664,1.3431144,0.58566034,0.5583295,0.5270943,0.4958591,0.46852827,0.43729305,0.38653582,0.3318742,0.28111696,0.22645533,0.1756981,0.16008049,0.14446288,0.12884527,0.113227665,0.10151446,0.80821127,1.5149081,2.2216048,2.9283018,3.638903,3.4241607,3.213323,2.998581,2.787743,2.5769055,2.5183394,2.4597735,2.4012074,2.3465457,2.2879796,4.0137253,5.735567,7.461313,9.187058,10.912805,11.888905,12.86891,13.845011,14.821111,15.801116,12.907954,10.018696,7.1294384,4.240181,1.3509232,1.3743496,1.4016805,1.4251068,1.4485333,1.475864,1.2142692,0.94876975,0.6871748,0.42557985,0.1639849,0.1678893,0.1717937,0.1756981,0.1835069,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.1717937,0.24597734,0.31625658,0.39044023,0.46071947,0.3709182,0.27721256,0.1835069,0.093705654,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.94096094,1.8819219,2.8189783,3.7599394,4.7009,4.2167544,3.736513,3.252367,2.7682211,2.2879796,1.9209659,1.5578566,1.1908426,0.8277333,0.46071947,1.756981,3.0532427,4.3455997,5.6418614,6.9381227,5.5989127,4.2557983,2.9165885,1.5773785,0.23816854,0.23035973,0.22255093,0.21474212,0.20693332,0.19912452,0.26940376,0.3357786,0.40215343,0.46852827,0.5388075,0.44119745,0.3474918,0.25378615,0.15617609,0.062470436,0.078088045,0.09761006,0.113227665,0.13274968,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06637484,0.13665408,0.20302892,0.26940376,0.3357786,0.39824903,0.46071947,0.5231899,0.58566034,0.6481308,0.95657855,1.261122,1.5656652,1.8702087,2.174752,2.0420024,1.9092526,1.7765031,1.6437533,1.5110037,1.7218413,1.9287747,2.135708,2.3426414,2.5495746,2.3699722,2.1903696,2.0107672,1.8311646,1.6515622,2.5066261,3.3616903,4.2167544,5.0718184,5.9268827,5.02887,4.1308575,3.232845,2.3348327,1.43682,1.2689307,1.1010414,0.93315214,0.76916724,0.60127795,0.7066968,0.8160201,0.92143893,1.0307622,1.1361811,0.9097257,0.6832704,0.45681506,0.22645533,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.23816854,0.44119745,0.6442264,0.8472553,1.0502841,0.9878138,0.92534333,0.8628729,0.80040246,0.737932,0.61689556,0.49195468,0.3709182,0.24597734,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.8394465,1.3782539,1.9209659,2.4597735,2.998581,2.8697357,2.7408905,2.6081407,2.4792955,2.35045,2.0107672,1.6710842,1.3314011,0.9917182,0.6481308,1.2064602,1.7608855,2.3153105,2.8697357,3.4241607,4.60329,5.7785153,6.957645,8.136774,9.311999,10.471607,11.62731,12.786918,13.94262,15.098324,12.892336,10.686349,8.476458,6.27047,4.0605783,3.6584249,3.2562714,2.854118,2.4519646,2.0498111,2.1200905,2.1903696,2.260649,2.330928,2.4012074,2.8658314,3.3343596,3.802888,4.271416,4.73604,5.618435,6.5008297,7.3832245,8.265619,9.151918,7.6135845,6.0752497,4.5369153,2.998581,1.4641509,1.2845483,1.1088502,0.92924774,0.75354964,0.57394713,0.698888,0.8238289,0.94876975,1.0737107,1.1986516,1.9756275,2.7486992,3.5256753,4.298747,5.0757227,4.7711797,4.4705405,4.165997,3.8653584,3.5608149,3.213323,2.8619268,2.514435,2.1630387,1.8116426,1.8350691,1.8584955,1.8819219,1.901444,1.9248703,2.6940374,3.4632049,4.2362766,5.0054436,5.774611,4.7711797,3.7716527,2.7682211,1.7647898,0.76135844,0.7223144,0.6832704,0.6442264,0.60127795,0.5622339,0.49195468,0.42167544,0.3513962,0.28111696,0.21083772,0.19131571,0.1717937,0.15227169,0.13274968,0.113227665,1.0619974,2.0068626,2.9556324,3.9044023,4.8492675,4.564246,4.2753205,3.9863946,3.7013733,3.4124475,3.1898966,2.9673457,2.7447948,2.522244,2.2996929,4.7009,7.098203,9.499411,11.900618,14.301826,15.020235,15.738646,16.46096,17.17937,17.901684,14.454097,11.010414,7.5667315,4.1191444,0.6754616,0.698888,0.7262188,0.74964523,0.77307165,0.80040246,0.6637484,0.5231899,0.38653582,0.24988174,0.113227665,0.14055848,0.1678893,0.19522011,0.22255093,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.175225,2.35045,3.5256753,4.7009,5.8761253,5.251421,4.6267166,3.998108,3.3734035,2.7486992,2.1981785,1.6515622,1.1010414,0.5505207,0.0,1.5110037,3.0259118,4.5369153,6.0518236,7.562827,6.0518236,4.5369153,3.0259118,1.5110037,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.31235218,0.37482262,0.43729305,0.4997635,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.27330816,0.42557985,0.57394713,0.7262188,0.8745861,0.8862993,0.9019169,0.9136301,0.92534333,0.93705654,1.0112402,1.0893283,1.1635119,1.2376955,1.3118792,1.6749885,2.0380979,2.4012074,2.7643168,3.1235218,2.8502135,2.5769055,2.2996929,2.0263848,1.7491722,1.4875772,1.2259823,0.96438736,0.698888,0.43729305,0.62470436,0.81211567,0.999527,1.1869383,1.3743496,1.1010414,0.8238289,0.5505207,0.27330816,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.47633708,0.57394713,0.6754616,0.77307165,0.8745861,0.7262188,0.57394713,0.42557985,0.27330816,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.6871748,1.3743496,2.0615244,2.7486992,3.435874,4.5876727,5.735567,6.8873653,8.039165,9.187058,11.037745,12.888432,14.739119,16.585901,18.436588,15.57466,12.712734,9.850807,6.98888,4.123049,3.5998588,3.076669,2.5495746,2.0263848,1.4992905,1.3743496,1.2494087,1.1244678,0.999527,0.8745861,1.6242313,2.3738766,3.1235218,3.873167,4.6267166,5.6379566,6.649197,7.6643414,8.675582,9.686822,7.812709,5.938596,4.0605783,2.1864653,0.31235218,0.28892577,0.26159495,0.23816854,0.21083772,0.18741131,0.28892577,0.38653582,0.48805028,0.58566034,0.6871748,1.7999294,2.912684,4.025439,5.138193,6.250948,5.8878384,5.5247293,5.1616197,4.7985106,4.4393053,3.7130866,2.9868677,2.260649,1.5383345,0.81211567,1.038571,1.261122,1.4875772,1.7140326,1.9365835,2.9868677,4.037152,5.087436,6.13772,7.1880045,5.938596,4.689187,3.435874,2.1864653,0.93705654,0.8862993,0.8394465,0.78868926,0.737932,0.6871748,0.60127795,0.5114767,0.42557985,0.3357786,0.24988174,0.22645533,0.19912452,0.1756981,0.14836729,0.12494087,1.3118792,2.4988174,3.6857557,4.8765984,6.0635366,5.700427,5.337318,4.9742084,4.6110992,4.251894,3.8614538,3.474918,3.0883822,2.7018464,2.3114061,5.388075,8.460839,11.537509,14.614178,17.686943,18.151566,18.612286,19.07691,19.537628,19.998348,16.00024,11.998228,8.00012,3.998108,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.113227665,0.1639849,0.21083772,0.26159495,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.94096094,1.8780174,2.8189783,3.7599394,4.7009,4.2089458,3.7130866,3.2211318,2.7291772,2.2372224,1.9092526,1.5773785,1.2494087,0.91753453,0.58566034,1.678893,2.7721257,3.8653584,4.958591,6.0518236,4.8570766,3.6662338,2.4714866,1.2806439,0.08589685,0.10932326,0.13274968,0.15617609,0.1756981,0.19912452,0.24988174,0.30063897,0.3513962,0.39824903,0.44900626,0.38653582,0.3240654,0.26159495,0.19912452,0.13665408,0.18741131,0.23816854,0.28892577,0.3357786,0.38653582,0.30844778,0.23426414,0.15617609,0.078088045,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.08199245,0.06637484,0.046852827,0.031235218,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.21864653,0.339683,0.46071947,0.58175594,0.698888,0.7106012,0.71841,0.7301232,0.7418364,0.74964523,0.8160201,0.8784905,0.94486535,1.0112402,1.0737107,1.3782539,1.678893,1.9834363,2.2840753,2.5886188,2.377781,2.1669433,1.9561055,1.7491722,1.5383345,1.3274968,1.116659,0.9058213,0.698888,0.48805028,0.63641757,0.78088045,0.92924774,1.077615,1.2259823,1.0073358,0.78868926,0.57394713,0.3553006,0.13665408,0.1639849,0.18741131,0.21083772,0.23816854,0.26159495,0.26940376,0.27721256,0.28502136,0.29283017,0.30063897,0.25378615,0.20693332,0.15617609,0.10932326,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.027330816,0.042948425,0.058566034,0.07418364,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.023426414,0.019522011,0.015617609,0.015617609,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.12103647,0.19131571,0.26159495,0.3318742,0.39824903,0.5270943,0.6559396,0.78088045,0.9097257,1.038571,0.8823949,0.7262188,0.57394713,0.41777104,0.26159495,0.21083772,0.15617609,0.10541886,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.08980125,0.093705654,0.093705654,0.09761006,0.10151446,0.14055848,0.1835069,0.22645533,0.26940376,0.31235218,0.28111696,0.25378615,0.22255093,0.19131571,0.1639849,0.19522011,0.22645533,0.26159495,0.29283017,0.3240654,0.29673457,0.26940376,0.24207294,0.21474212,0.18741131,0.7418364,1.2962615,1.8506867,2.4090161,2.9634414,3.8965936,4.83365,5.7668023,6.703859,7.6370106,9.093353,10.553599,12.009941,13.466284,14.92653,13.661504,12.400381,11.139259,9.874233,8.6131115,7.137247,5.661383,4.1894236,2.7135596,1.2376955,1.8116426,2.3816853,2.9556324,3.5256753,4.0996222,4.482254,4.8648853,5.2475166,5.630148,6.012779,6.969358,7.9259367,8.886419,9.8429985,10.799577,9.019169,7.238762,5.4583545,3.6818514,1.901444,1.7725986,1.6437533,1.5188124,1.3899672,1.261122,1.5461433,1.8272603,2.1083772,2.3933985,2.6745155,3.2484627,3.8185053,4.3924527,4.9663997,5.5364423,5.1616197,4.786797,4.4119744,4.037152,3.6623292,3.0610514,2.463678,1.8623998,1.261122,0.6637484,0.8394465,1.0190489,1.1947471,1.3743496,1.5500476,2.4714866,3.3890212,4.31046,5.2318993,6.1494336,5.6262436,5.099149,4.575959,4.0488653,3.5256753,2.9439192,2.358259,1.7765031,1.1947471,0.61299115,0.6715572,0.7340276,0.79259366,0.8511597,0.9136301,1.0580931,1.2064602,1.3548276,1.5031948,1.6515622,2.3153105,2.979059,3.6467118,4.31046,4.9742084,5.138193,5.298274,5.462259,5.6262436,5.786324,5.579391,5.368553,5.1577153,4.9468775,4.73604,6.98888,9.237816,11.486752,13.735687,15.988527,16.238409,16.492195,16.745981,16.995863,17.24965,14.329156,11.404759,8.484266,5.559869,2.639376,3.408543,4.181615,4.9546866,5.727758,6.5008297,6.3407493,6.180669,6.0205884,5.860508,5.700427,4.6657605,3.6349986,2.6042364,1.5695697,0.5388075,1.0854238,1.6320401,2.1786566,2.7291772,3.2757936,2.920493,2.5651922,2.2098918,1.8545911,1.4992905,1.261122,1.0190489,0.78088045,0.5388075,0.30063897,0.25378615,0.21083772,0.1639849,0.12103647,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7066968,1.4094892,2.1161861,2.8189783,3.5256753,3.1664703,2.803361,2.4441557,2.084951,1.7257458,1.6164225,1.5031948,1.3938715,1.2845483,1.175225,1.8467822,2.5183394,3.193801,3.8653584,4.5369153,3.6662338,2.7916477,1.9209659,1.0463798,0.1756981,0.1717937,0.1639849,0.16008049,0.15617609,0.14836729,0.18741131,0.22645533,0.26159495,0.30063897,0.3357786,0.3240654,0.31235218,0.30063897,0.28892577,0.27330816,0.3357786,0.39824903,0.46071947,0.5231899,0.58566034,0.46852827,0.3513962,0.23426414,0.11713207,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.06637484,0.05466163,0.046852827,0.03513962,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.1639849,0.25378615,0.3435874,0.43338865,0.5231899,0.5309987,0.5388075,0.5466163,0.5544251,0.5622339,0.61689556,0.6715572,0.7262188,0.78088045,0.8394465,1.0815194,1.3235924,1.5656652,1.8077383,2.0498111,1.9053483,1.7608855,1.6164225,1.4680552,1.3235924,1.1674163,1.0112402,0.8511597,0.6949836,0.5388075,0.6442264,0.75354964,0.8589685,0.96829176,1.0737107,0.9136301,0.75354964,0.59346914,0.43338865,0.27330816,0.30063897,0.3240654,0.3513962,0.37482262,0.39824903,0.42557985,0.45681506,0.48414588,0.5114767,0.5388075,0.45681506,0.3709182,0.28892577,0.20693332,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.05466163,0.08589685,0.113227665,0.14446288,0.1756981,0.14836729,0.12494087,0.10151446,0.07418364,0.05075723,0.046852827,0.039044023,0.03513962,0.031235218,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.1639849,0.23035973,0.29673457,0.359205,0.42557985,0.58175594,0.7340276,0.8902037,1.0463798,1.1986516,1.038571,0.8784905,0.71841,0.5583295,0.39824903,0.32016098,0.23816854,0.16008049,0.078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.1796025,0.1835069,0.19131571,0.19522011,0.19912452,0.21083772,0.21864653,0.23035973,0.23816854,0.24988174,0.26549935,0.28111696,0.29673457,0.30844778,0.3240654,0.3279698,0.3318742,0.3318742,0.3357786,0.3357786,0.3435874,0.3513962,0.359205,0.3670138,0.37482262,0.79649806,1.2181735,1.6437533,2.0654287,2.4871042,3.2094188,3.9278288,4.646239,5.368553,6.086963,7.152865,8.218767,9.280765,10.346666,11.412568,11.748346,12.08803,12.423808,12.763491,13.09927,10.674636,8.250002,5.825368,3.4007344,0.97610056,2.2450314,3.513962,4.786797,6.055728,7.3246584,7.3402762,7.355894,7.3715115,7.3832245,7.3988423,8.300759,9.20658,10.108498,11.010414,11.912332,10.22563,8.542832,6.8561306,5.173333,3.4866312,3.2562714,3.0259118,2.795552,2.5690966,2.338737,2.803361,3.2679846,3.7326086,4.1972322,4.661856,4.6930914,4.728231,4.759466,4.7907014,4.825841,4.4393053,4.0488653,3.6623292,3.2757936,2.8892577,2.4129205,1.9365835,1.4641509,0.9878138,0.5114767,0.6442264,0.77307165,0.9019169,1.0307622,1.1635119,1.9522011,2.7408905,3.533484,4.322173,5.1108627,5.3138914,5.5130157,5.7121406,5.911265,6.114294,4.997635,3.8809757,2.7682211,1.6515622,0.5388075,0.74574083,0.95267415,1.1596074,1.3665408,1.5734742,1.893635,2.2137961,2.533957,2.854118,3.174279,3.3187418,3.4593005,3.6037633,3.7443218,3.8887846,4.575959,5.263134,5.950309,6.6374836,7.3246584,7.2934237,7.2582836,7.2270484,7.195813,7.1606736,8.58578,10.010887,11.435994,12.861101,14.286208,14.329156,14.372105,14.415053,14.458001,14.50095,12.654168,10.81129,8.964508,7.1216297,5.2748475,6.79366,8.316377,9.835189,11.354002,12.8767185,12.568271,12.259823,11.951375,11.6468315,11.338385,9.2221985,7.1060123,4.9937305,2.8775444,0.76135844,1.9209659,3.076669,4.2362766,5.3919797,6.551587,5.840986,5.1303844,4.4197836,3.7091823,2.998581,2.5183394,2.0380979,1.5617609,1.0815194,0.60127795,0.5114767,0.42167544,0.3318742,0.23816854,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.46852827,0.94096094,1.4094892,1.8819219,2.35045,2.1239948,1.893635,1.6671798,1.4407244,1.2142692,1.3235924,1.4329157,1.542239,1.6515622,1.7608855,2.0146716,2.2684577,2.5183394,2.7721257,3.0259118,2.4714866,1.9209659,1.3665408,0.8160201,0.26159495,0.23035973,0.19912452,0.1639849,0.13274968,0.10151446,0.12494087,0.14836729,0.1756981,0.19912452,0.22645533,0.26159495,0.30063897,0.3357786,0.37482262,0.41386664,0.48805028,0.5622339,0.63641757,0.7106012,0.78868926,0.62860876,0.47243267,0.31625658,0.15617609,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.046852827,0.046852827,0.042948425,0.039044023,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.10932326,0.1717937,0.23035973,0.28892577,0.3513962,0.3553006,0.359205,0.3631094,0.3709182,0.37482262,0.42167544,0.46462387,0.5114767,0.5544251,0.60127795,0.78088045,0.96438736,1.1478943,1.3314011,1.5110037,1.4329157,1.3509232,1.2728351,1.1908426,1.1127546,1.0073358,0.9019169,0.79649806,0.6910792,0.58566034,0.6559396,0.7223144,0.78868926,0.8589685,0.92534333,0.8238289,0.71841,0.61689556,0.5153811,0.41386664,0.43729305,0.46071947,0.48805028,0.5114767,0.5388075,0.58566034,0.63251317,0.679366,0.7262188,0.77307165,0.6559396,0.5388075,0.42167544,0.30454338,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.08199245,0.12884527,0.1717937,0.21864653,0.26159495,0.22645533,0.18741131,0.14836729,0.113227665,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.21083772,0.26940376,0.3318742,0.39044023,0.44900626,0.63251317,0.8160201,0.9956226,1.1791295,1.3626363,1.1986516,1.0307622,0.8667773,0.7027924,0.5388075,0.42948425,0.3240654,0.21474212,0.10932326,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10541886,0.15617609,0.21083772,0.26159495,0.26940376,0.27721256,0.28502136,0.29283017,0.30063897,0.27721256,0.25378615,0.23426414,0.21083772,0.18741131,0.24597734,0.30844778,0.3670138,0.42557985,0.48805028,0.46071947,0.43338865,0.40605783,0.37872702,0.3513962,0.39434463,0.43338865,0.47633708,0.5192855,0.5622339,0.8511597,1.1439898,1.4329157,1.7218413,2.0107672,2.5183394,3.0220075,3.5256753,4.0332475,4.5369153,5.2084727,5.883934,6.5554914,7.2270484,7.898606,9.839094,11.775677,13.712261,15.648844,17.589333,14.212025,10.838621,7.461313,4.087909,0.7106012,2.67842,4.646239,6.6140575,8.581876,10.549695,10.198298,9.846903,9.491602,9.140205,8.78881,9.636065,10.48332,11.330575,12.177831,13.025085,11.435994,9.846903,8.253906,6.6648145,5.0757227,4.743849,4.40807,4.0761957,3.7443218,3.4124475,4.0605783,4.7087092,5.35684,6.001066,6.649197,6.141625,5.6340523,5.12648,4.618908,4.1113358,3.7130866,3.310933,2.912684,2.514435,2.1122816,1.7608855,1.4133936,1.0619974,0.7106012,0.3631094,0.44510186,0.5270943,0.60908675,0.6910792,0.77307165,1.43682,2.096664,2.7565079,3.416352,4.0761957,5.001539,5.9268827,6.8483214,7.773665,8.699008,7.0513506,5.4036927,3.7560349,2.1083772,0.46071947,0.8160201,1.1713207,1.5266213,1.8819219,2.2372224,2.7291772,3.2211318,3.7130866,4.2089458,4.7009,4.318269,3.9395418,3.5608149,3.1781836,2.7994564,4.0137253,5.22409,6.4383593,7.648724,8.862993,9.007456,9.151918,9.296382,9.440845,9.589212,10.186585,10.787864,11.389141,11.986515,12.587793,12.419904,12.252014,12.084125,11.916236,11.748346,10.983084,10.213917,9.448653,8.679486,7.914223,10.178777,12.447234,14.7156925,16.98415,19.248703,18.795792,18.338978,17.886066,17.429253,16.976341,13.778636,10.58093,7.3832245,4.185519,0.9878138,2.7565079,4.521298,6.289992,8.058686,9.823476,8.761478,7.6955767,6.629675,5.563773,4.5017757,3.7794614,3.0610514,2.338737,1.620327,0.9019169,0.76526284,0.62860876,0.4958591,0.359205,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23426414,0.46852827,0.7066968,0.94096094,1.175225,1.0815194,0.98390937,0.8902037,0.79649806,0.698888,1.0307622,1.358732,1.6906061,2.018576,2.35045,2.182561,2.0146716,1.8467822,1.678893,1.5110037,1.2806439,1.0463798,0.8160201,0.58175594,0.3513962,0.28892577,0.23035973,0.1717937,0.10932326,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.19912452,0.28892577,0.37482262,0.46071947,0.5505207,0.63641757,0.7262188,0.81211567,0.9019169,0.9878138,0.78868926,0.59346914,0.39434463,0.19912452,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.031235218,0.03513962,0.039044023,0.046852827,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.05466163,0.08589685,0.113227665,0.14446288,0.1756981,0.1756981,0.1796025,0.1835069,0.1835069,0.18741131,0.22255093,0.25769055,0.29283017,0.3279698,0.3631094,0.48414588,0.60908675,0.7301232,0.8511597,0.97610056,0.96048295,0.94486535,0.92924774,0.9136301,0.9019169,0.8472553,0.79649806,0.7418364,0.6910792,0.63641757,0.6637484,0.6910792,0.71841,0.74574083,0.77307165,0.7301232,0.6832704,0.64032197,0.59346914,0.5505207,0.57394713,0.60127795,0.62470436,0.6481308,0.6754616,0.7418364,0.80821127,0.8784905,0.94486535,1.0112402,0.8589685,0.7066968,0.5544251,0.40215343,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.10932326,0.1717937,0.23035973,0.28892577,0.3513962,0.30063897,0.24988174,0.19912452,0.14836729,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.25378615,0.30844778,0.3631094,0.42167544,0.47633708,0.6832704,0.8941081,1.1049459,1.3157835,1.5266213,1.3548276,1.1869383,1.0151446,0.8433509,0.6754616,0.5388075,0.40605783,0.26940376,0.13665408,0.0,0.0,0.0,0.0,0.0,0.0,0.07027924,0.14055848,0.21083772,0.28111696,0.3513962,0.359205,0.3709182,0.37872702,0.39044023,0.39824903,0.3435874,0.28892577,0.23426414,0.1796025,0.12494087,0.23035973,0.3357786,0.44119745,0.5466163,0.6481308,0.59346914,0.5349031,0.47633708,0.42167544,0.3631094,0.44119745,0.5192855,0.59346914,0.6715572,0.74964523,0.9058213,1.0659018,1.2220778,1.3782539,1.5383345,1.8272603,2.1161861,2.4090161,2.697942,2.9868677,3.2679846,3.5491016,3.8263142,4.1074314,4.388548,7.9259367,11.4633255,15.000713,18.538101,22.07549,17.749413,13.423335,9.101162,4.775084,0.44900626,3.1157131,5.7785153,8.445222,11.111929,13.774731,13.056321,12.334006,11.615597,10.893282,10.174872,10.967466,11.760059,12.552653,13.345247,14.13784,12.642454,11.147068,9.651682,8.156297,6.66091,6.2275214,5.794133,5.35684,4.9234514,4.4861584,5.3177958,6.1494336,6.9771667,7.8088045,8.636538,7.590158,6.5437784,5.493494,4.447114,3.4007344,2.9868677,2.5769055,2.1630387,1.7491722,1.33921,1.1127546,0.8862993,0.6637484,0.43729305,0.21083772,0.24597734,0.28111696,0.31625658,0.3513962,0.38653582,0.91753453,1.4485333,1.9756275,2.5066261,3.0376248,4.689187,6.336845,7.988407,9.636065,11.287627,9.108971,6.9264097,4.747753,2.5690966,0.38653582,0.8902037,1.3938715,1.893635,2.397303,2.900971,3.5647192,4.2284675,4.8961205,5.559869,6.223617,5.3217,4.4197836,3.5178664,2.6159496,1.7140326,3.4514916,5.1889505,6.9264097,8.663869,10.401327,10.721489,11.045554,11.365715,11.68978,12.013845,11.787391,11.560935,11.338385,11.111929,10.889378,10.510651,10.131924,9.753197,9.378374,8.999647,9.308095,9.620447,9.928895,10.241247,10.549695,13.563893,16.578093,19.596195,22.610394,25.624592,25.023314,24.422035,23.816854,23.215576,22.614298,18.33117,14.051944,9.772718,5.493494,1.2142692,3.59205,5.9659266,8.343708,10.721489,13.09927,11.678067,10.260769,8.839567,7.4183645,6.001066,5.040583,4.0801005,3.1196175,2.1591344,1.1986516,1.0190489,0.8394465,0.659844,0.48024148,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.737932,1.2884527,1.8389735,2.3855898,2.9361105,2.35045,1.7608855,1.175225,0.58566034,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.3513962,0.26159495,0.1756981,0.08589685,0.0,0.0,0.0,0.0,0.0,0.0,0.13665408,0.27330816,0.41386664,0.5505207,0.6871748,0.78868926,0.8862993,0.9878138,1.0893283,1.1869383,0.94876975,0.7106012,0.47633708,0.23816854,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.18741131,0.24988174,0.31235218,0.37482262,0.43729305,0.48805028,0.5388075,0.58566034,0.63641757,0.6871748,0.6871748,0.6871748,0.6871748,0.6871748,0.6871748,0.6754616,0.6637484,0.6481308,0.63641757,0.62470436,0.63641757,0.6481308,0.6637484,0.6754616,0.6871748,0.7106012,0.737932,0.76135844,0.78868926,0.81211567,0.9019169,0.9878138,1.0737107,1.1635119,1.2494087,1.0619974,0.8745861,0.6871748,0.4997635,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.13665408,0.21083772,0.28892577,0.3631094,0.43729305,0.37482262,0.31235218,0.24988174,0.18741131,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.30063897,0.3513962,0.39824903,0.44900626,0.4997635,0.737932,0.97610056,1.2142692,1.4485333,1.6867018,1.5110037,1.33921,1.1635119,0.9878138,0.81211567,0.6481308,0.48805028,0.3240654,0.1639849,0.0,0.0,0.0,0.0,0.0,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.44900626,0.46071947,0.47633708,0.48805028,0.4997635,0.41386664,0.3240654,0.23816854,0.14836729,0.062470436,0.21083772,0.3631094,0.5114767,0.6637484,0.81211567,0.7262188,0.63641757,0.5505207,0.46071947,0.37482262,0.48805028,0.60127795,0.7106012,0.8238289,0.93705654,0.96438736,0.9878138,1.0112402,1.038571,1.0619974,1.1361811,1.2142692,1.2884527,1.3626363,1.43682,1.3235924,1.2142692,1.1010414,0.9878138,0.8745861,6.012779,11.150972,16.289165,21.423454,26.56165,21.2868,16.011953,10.737106,5.462259,0.18741131,3.5491016,6.910792,10.276386,13.638077,16.999767,15.914344,14.825015,13.735687,12.650263,11.560935,12.298867,13.036799,13.774731,14.512663,15.250595,13.848915,12.4511385,11.0494585,9.651682,8.250002,7.7111945,7.1762915,6.6374836,6.098676,5.563773,6.575013,7.5862536,8.601398,9.612638,10.6238785,9.0386915,7.4495993,5.860508,4.2753205,2.6862288,2.260649,1.8389735,1.4133936,0.9878138,0.5622339,0.46071947,0.3631094,0.26159495,0.1639849,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.39824903,0.80040246,1.1986516,1.6008049,1.999054,4.376835,6.7507114,9.124588,11.498465,13.8762455,11.162686,8.449126,5.735567,3.0259118,0.31235218,0.96438736,1.6125181,2.260649,2.912684,3.5608149,4.4002614,5.2358036,6.0752497,6.910792,7.7502384,6.3251314,4.900025,3.474918,2.0498111,0.62470436,2.8892577,5.1499066,7.4144597,9.675109,11.935758,12.439425,12.939189,13.438952,13.938716,14.438479,13.388195,12.337912,11.287627,10.237343,9.187058,8.601398,8.011833,7.426173,6.8366084,6.250948,7.6370106,9.023073,10.413041,11.799104,13.189071,16.94901,20.712854,24.476698,28.236637,32.00048,31.250835,30.50119,29.751545,29.0019,28.24835,22.887606,17.526861,12.162213,6.801469,1.43682,4.423688,7.4105554,10.401327,13.388195,16.375063,14.59856,12.825961,11.0494585,9.276859,7.5003567,6.3017054,5.099149,3.900498,2.7018464,1.4992905,1.2767396,1.0502841,0.8238289,0.60127795,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.58956474,1.0307622,1.4680552,1.9092526,2.35045,1.8819219,1.4094892,0.94096094,0.46852827,0.0,0.07027924,0.14055848,0.21083772,0.28111696,0.3513962,0.28111696,0.21083772,0.14055848,0.07027924,0.0,0.0,0.0,0.0,0.0,0.0,0.10932326,0.21864653,0.3318742,0.44119745,0.5505207,0.62860876,0.7106012,0.78868926,0.8706817,0.94876975,0.76135844,0.5700427,0.37872702,0.19131571,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.10151446,0.1678893,0.23426414,0.29673457,0.3631094,0.28892577,0.21864653,0.14446288,0.07418364,0.0,0.046852827,0.093705654,0.14055848,0.19131571,0.23816854,0.27330816,0.31235218,0.3513962,0.38653582,0.42557985,0.339683,0.25378615,0.1717937,0.08589685,0.0,0.0,0.0,0.0,0.0,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.12884527,0.12103647,0.113227665,0.10932326,0.10151446,0.08199245,0.06637484,0.046852827,0.031235218,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.15227169,0.20693332,0.25769055,0.30844778,0.3631094,0.40996224,0.45681506,0.5036679,0.5544251,0.60127795,0.60518235,0.60908675,0.61689556,0.62079996,0.62470436,0.62079996,0.62079996,0.61689556,0.61689556,0.61299115,0.62079996,0.63251317,0.6442264,0.6520352,0.6637484,0.6910792,0.71841,0.74574083,0.77307165,0.80040246,0.8589685,0.9136301,0.97219616,1.0307622,1.0893283,0.96438736,0.8433509,0.71841,0.59737355,0.47633708,0.38653582,0.29673457,0.20693332,0.113227665,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.10932326,0.1717937,0.23035973,0.28892577,0.3513962,0.30063897,0.24988174,0.19912452,0.14836729,0.10151446,0.12103647,0.14446288,0.1678893,0.19131571,0.21083772,0.19131571,0.1717937,0.15227169,0.13274968,0.113227665,0.10932326,0.10932326,0.10541886,0.10151446,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.058566034,0.10932326,0.15617609,0.20302892,0.24988174,0.29673457,0.3435874,0.39434463,0.44119745,0.48805028,0.679366,0.8667773,1.0580931,1.2494087,1.43682,1.33921,1.2415999,1.1439898,1.0463798,0.94876975,0.8160201,0.6832704,0.5544251,0.42167544,0.28892577,0.24597734,0.20693332,0.1678893,0.12884527,0.08589685,0.14836729,0.20693332,0.26940376,0.3279698,0.38653582,0.42948425,0.47243267,0.5153811,0.5583295,0.60127795,0.4958591,0.39044023,0.28502136,0.1796025,0.07418364,0.19912452,0.32016098,0.44119745,0.5661383,0.6871748,0.61689556,0.5427119,0.46852827,0.39824903,0.3240654,0.41386664,0.5036679,0.59346914,0.6832704,0.77307165,0.78868926,0.80430686,0.8199245,0.8355421,0.8511597,0.93705654,1.0268579,1.1127546,1.1986516,1.2884527,1.1791295,1.0737107,0.96438736,0.8589685,0.74964523,5.0640097,9.37447,13.688834,17.999294,22.31366,17.96025,13.610746,9.261242,4.911738,0.5622339,3.1859922,5.813655,8.437413,11.061172,13.688834,12.802535,11.916236,11.033841,10.147541,9.261242,9.86252,10.4637985,11.061172,11.66245,12.263727,11.143164,10.0265045,8.909846,7.793187,6.676528,6.2314262,5.786324,5.3412223,4.8961205,4.4510183,5.3217,6.196286,7.066968,7.941554,8.812236,7.5081654,6.2040954,4.8961205,3.59205,2.2879796,1.9209659,1.5539521,1.183034,0.8160201,0.44900626,0.3709182,0.28892577,0.21083772,0.12884527,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.32016098,0.64032197,0.96048295,1.2806439,1.6008049,3.513962,5.423215,7.336372,9.249529,11.162686,9.190963,7.2192397,5.2436123,3.2718892,1.3001659,1.756981,2.2137961,2.6706111,3.1313305,3.5881457,4.181615,4.7711797,5.364649,5.958118,6.551587,5.7316628,4.9156423,4.095718,3.279698,2.463678,4.5837684,6.703859,8.823949,10.944039,13.06413,12.911859,12.763491,12.611219,12.4628525,12.31058,11.326671,10.342762,9.358852,8.371038,7.387129,7.164578,6.942027,6.719476,6.4969254,6.2743745,7.1606736,8.050878,8.937177,9.823476,10.71368,14.087084,17.456583,20.829987,24.20339,27.576794,26.90914,26.245392,25.581644,24.91399,24.250242,20.705046,17.159847,13.614651,10.069453,6.524256,8.32809,10.131924,11.931853,13.735687,15.535617,13.735687,11.935758,10.135828,8.335898,6.5359693,5.4856853,4.4314966,3.3812122,2.3270237,1.2767396,1.1322767,0.9917182,0.8472553,0.7066968,0.5622339,0.6832704,0.80821127,0.92924774,1.0541886,1.175225,0.96829176,0.76526284,0.5583295,0.3553006,0.14836729,0.12884527,0.10932326,0.08980125,0.07027924,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.44119745,0.77307165,1.1010414,1.4329157,1.7608855,1.4094892,1.0580931,0.7066968,0.3513962,0.0,0.05075723,0.10541886,0.15617609,0.21083772,0.26159495,0.21083772,0.15617609,0.10541886,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.08199245,0.1639849,0.24597734,0.3318742,0.41386664,0.47243267,0.5309987,0.59346914,0.6520352,0.7106012,0.5700427,0.42557985,0.28502136,0.14055848,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.19131571,0.30844778,0.42557985,0.5466163,0.6637484,0.5309987,0.39824903,0.26549935,0.13274968,0.0,0.093705654,0.19131571,0.28502136,0.37872702,0.47633708,0.5505207,0.62470436,0.698888,0.77307165,0.8511597,0.679366,0.5114767,0.339683,0.1717937,0.0,0.0,0.0,0.0,0.0,0.0,0.05466163,0.10932326,0.1639849,0.21864653,0.27330816,0.26159495,0.24597734,0.23035973,0.21474212,0.19912452,0.1639849,0.12884527,0.093705654,0.058566034,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.11713207,0.16008049,0.20302892,0.24597734,0.28892577,0.3318742,0.37872702,0.42167544,0.46852827,0.5114767,0.5231899,0.5309987,0.5427119,0.5544251,0.5622339,0.5700427,0.57785153,0.58566034,0.59346914,0.60127795,0.60908675,0.61689556,0.62079996,0.62860876,0.63641757,0.6676528,0.698888,0.7262188,0.75745404,0.78868926,0.8160201,0.8433509,0.8706817,0.8980125,0.92534333,0.8667773,0.80821127,0.75354964,0.6949836,0.63641757,0.5192855,0.40215343,0.28502136,0.1678893,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.08199245,0.12884527,0.1717937,0.21864653,0.26159495,0.22645533,0.18741131,0.14836729,0.113227665,0.07418364,0.13274968,0.19131571,0.24597734,0.30454338,0.3631094,0.3240654,0.28111696,0.24207294,0.20302892,0.1639849,0.1717937,0.1756981,0.1835069,0.19131571,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.07027924,0.113227665,0.16008049,0.20693332,0.24988174,0.29673457,0.339683,0.38653582,0.42948425,0.47633708,0.61689556,0.76135844,0.9019169,1.0463798,1.1869383,1.1674163,1.1478943,1.1283722,1.1088502,1.0893283,0.98390937,0.8823949,0.78088045,0.679366,0.57394713,0.4958591,0.41386664,0.3357786,0.25378615,0.1756981,0.20693332,0.23816854,0.27330816,0.30454338,0.3357786,0.40996224,0.48414588,0.5544251,0.62860876,0.698888,0.57785153,0.45681506,0.3318742,0.21083772,0.08589685,0.1835069,0.27721256,0.3709182,0.46852827,0.5622339,0.5036679,0.44900626,0.39044023,0.3318742,0.27330816,0.3435874,0.40996224,0.47633708,0.5466163,0.61299115,0.61689556,0.62079996,0.62860876,0.63251317,0.63641757,0.737932,0.8394465,0.93705654,1.038571,1.1361811,1.0346665,0.93315214,0.8316377,0.7262188,0.62470436,4.1113358,7.5979667,11.088503,14.575133,18.061766,14.637604,11.213444,7.7892823,4.3612175,0.93705654,2.8267872,4.7126136,6.5984397,8.488171,10.373997,9.690726,9.01136,8.32809,7.6448197,6.9615493,7.426173,7.8868923,8.351517,8.812236,9.276859,8.441318,7.605776,6.7702336,5.9346914,5.099149,4.747753,4.396357,4.041056,3.68966,3.338264,4.068387,4.802415,5.5364423,6.266566,7.000593,5.9776397,4.9546866,3.9317331,2.9087796,1.8858263,1.5773785,1.2689307,0.95657855,0.6481308,0.3357786,0.27721256,0.21864653,0.15617609,0.09761006,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.23816854,0.48024148,0.71841,0.96048295,1.1986516,2.6510892,4.0996222,5.548156,7.000593,8.449126,7.2192397,5.985449,4.7516575,3.521771,2.2879796,2.5534792,2.8189783,3.0805733,3.3460727,3.611572,3.959064,4.3065557,4.6540475,5.001539,5.349031,5.138193,4.93126,4.7204223,4.5095844,4.298747,6.278279,8.253906,10.2334385,12.209065,14.188598,13.388195,12.587793,11.787391,10.986988,10.186585,9.269051,8.347612,7.426173,6.5086384,5.5871997,5.7316628,5.872221,6.016684,6.1572423,6.3017054,6.688241,7.0747766,7.461313,7.8517528,8.238289,11.221252,14.204215,17.183275,20.166237,23.1492,22.57135,21.989594,21.411741,20.829987,20.24823,18.522484,16.796738,15.067088,13.341343,11.611692,12.228588,12.849388,13.466284,14.0831785,14.700074,12.8767185,11.0494585,9.226103,7.3988423,5.575486,4.6696653,3.7638438,2.8580225,1.9561055,1.0502841,0.9917182,0.92924774,0.8706817,0.80821127,0.74964523,1.0698062,1.3899672,1.7101282,2.0302892,2.35045,1.9404879,1.5305257,1.1205635,0.7106012,0.30063897,0.26159495,0.21864653,0.1796025,0.14055848,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.29673457,0.5153811,0.7340276,0.95657855,1.175225,0.94096094,0.7066968,0.46852827,0.23426414,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.0,0.0,0.0,0.0,0.0,0.05466163,0.10932326,0.1639849,0.21864653,0.27330816,0.31625658,0.3553006,0.39434463,0.43338865,0.47633708,0.37872702,0.28502136,0.19131571,0.093705654,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.28111696,0.45291066,0.62079996,0.79259366,0.96438736,0.76916724,0.57785153,0.38653582,0.19131571,0.0,0.14055848,0.28502136,0.42557985,0.5700427,0.7106012,0.8238289,0.93705654,1.0502841,1.1635119,1.2767396,1.0190489,0.76526284,0.5114767,0.25378615,0.0,0.0,0.0,0.0,0.0,0.0,0.08199245,0.1639849,0.24597734,0.3318742,0.41386664,0.39044023,0.3670138,0.3435874,0.3240654,0.30063897,0.24597734,0.19522011,0.14055848,0.08980125,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.08199245,0.113227665,0.14836729,0.1796025,0.21083772,0.25378615,0.29673457,0.339683,0.38263142,0.42557985,0.44119745,0.45681506,0.46852827,0.48414588,0.4997635,0.5192855,0.5349031,0.5544251,0.5700427,0.58566034,0.59346914,0.59737355,0.60127795,0.60908675,0.61299115,0.6442264,0.679366,0.7106012,0.7418364,0.77307165,0.77307165,0.76916724,0.76916724,0.76526284,0.76135844,0.76916724,0.77697605,0.78478485,0.79259366,0.80040246,0.6559396,0.5114767,0.3631094,0.21864653,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.05466163,0.08589685,0.113227665,0.14446288,0.1756981,0.14836729,0.12494087,0.10151446,0.07418364,0.05075723,0.14055848,0.23426414,0.3279698,0.42167544,0.5114767,0.45291066,0.39434463,0.3318742,0.27330816,0.21083772,0.23035973,0.24597734,0.26549935,0.28111696,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.078088045,0.12103647,0.1639849,0.20693332,0.24988174,0.29283017,0.3357786,0.37872702,0.42167544,0.46071947,0.5583295,0.6520352,0.74574083,0.8433509,0.93705654,0.9956226,1.0541886,1.1088502,1.1674163,1.2259823,1.1517987,1.0815194,1.0073358,0.93315214,0.8628729,0.7418364,0.62079996,0.5036679,0.38263142,0.26159495,0.26940376,0.27330816,0.27721256,0.28111696,0.28892577,0.39044023,0.49195468,0.59346914,0.698888,0.80040246,0.659844,0.5192855,0.37872702,0.23816854,0.10151446,0.1678893,0.23426414,0.30063897,0.3709182,0.43729305,0.39434463,0.3513962,0.30844778,0.26940376,0.22645533,0.26940376,0.31625658,0.359205,0.40605783,0.44900626,0.44510186,0.44119745,0.43338865,0.42948425,0.42557985,0.5388075,0.6481308,0.76135844,0.8745861,0.9878138,0.8902037,0.79259366,0.6949836,0.59737355,0.4997635,3.1625657,5.825368,8.488171,11.150972,13.813775,11.311053,8.812236,6.3134184,3.8106966,1.3118792,2.463678,3.611572,4.7633705,5.911265,7.0630636,6.5828223,6.1025805,5.6223392,5.142098,4.661856,4.985922,5.3138914,5.6379566,5.9620223,6.2860875,5.735567,5.181142,4.630621,4.0761957,3.5256753,3.2640803,3.0063896,2.7447948,2.4831998,2.2255092,2.8189783,3.408543,4.0020123,4.5954814,5.1889505,4.447114,3.7091823,2.9673457,2.2294137,1.4875772,1.2337911,0.98390937,0.7301232,0.47633708,0.22645533,0.1835069,0.14446288,0.10541886,0.06637484,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.16008049,0.32016098,0.48024148,0.64032197,0.80040246,1.7882162,2.77603,3.7638438,4.7516575,5.7394714,5.2436123,4.7516575,4.2597027,3.767748,3.2757936,3.3460727,3.4202564,3.49444,3.5647192,3.638903,3.7404175,3.8419318,3.9434462,4.0488653,4.1503797,4.548629,4.9468775,5.3412223,5.7394714,6.13772,7.9727893,9.807858,11.642927,13.477997,15.313066,13.860628,12.412095,10.963562,9.511124,8.062591,7.2075267,6.3524623,5.4973984,4.6423345,3.78727,4.2948427,4.802415,5.309987,5.8175592,6.3251314,6.211904,6.098676,5.989353,5.8761253,5.7628975,8.355421,10.947944,13.540467,16.13299,18.725513,18.229654,17.733795,17.24184,16.745981,16.250122,16.339924,16.429726,16.519526,16.609327,16.69913,16.13299,15.566852,14.996809,14.430671,13.860628,12.013845,10.163159,8.312472,6.461786,4.6110992,3.853645,3.096191,2.338737,1.5812829,0.8238289,0.8472553,0.8706817,0.8941081,0.9136301,0.93705654,1.456342,1.9717231,2.4910088,3.0063896,3.5256753,2.9087796,2.2957885,1.678893,1.0659018,0.44900626,0.39044023,0.3318742,0.26940376,0.21083772,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.14836729,0.25769055,0.3670138,0.47633708,0.58566034,0.46852827,0.3513962,0.23426414,0.11713207,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.15617609,0.1756981,0.19912452,0.21864653,0.23816854,0.19131571,0.14055848,0.093705654,0.046852827,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.3709182,0.59346914,0.8160201,1.038571,1.261122,1.0112402,0.75745404,0.5036679,0.25378615,0.0,0.19131571,0.37872702,0.5700427,0.76135844,0.94876975,1.1010414,1.2494087,1.4016805,1.5500476,1.698415,1.358732,1.0190489,0.679366,0.339683,0.0,0.0,0.0,0.0,0.0,0.0,0.10932326,0.21864653,0.3318742,0.44119745,0.5505207,0.5192855,0.49195468,0.46071947,0.42948425,0.39824903,0.3318742,0.26159495,0.19131571,0.12103647,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.046852827,0.07027924,0.093705654,0.113227665,0.13665408,0.1756981,0.21864653,0.25769055,0.29673457,0.3357786,0.359205,0.37872702,0.39824903,0.41777104,0.43729305,0.46462387,0.49195468,0.5192855,0.5466163,0.57394713,0.57785153,0.58175594,0.58175594,0.58566034,0.58566034,0.62079996,0.6559396,0.6910792,0.7262188,0.76135844,0.7301232,0.698888,0.6637484,0.63251317,0.60127795,0.6715572,0.74574083,0.8160201,0.8902037,0.96438736,0.78868926,0.61689556,0.44510186,0.27330816,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.027330816,0.042948425,0.058566034,0.07418364,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.15227169,0.28111696,0.40605783,0.5349031,0.6637484,0.58175594,0.5036679,0.42167544,0.3435874,0.26159495,0.28892577,0.31625658,0.3435874,0.3709182,0.39824903,0.32016098,0.23816854,0.16008049,0.078088045,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.08980125,0.12884527,0.1717937,0.21083772,0.24988174,0.28892577,0.3318742,0.3709182,0.40996224,0.44900626,0.4958591,0.5466163,0.59346914,0.64032197,0.6871748,0.8238289,0.95657855,1.0932326,1.2259823,1.3626363,1.319688,1.2767396,1.2337911,1.1908426,1.1517987,0.9917182,0.8316377,0.6715572,0.5114767,0.3513962,0.3279698,0.30454338,0.28111696,0.26159495,0.23816854,0.3709182,0.5036679,0.63641757,0.76916724,0.9019169,0.7418364,0.58566034,0.42557985,0.26940376,0.113227665,0.15227169,0.19131571,0.23426414,0.27330816,0.31235218,0.28502136,0.25769055,0.23035973,0.20302892,0.1756981,0.19912452,0.21864653,0.24207294,0.26549935,0.28892577,0.27330816,0.25769055,0.24207294,0.22645533,0.21083772,0.3357786,0.46071947,0.58566034,0.7106012,0.8394465,0.74574083,0.6520352,0.5583295,0.46852827,0.37482262,2.2137961,4.0488653,5.8878384,7.726812,9.561881,7.988407,6.4110284,4.8375545,3.2640803,1.6867018,2.1005683,2.5105307,2.9243972,3.338264,3.7482262,3.4710135,3.193801,2.9165885,2.639376,2.3621633,2.5495746,2.736986,2.9243972,3.1118085,3.2992198,3.0298162,2.7604125,2.4910088,2.2216048,1.9482968,1.7843118,1.6164225,1.4485333,1.2806439,1.1127546,1.5656652,2.018576,2.4714866,2.9243972,3.3734035,2.9165885,2.4597735,2.0029583,1.5461433,1.0893283,0.8941081,0.698888,0.5036679,0.30844778,0.113227665,0.093705654,0.07418364,0.05075723,0.031235218,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,0.92534333,1.4485333,1.9756275,2.4988174,3.0259118,3.2718892,3.521771,3.767748,4.0137253,4.263607,4.142571,4.0215344,3.9044023,3.7833657,3.6623292,3.521771,3.377308,3.2367494,3.0922866,2.951728,3.9551594,4.958591,5.9659266,6.969358,7.9766936,9.6673,11.361811,13.052417,14.746927,16.437534,14.336966,12.236397,10.135828,8.039165,5.938596,5.1460023,4.357313,3.5686235,2.77603,1.9873407,2.8619268,3.7326086,4.60329,5.477876,6.348558,5.735567,5.12648,4.513489,3.900498,3.2875066,5.4895897,7.6916723,9.893755,12.095839,14.301826,13.887959,13.477997,13.068034,12.658072,12.24811,14.157363,16.066616,17.971964,19.881216,21.786564,20.033487,18.284315,16.531239,14.778163,13.025085,11.150972,9.276859,7.3988423,5.5247293,3.6506162,3.0415294,2.4285383,1.8194515,1.2103647,0.60127795,0.7066968,0.80821127,0.9136301,1.0190489,1.1244678,1.8389735,2.5534792,3.2718892,3.9863946,4.7009,3.8809757,3.0610514,2.241127,1.4212024,0.60127795,0.5192855,0.44119745,0.359205,0.28111696,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.46071947,0.737932,1.0112402,1.2884527,1.5617609,1.2494087,0.93705654,0.62470436,0.31235218,0.0,0.23816854,0.47633708,0.7106012,0.94876975,1.1869383,1.3743496,1.5617609,1.7491722,1.9365835,2.1239948,1.698415,1.2767396,0.8511597,0.42557985,0.0,0.0,0.0,0.0,0.0,0.0,0.13665408,0.27330816,0.41386664,0.5505207,0.6871748,0.6481308,0.61299115,0.57394713,0.5388075,0.4997635,0.41386664,0.3240654,0.23816854,0.14836729,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.10151446,0.13665408,0.1756981,0.21083772,0.24988174,0.27330816,0.30063897,0.3240654,0.3513962,0.37482262,0.41386664,0.44900626,0.48805028,0.5231899,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.60127795,0.63641757,0.6754616,0.7106012,0.74964523,0.6871748,0.62470436,0.5622339,0.4997635,0.43729305,0.57394713,0.7106012,0.8511597,0.9878138,1.1244678,0.92534333,0.7262188,0.5231899,0.3240654,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1639849,0.3240654,0.48805028,0.6481308,0.81211567,0.7106012,0.61299115,0.5114767,0.41386664,0.31235218,0.3513962,0.38653582,0.42557985,0.46071947,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.10151446,0.13665408,0.1756981,0.21083772,0.24988174,0.28892577,0.3240654,0.3631094,0.39824903,0.43729305,0.43729305,0.43729305,0.43729305,0.43729305,0.43729305,0.6481308,0.8628729,1.0737107,1.2884527,1.4992905,1.4875772,1.475864,1.4641509,1.4485333,1.43682,1.2376955,1.038571,0.8355421,0.63641757,0.43729305,0.38653582,0.3357786,0.28892577,0.23816854,0.18741131,0.3513962,0.5114767,0.6754616,0.8394465,0.999527,0.8238289,0.6481308,0.47633708,0.30063897,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.13665408,0.27330816,0.41386664,0.5505207,0.6871748,0.60127795,0.5114767,0.42557985,0.3357786,0.24988174,1.261122,2.2762666,3.2875066,4.298747,5.3138914,4.661856,4.0137253,3.3616903,2.7135596,2.0615244,1.737459,1.4133936,1.0893283,0.76135844,0.43729305,0.3631094,0.28892577,0.21083772,0.13665408,0.062470436,0.113227665,0.1639849,0.21083772,0.26159495,0.31235218,0.3240654,0.3357786,0.3513962,0.3631094,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.31235218,0.62470436,0.93705654,1.2494087,1.5617609,1.3860629,1.2142692,1.038571,0.8628729,0.6871748,0.5505207,0.41386664,0.27330816,0.13665408,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,1.3001659,2.2879796,3.2757936,4.263607,5.251421,4.939069,4.6267166,4.3143644,3.998108,3.6857557,3.2992198,2.912684,2.5261483,2.135708,1.7491722,3.3616903,4.9742084,6.5867267,8.1992445,9.811763,11.361811,12.911859,14.461906,16.011953,17.562002,14.813302,12.0606985,9.311999,6.5633,3.8106966,3.0883822,2.3621633,1.6359446,0.9136301,0.18741131,1.4251068,2.6628022,3.900498,5.138193,6.375889,5.263134,4.1503797,3.0376248,1.9248703,0.81211567,2.6237583,4.4393053,6.250948,8.062591,9.874233,9.550168,9.226103,8.898132,8.574067,8.250002,11.974802,15.699601,19.4244,23.1492,26.874,23.937891,21.00178,18.061766,15.125654,12.185639,10.2881,8.386656,6.4891167,4.5876727,2.6862288,2.2255092,1.7608855,1.3001659,0.8394465,0.37482262,0.5622339,0.74964523,0.93705654,1.1244678,1.3118792,2.2255092,3.1391394,4.0488653,4.9624953,5.8761253,4.8492675,3.8263142,2.7994564,1.7765031,0.74964523,0.6481308,0.5505207,0.44900626,0.3513962,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.37872702,0.60518235,0.8316377,1.0580931,1.2884527,1.1010414,0.91753453,0.7340276,0.5466163,0.3631094,0.679366,0.9917182,1.3079748,1.6242313,1.9365835,1.8897307,1.8428779,1.796025,1.7491722,1.698415,1.358732,1.0190489,0.679366,0.339683,0.0,0.0,0.0,0.0,0.0,0.0,0.10932326,0.21864653,0.3318742,0.44119745,0.5505207,0.59346914,0.64032197,0.6832704,0.7301232,0.77307165,0.7262188,0.6754616,0.62470436,0.57394713,0.5231899,0.43338865,0.339683,0.24597734,0.15617609,0.062470436,0.05466163,0.046852827,0.039044023,0.031235218,0.023426414,0.023426414,0.019522011,0.015617609,0.015617609,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.08199245,0.113227665,0.14836729,0.1796025,0.21083772,0.23426414,0.25378615,0.27330816,0.29283017,0.31235218,0.339683,0.3670138,0.39434463,0.42167544,0.44900626,0.45291066,0.45681506,0.45681506,0.46071947,0.46071947,0.48805028,0.5192855,0.5466163,0.57394713,0.60127795,0.5700427,0.5388075,0.5114767,0.48024148,0.44900626,0.5583295,0.6637484,0.77307165,0.8784905,0.9878138,0.81211567,0.63641757,0.46071947,0.28892577,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.24988174,0.3240654,0.39824903,0.47633708,0.5505207,0.45681506,0.3631094,0.27330816,0.1796025,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13274968,0.26549935,0.39824903,0.5309987,0.6637484,0.60127795,0.5388075,0.47633708,0.41386664,0.3513962,0.38653582,0.42557985,0.46071947,0.4997635,0.5388075,0.44119745,0.3474918,0.25378615,0.15617609,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.093705654,0.12103647,0.15227169,0.1835069,0.21083772,0.24207294,0.27330816,0.30063897,0.3318742,0.3631094,0.3631094,0.3670138,0.3709182,0.3709182,0.37482262,0.5505207,0.7262188,0.9019169,1.0737107,1.2494087,1.2806439,1.3118792,1.33921,1.3704453,1.4016805,1.2337911,1.0659018,0.8980125,0.7301232,0.5622339,0.5075723,0.45291066,0.39824903,0.3435874,0.28892577,0.39434463,0.4958591,0.60127795,0.7066968,0.81211567,0.6949836,0.57785153,0.46071947,0.3435874,0.22645533,0.22255093,0.21864653,0.21864653,0.21474212,0.21083772,0.19131571,0.1678893,0.14446288,0.12103647,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.10932326,0.21864653,0.3318742,0.44119745,0.5505207,0.48414588,0.41386664,0.3474918,0.28111696,0.21083772,1.0268579,1.8428779,2.6588979,3.4710135,4.2870336,3.8106966,3.3343596,2.854118,2.377781,1.901444,1.6125181,1.3235924,1.038571,0.74964523,0.46071947,0.38653582,0.31235218,0.23816854,0.1639849,0.08589685,0.15617609,0.22645533,0.29673457,0.3670138,0.43729305,0.41386664,0.38653582,0.3631094,0.3357786,0.31235218,0.25378615,0.19131571,0.13274968,0.07418364,0.011713207,0.26159495,0.5075723,0.75354964,1.0034313,1.2494087,1.1088502,0.96829176,0.8316377,0.6910792,0.5505207,0.44119745,0.3318742,0.21864653,0.10932326,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,1.038571,1.8311646,2.619854,3.408543,4.2011366,3.978586,3.7560349,3.533484,3.310933,3.0883822,2.8970666,2.7057507,2.5183394,2.3270237,2.135708,3.4827268,4.825841,6.17286,7.5159745,8.862993,10.198298,11.537509,12.8767185,14.212025,15.551234,13.329629,11.111929,8.890324,6.6687193,4.4510183,3.9161155,3.3812122,2.8463092,2.3114061,1.7765031,2.7643168,3.7482262,4.73604,5.7238536,6.7116675,5.6809053,4.6540475,3.6232853,2.592523,1.5617609,2.8892577,4.2167544,5.5442514,6.871748,8.1992445,7.929841,7.660437,7.3910336,7.1216297,6.8483214,10.069453,13.2905855,16.511717,19.728945,22.950077,20.31851,17.686943,15.051471,12.419904,9.788337,9.347139,8.905942,8.468649,8.027451,7.5862536,6.211904,4.8375545,3.4632049,2.0888553,0.7106012,0.92924774,1.1478943,1.3665408,1.5812829,1.7999294,2.7252727,3.6506162,4.575959,5.5013027,6.426646,5.6926184,4.958591,4.2284675,3.49444,2.7643168,2.7291772,2.6940374,2.6588979,2.6237583,2.5886188,2.182561,1.7765031,1.3743496,0.96829176,0.5622339,0.46071947,0.3631094,0.26159495,0.1639849,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.29283017,0.47243267,0.6520352,0.8316377,1.0112402,0.95657855,0.8980125,0.8394465,0.78088045,0.7262188,1.116659,1.5110037,1.901444,2.2957885,2.6862288,2.4051118,2.1239948,1.8389735,1.5578566,1.2767396,1.0190489,0.76526284,0.5114767,0.25378615,0.0,0.0,0.0,0.0,0.0,0.0,0.08199245,0.1639849,0.24597734,0.3318742,0.41386664,0.5388075,0.6676528,0.79649806,0.92143893,1.0502841,1.038571,1.0268579,1.0112402,0.999527,0.9878138,0.8160201,0.6442264,0.46852827,0.29673457,0.12494087,0.10932326,0.093705654,0.078088045,0.06637484,0.05075723,0.046852827,0.039044023,0.03513962,0.031235218,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.06637484,0.093705654,0.12103647,0.14836729,0.1756981,0.19131571,0.20693332,0.21864653,0.23426414,0.24988174,0.26940376,0.28502136,0.30063897,0.32016098,0.3357786,0.3435874,0.3474918,0.3513962,0.359205,0.3631094,0.37872702,0.39824903,0.41386664,0.43338865,0.44900626,0.45291066,0.45681506,0.45681506,0.46071947,0.46071947,0.5388075,0.61689556,0.6949836,0.77307165,0.8511597,0.698888,0.5505207,0.39824903,0.24988174,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.07027924,0.14055848,0.21083772,0.28111696,0.3513962,0.4997635,0.6481308,0.80040246,0.94876975,1.1010414,0.9136301,0.7301232,0.5466163,0.359205,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.20693332,0.30844778,0.40996224,0.5114767,0.48805028,0.46071947,0.43729305,0.41386664,0.38653582,0.42557985,0.46071947,0.4997635,0.5388075,0.57394713,0.48414588,0.39434463,0.30454338,0.21474212,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.08589685,0.10932326,0.12884527,0.15227169,0.1756981,0.19912452,0.21864653,0.24207294,0.26549935,0.28892577,0.29283017,0.29673457,0.30063897,0.30844778,0.31235218,0.44900626,0.58566034,0.7262188,0.8628729,0.999527,1.0737107,1.1439898,1.2181735,1.2884527,1.3626363,1.2259823,1.0932326,0.95657855,0.8238289,0.6871748,0.62860876,0.5661383,0.5075723,0.44900626,0.38653582,0.43338865,0.48414588,0.5309987,0.57785153,0.62470436,0.5661383,0.5036679,0.44510186,0.38653582,0.3240654,0.30844778,0.28892577,0.27330816,0.25378615,0.23816854,0.20693332,0.1717937,0.14055848,0.10932326,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.08199245,0.1639849,0.24597734,0.3318742,0.41386664,0.3631094,0.31625658,0.26940376,0.22255093,0.1756981,0.79259366,1.4094892,2.0263848,2.6432803,3.2640803,2.9556324,2.6510892,2.3465457,2.0420024,1.737459,1.4875772,1.2376955,0.9878138,0.737932,0.48805028,0.41386664,0.3357786,0.26159495,0.18741131,0.113227665,0.20302892,0.29283017,0.38263142,0.47243267,0.5622339,0.4997635,0.43729305,0.37482262,0.31235218,0.24988174,0.20693332,0.16008049,0.113227665,0.07027924,0.023426414,0.20693332,0.39044023,0.57394713,0.75354964,0.93705654,0.8316377,0.7262188,0.62079996,0.5192855,0.41386664,0.3318742,0.24597734,0.1639849,0.08199245,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.78088045,1.3743496,1.9639144,2.5573835,3.1508527,3.018103,2.8853533,2.7526035,2.619854,2.4871042,2.494913,2.5027218,2.5105307,2.5183394,2.5261483,3.6037633,4.6813784,5.758993,6.8366084,7.914223,9.0386915,10.163159,11.287627,12.412095,13.536563,11.845957,10.159255,8.468649,6.7780423,5.087436,4.743849,4.396357,4.0527697,3.7091823,3.3616903,4.0996222,4.8375545,5.575486,6.3134184,7.0513506,6.1025805,5.153811,4.2089458,3.260176,2.3114061,3.154757,3.998108,4.841459,5.6809053,6.524256,6.309514,6.094772,5.8800297,5.6652875,5.4505453,8.164105,10.881569,13.595129,16.30869,19.026152,16.69913,14.3682,12.041177,9.714153,7.387129,8.406178,9.4291315,10.44818,11.46723,12.486279,10.198298,7.914223,5.6262436,3.338264,1.0502841,1.2962615,1.5461433,1.7921207,2.0380979,2.2879796,3.2250361,4.1620927,5.099149,6.036206,6.9732623,6.5359693,6.094772,5.6535745,5.2162814,4.775084,4.806319,4.83365,4.8648853,4.8961205,4.9234514,4.165997,3.4046388,2.6432803,1.8858263,1.1244678,0.92534333,0.7262188,0.5231899,0.3240654,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.20693332,0.339683,0.47243267,0.60518235,0.737932,0.80821127,0.8784905,0.94876975,1.0190489,1.0893283,1.5578566,2.0263848,2.4988174,2.9673457,3.435874,2.920493,2.4012074,1.8858263,1.3665408,0.8511597,0.679366,0.5114767,0.339683,0.1717937,0.0,0.0,0.0,0.0,0.0,0.0,0.05466163,0.10932326,0.1639849,0.21864653,0.27330816,0.48414588,0.6949836,0.9058213,1.116659,1.3235924,1.3509232,1.3743496,1.4016805,1.4251068,1.4485333,1.1986516,0.94486535,0.6910792,0.44119745,0.18741131,0.1639849,0.14055848,0.12103647,0.09761006,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.046852827,0.07027924,0.093705654,0.113227665,0.13665408,0.14836729,0.15617609,0.1678893,0.1756981,0.18741131,0.19522011,0.20302892,0.21083772,0.21864653,0.22645533,0.23426414,0.23816854,0.24597734,0.25378615,0.26159495,0.26940376,0.27721256,0.28502136,0.29283017,0.30063897,0.3357786,0.3709182,0.40605783,0.44119745,0.47633708,0.5231899,0.5700427,0.61689556,0.6637484,0.7106012,0.58566034,0.46071947,0.3357786,0.21083772,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.10541886,0.21083772,0.31625658,0.42167544,0.5231899,0.74964523,0.97610056,1.1986516,1.4251068,1.6515622,1.3743496,1.0932326,0.8160201,0.5388075,0.26159495,0.21083772,0.15617609,0.10541886,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14446288,0.21864653,0.28892577,0.3631094,0.37482262,0.38653582,0.39824903,0.41386664,0.42557985,0.46071947,0.4997635,0.5388075,0.57394713,0.61299115,0.5270943,0.44119745,0.359205,0.27330816,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.078088045,0.093705654,0.10932326,0.12103647,0.13665408,0.15227169,0.1678893,0.1835069,0.19912452,0.21083772,0.21864653,0.22645533,0.23426414,0.24207294,0.24988174,0.3513962,0.44900626,0.5505207,0.6481308,0.74964523,0.8667773,0.98000497,1.0932326,1.2103647,1.3235924,1.2220778,1.1205635,1.0190489,0.9136301,0.81211567,0.74574083,0.6832704,0.61689556,0.5544251,0.48805028,0.47633708,0.46852827,0.45681506,0.44900626,0.43729305,0.43338865,0.43338865,0.42948425,0.42557985,0.42557985,0.39434463,0.359205,0.3279698,0.29673457,0.26159495,0.21864653,0.1756981,0.13665408,0.093705654,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.05466163,0.10932326,0.1639849,0.21864653,0.27330816,0.24597734,0.21864653,0.19131571,0.1639849,0.13665408,0.5583295,0.97610056,1.397776,1.8194515,2.2372224,2.1044729,1.9717231,1.8389735,1.7062237,1.5734742,1.3626363,1.1517987,0.93705654,0.7262188,0.5114767,0.43729305,0.3631094,0.28892577,0.21083772,0.13665408,0.24597734,0.359205,0.46852827,0.57785153,0.6871748,0.58566034,0.48805028,0.38653582,0.28892577,0.18741131,0.15617609,0.12884527,0.09761006,0.06637484,0.039044023,0.15617609,0.27330816,0.39044023,0.5075723,0.62470436,0.5544251,0.48414588,0.41386664,0.3435874,0.27330816,0.21864653,0.1639849,0.10932326,0.05466163,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.5192855,0.9136301,1.3118792,1.7062237,2.1005683,2.05762,2.0146716,1.9717231,1.9287747,1.8858263,2.0927596,2.2957885,2.5027218,2.7057507,2.912684,3.7208953,4.533011,5.3412223,6.153338,6.9615493,7.8751793,8.78881,9.698535,10.612165,11.525795,10.366188,9.20658,8.043069,6.883461,5.7238536,5.571582,5.4154058,5.2592297,5.1030536,4.950782,5.4388323,5.9268827,6.4110284,6.899079,7.387129,6.524256,5.657479,4.7907014,3.9278288,3.0610514,3.4202564,3.775557,4.134762,4.493967,4.8492675,4.689187,4.5291066,4.369026,4.2089458,4.0488653,6.2587566,8.468649,10.67854,12.888432,15.098324,13.075843,11.053363,9.030883,7.008402,4.985922,7.4691215,9.948417,12.427712,14.907008,17.386303,14.188598,10.986988,7.7892823,4.5876727,1.3860629,1.6632754,1.9443923,2.2216048,2.4988174,2.77603,3.7247996,4.6735697,5.6262436,6.575013,7.523783,7.37932,7.230953,7.082586,6.9342184,6.785851,6.883461,6.9771667,7.0708723,7.168483,7.262188,6.1455293,5.0327744,3.9161155,2.803361,1.6867018,1.3860629,1.0893283,0.78868926,0.48805028,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.12103647,0.20693332,0.29283017,0.37872702,0.46071947,0.659844,0.8589685,1.0541886,1.2533131,1.4485333,1.999054,2.5456703,3.0922866,3.638903,4.1894236,3.435874,2.6823244,1.9287747,1.1791295,0.42557985,0.339683,0.25378615,0.1717937,0.08589685,0.0,0.0,0.0,0.0,0.0,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.42948425,0.7223144,1.0151446,1.3079748,1.6008049,1.6632754,1.7257458,1.7882162,1.8506867,1.9131571,1.5812829,1.2494087,0.9136301,0.58175594,0.24988174,0.21864653,0.19131571,0.16008049,0.12884527,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.031235218,0.046852827,0.06637484,0.08199245,0.10151446,0.10541886,0.10932326,0.113227665,0.12103647,0.12494087,0.12103647,0.12103647,0.11713207,0.113227665,0.113227665,0.12103647,0.13274968,0.14055848,0.15227169,0.1639849,0.16008049,0.15617609,0.15617609,0.15227169,0.14836729,0.21864653,0.28502136,0.3513962,0.42167544,0.48805028,0.5036679,0.5231899,0.5388075,0.5583295,0.57394713,0.47633708,0.37482262,0.27330816,0.1756981,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.14055848,0.28111696,0.42167544,0.5583295,0.698888,0.999527,1.3001659,1.6008049,1.901444,2.1981785,1.8311646,1.4602464,1.0893283,0.71841,0.3513962,0.28111696,0.21083772,0.14055848,0.07027924,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.042948425,0.08589685,0.12884527,0.1717937,0.21083772,0.26159495,0.31235218,0.3631094,0.41386664,0.46071947,0.4997635,0.5388075,0.57394713,0.61299115,0.6481308,0.5700427,0.49195468,0.40996224,0.3318742,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,0.07027924,0.078088045,0.08589685,0.093705654,0.10151446,0.10932326,0.113227665,0.12103647,0.12884527,0.13665408,0.14836729,0.15617609,0.1678893,0.1756981,0.18741131,0.24988174,0.31235218,0.37482262,0.43729305,0.4997635,0.6559396,0.8160201,0.97219616,1.1283722,1.2884527,1.2181735,1.1478943,1.077615,1.0073358,0.93705654,0.8667773,0.79649806,0.7262188,0.6559396,0.58566034,0.5192855,0.45291066,0.38653582,0.31625658,0.24988174,0.30454338,0.359205,0.41386664,0.46852827,0.5231899,0.47633708,0.42948425,0.38263142,0.3357786,0.28892577,0.23426414,0.1835069,0.12884527,0.078088045,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.12884527,0.12103647,0.113227665,0.10932326,0.10151446,0.3240654,0.5466163,0.76916724,0.9917182,1.2142692,1.2533131,1.2923572,1.3314011,1.3743496,1.4133936,1.2376955,1.0619974,0.8862993,0.7106012,0.5388075,0.46071947,0.38653582,0.31235218,0.23816854,0.1639849,0.29283017,0.42167544,0.5544251,0.6832704,0.81211567,0.6754616,0.5388075,0.39824903,0.26159495,0.12494087,0.10932326,0.093705654,0.078088045,0.06637484,0.05075723,0.10151446,0.15617609,0.20693332,0.26159495,0.31235218,0.27721256,0.24207294,0.20693332,0.1717937,0.13665408,0.10932326,0.08199245,0.05466163,0.027330816,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.26159495,0.45681506,0.6559396,0.8511597,1.0502841,1.097137,1.1439898,1.1908426,1.2415999,1.2884527,1.6906061,2.0927596,2.494913,2.8970666,3.2992198,3.8419318,4.3846436,4.927356,5.4700675,6.012779,6.7116675,7.4105554,8.113348,8.812236,9.511124,8.882515,8.253906,7.621393,6.9927845,6.364176,6.3993154,6.434455,6.46569,6.5008297,6.5359693,6.774138,7.012306,7.250475,7.4886436,7.726812,6.942027,6.1611466,5.376362,4.5954814,3.8106966,3.6857557,3.5569105,3.4280653,3.3031244,3.174279,3.06886,2.9634414,2.8580225,2.7565079,2.6510892,4.3534083,6.0596323,7.7658563,9.468176,11.174399,9.456462,7.7385254,6.0205884,4.3065557,2.5886188,6.5281606,10.467703,14.407245,18.346786,22.286327,18.174992,14.063657,9.948417,5.8370814,1.7257458,2.0341935,2.338737,2.6471848,2.9556324,3.2640803,4.224563,5.1889505,6.1494336,7.113821,8.074304,8.218767,8.36323,8.511597,8.65606,8.800523,8.960603,9.120684,9.280765,9.440845,9.600925,8.128965,6.66091,5.1889505,3.7208953,2.2489357,1.8506867,1.4485333,1.0502841,0.6481308,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.5114767,0.8355421,1.1635119,1.4875772,1.8116426,2.436347,3.0610514,3.6857557,4.3143644,4.939069,3.951255,2.9634414,1.9756275,0.9878138,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.37482262,0.74964523,1.1244678,1.4992905,1.8741131,1.9756275,2.0732377,2.174752,2.2762666,2.3738766,1.9639144,1.5500476,1.1361811,0.7262188,0.31235218,0.27330816,0.23816854,0.19912452,0.1639849,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.48805028,0.47633708,0.46071947,0.44900626,0.43729305,0.3631094,0.28892577,0.21083772,0.13665408,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.1756981,0.3513962,0.5231899,0.698888,0.8745861,1.2494087,1.6242313,1.999054,2.3738766,2.7486992,2.2879796,1.8233559,1.3626363,0.9019169,0.43729305,0.3513962,0.26159495,0.1756981,0.08589685,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.14836729,0.23816854,0.3240654,0.41386664,0.4997635,0.5388075,0.57394713,0.61299115,0.6481308,0.6871748,0.61299115,0.5388075,0.46071947,0.38653582,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.14836729,0.1756981,0.19912452,0.22645533,0.24988174,0.44900626,0.6481308,0.8511597,1.0502841,1.2494087,1.2142692,1.175225,1.1361811,1.1010414,1.0619974,0.9878138,0.9136301,0.8394465,0.76135844,0.6871748,0.5622339,0.43729305,0.31235218,0.18741131,0.062470436,0.1756981,0.28892577,0.39824903,0.5114767,0.62470436,0.5622339,0.4997635,0.43729305,0.37482262,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.39824903,0.61299115,0.8238289,1.038571,1.2494087,1.1127546,0.97610056,0.8394465,0.698888,0.5622339,0.48805028,0.41386664,0.3357786,0.26159495,0.18741131,0.3357786,0.48805028,0.63641757,0.78868926,0.93705654,0.76135844,0.58566034,0.41386664,0.23816854,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13665408,0.27330816,0.41386664,0.5505207,0.6871748,1.2884527,1.8858263,2.4871042,3.0883822,3.6857557,3.9629683,4.2362766,4.513489,4.786797,5.0640097,5.548156,6.036206,6.524256,7.012306,7.5003567,7.3988423,7.3012323,7.1997175,7.098203,7.000593,7.223144,7.4495993,7.676055,7.898606,8.125061,8.113348,8.101635,8.086017,8.074304,8.062591,7.363703,6.66091,5.9620223,5.263134,4.564246,3.951255,3.338264,2.7252727,2.1122816,1.4992905,1.4485333,1.4016805,1.3509232,1.3001659,1.2494087,2.4519646,3.6506162,4.8492675,6.0518236,7.250475,5.8370814,4.423688,3.0141985,1.6008049,0.18741131,5.5871997,10.986988,16.386776,21.786564,27.186354,22.161386,17.136421,12.111456,7.08649,2.0615244,2.4012074,2.736986,3.076669,3.4124475,3.7482262,4.7243266,5.700427,6.676528,7.648724,8.624825,9.062118,9.499411,9.936704,10.373997,10.81129,11.037745,11.2642,11.486752,11.713207,11.935758,10.112402,8.289046,6.461786,4.6384296,2.8111696,2.3114061,1.8116426,1.3118792,0.81211567,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3279698,0.6559396,0.98390937,1.3118792,1.6359446,1.3157835,0.9917182,0.6715572,0.3474918,0.023426414,0.023426414,0.019522011,0.015617609,0.015617609,0.011713207,0.031235218,0.05075723,0.07418364,0.093705654,0.113227665,0.13665408,0.1639849,0.18741131,0.21083772,0.23816854,0.19131571,0.14055848,0.093705654,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.93315214,1.815547,2.697942,3.5803368,4.462732,4.6657605,4.872694,5.0757227,5.282656,5.4856853,4.7633705,4.041056,3.3187418,2.5964274,1.8741131,1.7257458,1.5812829,1.4329157,1.2845483,1.1361811,1.2259823,1.3118792,1.4016805,1.4875772,1.5734742,1.9248703,2.2762666,2.6237583,2.9751544,3.3265507,3.5842414,3.8458362,4.1035266,4.365122,4.6267166,3.9434462,3.260176,2.5769055,1.893635,1.2142692,2.182561,3.1508527,4.123049,5.0913405,6.0635366,7.0357327,8.011833,8.987934,9.964035,10.936231,10.249056,9.561881,8.874706,8.187531,7.5003567,6.559396,5.6145306,4.6735697,3.7287042,2.787743,2.7526035,2.717464,2.6823244,2.6471848,2.612045,2.2645533,1.9170616,1.5695697,1.2220778,0.8745861,0.79649806,0.7145056,0.63641757,0.5544251,0.47633708,0.39044023,0.30454338,0.21864653,0.13665408,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.07027924,0.08980125,0.10932326,0.12884527,0.14836729,0.3318742,0.5114767,0.6910792,0.8706817,1.0502841,0.94486535,0.8394465,0.7340276,0.62860876,0.5231899,0.5427119,0.5583295,0.57785153,0.59346914,0.61299115,0.59737355,0.58175594,0.5661383,0.5544251,0.5388075,0.5700427,0.60127795,0.63641757,0.6676528,0.698888,0.999527,1.3001659,1.6008049,1.901444,2.1981785,1.8584955,1.5149081,1.1713207,0.8316377,0.48805028,0.39044023,0.29283017,0.19522011,0.09761006,0.0,0.07418364,0.14446288,0.21864653,0.28892577,0.3631094,0.46462387,0.5661383,0.6715572,0.77307165,0.8745861,0.79259366,0.7106012,0.62860876,0.5466163,0.46071947,0.5309987,0.60127795,0.6715572,0.7418364,0.81211567,0.7106012,0.61299115,0.5114767,0.41386664,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.12103647,0.19131571,0.26159495,0.3318742,0.39824903,0.43338865,0.46462387,0.4958591,0.5309987,0.5622339,0.4997635,0.43729305,0.37482262,0.31235218,0.24988174,0.21083772,0.1717937,0.12884527,0.08980125,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.058566034,0.07027924,0.078088045,0.08980125,0.10151446,0.12103647,0.14055848,0.16008049,0.1796025,0.19912452,0.359205,0.5192855,0.679366,0.8394465,0.999527,0.96829176,0.94096094,0.9097257,0.8784905,0.8511597,0.78868926,0.7301232,0.6715572,0.60908675,0.5505207,0.44900626,0.3513962,0.24988174,0.14836729,0.05075723,0.14055848,0.23035973,0.32016098,0.40996224,0.4997635,0.44900626,0.39824903,0.3513962,0.30063897,0.24988174,0.20302892,0.15617609,0.10932326,0.058566034,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.023426414,0.031235218,0.042948425,0.05075723,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.359205,0.5309987,0.7066968,0.8784905,1.0502841,0.95657855,0.8667773,0.77307165,0.679366,0.58566034,0.5466163,0.5075723,0.46852827,0.42557985,0.38653582,0.48024148,0.57394713,0.6637484,0.75745404,0.8511597,0.7066968,0.5661383,0.42167544,0.28111696,0.13665408,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10932326,0.21864653,0.3318742,0.44119745,0.5505207,1.0307622,1.5110037,1.9912452,2.4714866,2.951728,3.1781836,3.408543,3.638903,3.8692627,4.0996222,4.572055,5.044488,5.5169206,5.989353,6.461786,6.4500723,6.4383593,6.426646,6.4110284,6.3993154,6.5437784,6.6843367,6.8287997,6.969358,7.113821,7.2582836,7.406651,7.5550184,7.703386,7.8517528,7.2192397,6.590631,5.958118,5.3295093,4.7009,4.1464753,3.5881457,3.0337205,2.4792955,1.9248703,2.0810463,2.233318,2.3894942,2.5456703,2.7018464,3.5491016,4.4002614,5.251421,6.098676,6.949836,6.774138,6.5945354,6.4188375,6.239235,6.0635366,9.276859,12.486279,15.699601,18.912924,22.126247,18.124235,14.126127,10.124115,6.126007,2.1239948,2.5534792,2.9868677,3.416352,3.8458362,4.2753205,5.2358036,6.196286,7.1567693,8.113348,9.073831,9.265146,9.456462,9.643873,9.835189,10.0265045,10.541886,11.053363,11.568744,12.084125,12.599506,10.932326,9.265146,7.5979667,5.930787,4.263607,3.814601,3.3694992,2.920493,2.4714866,2.0263848,1.999054,1.9756275,1.9482968,1.9248703,1.901444,1.6632754,1.4251068,1.1869383,0.94876975,0.7106012,0.5700427,0.42557985,0.28502136,0.14446288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6559396,1.3118792,1.9639144,2.619854,3.2757936,2.631567,1.9834363,1.33921,0.6949836,0.05075723,0.046852827,0.039044023,0.03513962,0.031235218,0.023426414,0.039044023,0.05466163,0.07027924,0.08589685,0.10151446,0.1756981,0.24988174,0.3240654,0.39824903,0.47633708,0.37872702,0.28502136,0.19131571,0.093705654,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,1.8663043,3.631094,5.395884,7.1606736,8.925464,9.335425,9.745388,10.155351,10.565312,10.975275,9.530646,8.086017,6.6413884,5.196759,3.7482262,3.455396,3.1586614,2.8658314,2.5690966,2.2762666,2.4129205,2.5495746,2.6862288,2.8267872,2.9634414,3.338264,3.7130866,4.087909,4.462732,4.8375545,4.732136,4.6267166,4.521298,4.415879,4.3143644,3.9356375,3.5569105,3.1781836,2.803361,2.4246337,4.365122,6.3056097,8.246098,10.186585,12.123169,14.07537,16.023666,17.975868,19.924164,21.876366,20.502016,19.123762,17.749413,16.375063,15.000713,12.740065,10.479416,8.218767,5.958118,3.7013733,3.5295796,3.3616903,3.1898966,3.018103,2.8502135,2.5690966,2.2840753,2.0029583,1.7218413,1.43682,1.3157835,1.1908426,1.0698062,0.94876975,0.8238289,0.6676528,0.5114767,0.3513962,0.19522011,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.08980125,0.14055848,0.19522011,0.24597734,0.30063897,0.5583295,0.8199245,1.0815194,1.33921,1.6008049,1.4016805,1.2064602,1.0073358,0.80821127,0.61299115,0.7223144,0.8316377,0.94096094,1.0541886,1.1635119,1.1439898,1.1283722,1.1088502,1.0932326,1.0737107,0.96438736,0.8550641,0.74574083,0.63641757,0.5231899,0.74964523,0.97610056,1.1986516,1.4251068,1.6515622,1.4290112,1.2064602,0.98390937,0.76135844,0.5388075,0.42948425,0.3240654,0.21474212,0.10932326,0.0,0.14446288,0.28892577,0.43338865,0.58175594,0.7262188,0.8784905,1.0346665,1.1908426,1.3431144,1.4992905,1.3860629,1.2689307,1.1557031,1.038571,0.92534333,1.0659018,1.2064602,1.3431144,1.4836729,1.6242313,1.4251068,1.2259823,1.0268579,0.8238289,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.08980125,0.14055848,0.19522011,0.24597734,0.30063897,0.3279698,0.3553006,0.38263142,0.40996224,0.43729305,0.38653582,0.3357786,0.28892577,0.23816854,0.18741131,0.15617609,0.12884527,0.09761006,0.06637484,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.046852827,0.05075723,0.058566034,0.06637484,0.07418364,0.08980125,0.10541886,0.12103647,0.13665408,0.14836729,0.26940376,0.39044023,0.5114767,0.62860876,0.74964523,0.7262188,0.7066968,0.6832704,0.659844,0.63641757,0.59346914,0.5466163,0.5036679,0.45681506,0.41386664,0.3357786,0.26159495,0.18741131,0.113227665,0.039044023,0.10541886,0.1717937,0.23816854,0.30844778,0.37482262,0.3357786,0.30063897,0.26159495,0.22645533,0.18741131,0.15617609,0.12103647,0.08980125,0.058566034,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.031235218,0.039044023,0.046852827,0.05466163,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.32016098,0.45291066,0.58566034,0.71841,0.8511597,0.80430686,0.75354964,0.7066968,0.659844,0.61299115,0.60908675,0.60127795,0.59737355,0.59346914,0.58566034,0.62079996,0.6559396,0.6910792,0.7262188,0.76135844,0.6520352,0.5427119,0.43338865,0.3240654,0.21083772,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08199245,0.1639849,0.24597734,0.3318742,0.41386664,0.77307165,1.1322767,1.4914817,1.8506867,2.2137961,2.397303,2.5808098,2.7682211,2.951728,3.1391394,3.5959544,4.0527697,4.5095844,4.9663997,5.423215,5.5013027,5.575486,5.64967,5.7238536,5.801942,5.860508,5.919074,5.9815445,6.04011,6.098676,6.407124,6.715572,7.0240197,7.328563,7.6370106,7.0786815,6.5164475,5.958118,5.395884,4.8375545,4.3416953,3.8419318,3.3460727,2.8463092,2.35045,2.7096553,3.06886,3.4319696,3.7911747,4.1503797,4.650143,5.1499066,5.64967,6.1494336,6.649197,7.70729,8.765383,9.823476,10.881569,11.935758,12.962616,13.985569,15.012426,16.039284,17.062239,14.087084,11.111929,8.136774,5.1616197,2.1864653,2.7096553,3.232845,3.7560349,4.279225,4.7985106,5.743376,6.688241,7.633106,8.581876,9.526741,9.468176,9.40961,9.351044,9.296382,9.237816,10.042123,10.84643,11.650736,12.458947,13.263254,11.752251,10.241247,8.734148,7.223144,5.7121406,5.3177958,4.9234514,4.5291066,4.1308575,3.736513,3.7482262,3.7638438,3.775557,3.78727,3.7989833,3.3265507,2.8502135,2.3738766,1.901444,1.4251068,1.1400855,0.8550641,0.5700427,0.28502136,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.98390937,1.9639144,2.9478238,3.9317331,4.911738,3.9434462,2.979059,2.0107672,1.0424755,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.046852827,0.058566034,0.06637484,0.078088045,0.08589685,0.21083772,0.3357786,0.46071947,0.58566034,0.7106012,0.5700427,0.42557985,0.28502136,0.14055848,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,2.795552,5.446641,8.093826,10.741011,13.388195,14.001186,14.618082,15.231073,15.847969,16.46096,14.294017,12.127073,9.96013,7.793187,5.6262436,5.181142,4.7399445,4.298747,3.853645,3.4124475,3.5998588,3.78727,3.9746814,4.1620927,4.349504,4.7516575,5.1499066,5.548156,5.950309,6.348558,5.8800297,5.4115014,4.939069,4.4705405,3.998108,3.9278288,3.853645,3.7833657,3.7091823,3.638903,6.547683,9.456462,12.369146,15.277926,18.186707,21.111103,24.0355,26.963802,29.888199,32.812595,30.751072,28.685644,26.624119,24.562595,22.50107,18.920732,15.344301,11.767868,8.191436,4.6110992,4.3065557,4.0020123,3.697469,3.3929255,3.0883822,2.8697357,2.6510892,2.436347,2.2177005,1.999054,1.8350691,1.6710842,1.5031948,1.33921,1.175225,0.94486535,0.7145056,0.48414588,0.25378615,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.10932326,0.19522011,0.28111696,0.3631094,0.44900626,0.78868926,1.1283722,1.4719596,1.8116426,2.1513257,1.8584955,1.5695697,1.2806439,0.9917182,0.698888,0.9019169,1.1049459,1.3079748,1.5110037,1.7140326,1.6906061,1.6710842,1.6515622,1.6320401,1.6125181,1.358732,1.1088502,0.8550641,0.60127795,0.3513962,0.4997635,0.6481308,0.80040246,0.94876975,1.1010414,0.9956226,0.8941081,0.79259366,0.6910792,0.58566034,0.46852827,0.3513962,0.23426414,0.11713207,0.0,0.21864653,0.43338865,0.6520352,0.8706817,1.0893283,1.2962615,1.5031948,1.7101282,1.9170616,2.1239948,1.9756275,1.8311646,1.6827974,1.53443,1.3860629,1.5969005,1.8077383,2.018576,2.2294137,2.436347,2.135708,1.8389735,1.5383345,1.2376955,0.93705654,0.74964523,0.5622339,0.37482262,0.18741131,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.058566034,0.093705654,0.12884527,0.1639849,0.19912452,0.22255093,0.24597734,0.26940376,0.28892577,0.31235218,0.27330816,0.23816854,0.19912452,0.1639849,0.12494087,0.10541886,0.08589685,0.06637484,0.046852827,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.031235218,0.03513962,0.039044023,0.046852827,0.05075723,0.058566034,0.07027924,0.078088045,0.08980125,0.10151446,0.1796025,0.26159495,0.339683,0.42167544,0.4997635,0.48414588,0.46852827,0.45681506,0.44119745,0.42557985,0.39434463,0.3631094,0.3357786,0.30454338,0.27330816,0.22645533,0.1756981,0.12494087,0.07418364,0.023426414,0.07027924,0.113227665,0.16008049,0.20693332,0.24988174,0.22645533,0.19912452,0.1756981,0.14836729,0.12494087,0.10932326,0.08980125,0.07418364,0.05466163,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.042948425,0.046852827,0.05075723,0.058566034,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.28111696,0.3709182,0.46462387,0.5583295,0.6481308,0.6481308,0.6442264,0.6442264,0.64032197,0.63641757,0.6676528,0.698888,0.7262188,0.75745404,0.78868926,0.76526284,0.7418364,0.71841,0.698888,0.6754616,0.59737355,0.5192855,0.44119745,0.3631094,0.28892577,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05466163,0.10932326,0.1639849,0.21864653,0.27330816,0.5153811,0.75354964,0.9956226,1.2337911,1.475864,1.6164225,1.7530766,1.893635,2.0341935,2.174752,2.6159496,3.0610514,3.5022488,3.9434462,4.388548,4.548629,4.7126136,4.8765984,5.036679,5.2006636,5.1772375,5.153811,5.134289,5.1108627,5.087436,5.5559645,6.0205884,6.4891167,6.957645,7.426173,6.9342184,6.446168,5.9542136,5.466163,4.9742084,4.5369153,4.095718,3.6545205,3.213323,2.77603,3.338264,3.9044023,4.4705405,5.036679,5.5989127,5.7511845,5.899552,6.0518236,6.2001905,6.348558,8.644346,10.936231,13.228115,15.519999,17.811884,16.64837,15.488764,14.325252,13.16174,11.998228,10.049932,8.101635,6.1494336,4.2011366,2.2489357,2.8658314,3.4788225,4.095718,4.7087092,5.3256044,6.2548523,7.1841,8.113348,9.0465,9.975748,9.671205,9.366661,9.058213,8.75367,8.449126,9.546264,10.639496,11.736633,12.829865,13.923099,12.572175,11.221252,9.866425,8.515501,7.1606736,6.8209906,6.477403,6.133816,5.794133,5.4505453,5.5013027,5.548156,5.5989127,5.64967,5.700427,4.985922,4.2753205,3.5608149,2.8502135,2.135708,1.7101282,1.2806439,0.8550641,0.42557985,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.3118792,2.619854,3.9317331,5.239708,6.551587,5.2592297,3.970777,2.67842,1.3899672,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.05466163,0.058566034,0.06637484,0.07027924,0.07418364,0.24988174,0.42557985,0.60127795,0.77307165,0.94876975,0.76135844,0.5700427,0.37872702,0.19131571,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,3.7287042,7.2582836,10.791768,14.321347,17.850927,18.67085,19.490776,20.310701,21.130625,21.95055,19.061293,16.172033,13.2788725,10.389614,7.5003567,6.910792,6.321227,5.7316628,5.138193,4.548629,4.786797,5.024966,5.263134,5.5013027,5.7394714,6.1611466,6.5867267,7.012306,7.437886,7.8634663,7.027924,6.192382,5.35684,4.521298,3.6857557,3.9200199,4.154284,4.3846436,4.618908,4.8492675,8.730244,12.611219,16.48829,20.369267,24.250242,28.15074,32.05124,35.951736,39.848328,43.74883,41.00013,38.25143,35.498825,32.750126,30.001427,25.105307,20.209187,15.313066,10.42085,5.5247293,5.083532,4.646239,4.2050414,3.7638438,3.3265507,3.174279,3.018103,2.8658314,2.7135596,2.5612879,2.3543546,2.1474214,1.9404879,1.7335546,1.5266213,1.2220778,0.92143893,0.61689556,0.31625658,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.12884527,0.24597734,0.3631094,0.48414588,0.60127795,1.0190489,1.4407244,1.8584955,2.280171,2.7018464,2.3192148,1.9365835,1.5539521,1.1713207,0.78868926,1.0815194,1.3782539,1.6710842,1.9678187,2.260649,2.241127,2.2177005,2.194274,2.1708477,2.1513257,1.7530766,1.358732,0.96438736,0.5700427,0.1756981,0.24988174,0.3240654,0.39824903,0.47633708,0.5505207,0.5661383,0.58566034,0.60127795,0.62079996,0.63641757,0.5114767,0.38263142,0.25378615,0.12884527,0.0,0.28892577,0.58175594,0.8706817,1.1596074,1.4485333,1.7101282,1.9717231,2.2294137,2.4910088,2.7486992,2.5690966,2.3894942,2.2098918,2.0302892,1.8506867,2.1318035,2.4090161,2.690133,2.97125,3.2484627,2.8502135,2.4519646,2.0498111,1.6515622,1.2494087,0.999527,0.74964523,0.4997635,0.24988174,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.031235218,0.046852827,0.06637484,0.08199245,0.10151446,0.11713207,0.13665408,0.15227169,0.1717937,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.05075723,0.042948425,0.031235218,0.023426414,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.015617609,0.015617609,0.019522011,0.023426414,0.023426414,0.031235218,0.03513962,0.039044023,0.046852827,0.05075723,0.08980125,0.12884527,0.1717937,0.21083772,0.24988174,0.24207294,0.23426414,0.22645533,0.21864653,0.21083772,0.19912452,0.1835069,0.1678893,0.15227169,0.13665408,0.113227665,0.08589685,0.062470436,0.039044023,0.011713207,0.03513962,0.058566034,0.078088045,0.10151446,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.058566034,0.058566034,0.05466163,0.05075723,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05466163,0.058566034,0.058566034,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.23816854,0.29283017,0.3435874,0.39824903,0.44900626,0.49195468,0.5349031,0.57785153,0.62079996,0.6637484,0.7262188,0.79259366,0.8589685,0.92143893,0.9878138,0.9058213,0.8277333,0.74574083,0.6676528,0.58566034,0.5427119,0.4958591,0.45291066,0.40605783,0.3631094,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.25769055,0.37872702,0.4958591,0.61689556,0.737932,0.8316377,0.92924774,1.0229534,1.116659,1.2142692,1.639849,2.069333,2.494913,2.9243972,3.349977,3.5998588,3.8497405,4.0996222,4.349504,4.5993857,4.493967,4.388548,4.283129,4.181615,4.0761957,4.7009,5.3295093,5.958118,6.5867267,7.211431,6.79366,6.3719845,5.9542136,5.532538,5.1108627,4.728231,4.3455997,3.9668727,3.5842414,3.2016098,3.970777,4.7399445,5.5091114,6.278279,7.0513506,6.8483214,6.649197,6.4500723,6.250948,6.0518236,9.577498,13.103174,16.632753,20.158428,23.68801,20.338032,16.988054,13.638077,10.2881,6.9381227,6.012779,5.087436,4.1620927,3.2367494,2.3114061,3.018103,3.7287042,4.435401,5.142098,5.8487945,6.7663293,7.6799593,8.59359,9.511124,10.424754,9.874233,9.319808,8.769287,8.214863,7.6643414,9.0465,10.432563,11.818625,13.200784,14.586847,13.392099,12.197352,11.002605,9.807858,8.6131115,8.324185,8.031356,7.7424297,7.453504,7.1606736,7.250475,7.336372,7.426173,7.5120697,7.601871,6.649197,5.700427,4.7516575,3.7989833,2.8502135,2.280171,1.7101282,1.1400855,0.5700427,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.6359446,3.2757936,4.911738,6.551587,8.187531,6.575013,4.9624953,3.349977,1.737459,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.28892577,0.5114767,0.737932,0.96438736,1.1869383,0.94876975,0.7106012,0.47633708,0.23816854,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,4.661856,9.073831,13.4858055,17.901684,22.31366,23.336613,24.36347,25.386423,26.41328,27.436235,23.824663,20.21309,16.601519,12.986042,9.37447,8.636538,7.898606,7.1606736,6.426646,5.688714,5.9737353,6.262661,6.551587,6.8366084,7.125534,7.57454,8.023546,8.476458,8.925464,9.37447,8.175818,6.9732623,5.774611,4.575959,3.3734035,3.912211,4.4510183,4.985922,5.5247293,6.0635366,10.912805,15.762072,20.61134,25.464512,30.31378,35.186474,40.063072,44.935764,49.812363,54.68896,51.249184,47.81331,44.37353,40.937656,37.501785,31.285975,25.074072,18.862167,12.650263,6.4383593,5.8644123,5.2865605,4.7126136,4.138666,3.5608149,3.474918,3.3890212,3.2992198,3.213323,3.1235218,2.87364,2.6237583,2.3738766,2.1239948,1.8741131,1.4992905,1.1244678,0.74964523,0.37482262,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14836729,0.30063897,0.44900626,0.60127795,0.74964523,1.2494087,1.7491722,2.2489357,2.7486992,3.2484627,2.77603,2.2996929,1.8233559,1.3509232,0.8745861,1.261122,1.6515622,2.0380979,2.4246337,2.8111696,2.787743,2.7643168,2.736986,2.7135596,2.6862288,2.1513257,1.6125181,1.0737107,0.5388075,0.0,0.0,0.0,0.0,0.0,0.0,0.13665408,0.27330816,0.41386664,0.5505207,0.6871748,0.5505207,0.41386664,0.27330816,0.13665408,0.0,0.3631094,0.7262188,1.0893283,1.4485333,1.8116426,2.1239948,2.436347,2.7486992,3.0610514,3.3734035,3.1625657,2.951728,2.736986,2.5261483,2.3114061,2.6628022,3.0141985,3.3616903,3.7130866,4.0605783,3.5608149,3.0610514,2.5612879,2.0615244,1.5617609,1.2494087,0.93705654,0.62470436,0.31235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,0.3357786,0.42557985,0.5114767,0.60127795,0.6871748,0.78868926,0.8862993,0.9878138,1.0893283,1.1869383,1.0502841,0.9136301,0.77307165,0.63641757,0.4997635,0.48805028,0.47633708,0.46071947,0.44900626,0.43729305,0.37482262,0.31235218,0.24988174,0.18741131,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.6637484,1.0737107,1.4875772,1.901444,2.3114061,2.6510892,2.9868677,3.3265507,3.6623292,3.998108,3.8106966,3.6232853,3.435874,3.2484627,3.0610514,3.8497405,4.6384296,5.423215,6.211904,7.000593,6.649197,6.3017054,5.950309,5.5989127,5.251421,4.9234514,4.5993857,4.2753205,3.951255,3.6232853,4.5993857,5.575486,6.551587,7.523783,8.499884,7.9493628,7.3988423,6.8483214,6.3017054,5.7511845,10.514555,15.274021,20.037392,24.800762,29.564135,24.023787,18.487345,12.950902,7.4144597,1.8741131,1.9756275,2.0732377,2.174752,2.2762666,2.3738766,3.174279,3.9746814,4.775084,5.575486,6.375889,7.2739015,8.175818,9.073831,9.975748,10.87376,10.073358,9.276859,8.476458,7.676055,6.8756523,8.550641,10.22563,11.900618,13.575606,15.250595,14.212025,13.173453,12.138786,11.100216,10.061645,9.823476,9.589212,9.351044,9.112875,8.874706,8.999647,9.124588,9.249529,9.37447,9.499411,8.312472,7.125534,5.938596,4.7516575,3.5608149,2.8502135,2.135708,1.4251068,0.7106012,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.3118792,2.619854,3.9317331,5.239708,6.551587,5.2592297,3.970777,2.67842,1.3899672,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.20693332,0.3631094,0.5231899,0.679366,0.8394465,0.98000497,1.1205635,1.2650263,1.4055848,1.5500476,1.5929961,1.6359446,1.678893,1.7218413,1.7608855,2.0927596,2.4207294,2.7526035,3.084478,3.4124475,3.474918,3.5373883,3.5998588,3.6623292,3.7247996,6.590631,9.460366,12.326198,15.195933,18.061766,18.838741,19.615717,20.396597,21.173573,21.95055,19.061293,16.168129,13.2788725,10.389614,7.5003567,6.910792,6.321227,5.7316628,5.138193,4.548629,4.7789884,5.009348,5.239708,5.4700675,5.700427,6.0596323,6.4188375,6.7780423,7.141152,7.5003567,6.7116675,5.919074,5.1303844,4.3416953,3.5491016,4.095718,4.646239,5.192855,5.7394714,6.2860875,10.03041,13.770826,17.515148,21.255566,24.999887,29.130745,33.265507,37.396366,41.531128,45.661983,42.975754,40.28562,37.599392,34.913166,32.22303,27.401094,22.575254,17.749413,12.923572,8.101635,8.031356,7.9610763,7.890797,7.8205175,7.7502384,8.101635,8.456935,8.8083315,9.159728,9.511124,9.347139,9.183154,9.019169,8.85128,8.687295,8.484266,8.281238,8.082112,7.8790836,7.676055,7.57454,7.47693,7.375416,7.2739015,7.1762915,6.9068875,6.6413884,6.3719845,6.1064854,5.8370814,5.3021784,4.7672753,4.2323723,3.697469,3.1625657,2.8658314,2.5690966,2.2684577,1.9717231,1.6749885,1.3782539,1.0815194,0.78088045,0.48414588,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.058566034,0.058566034,0.05466163,0.05075723,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.09761006,0.093705654,0.093705654,0.08980125,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.12103647,0.23816854,0.359205,0.48024148,0.60127795,1.0112402,1.4212024,1.8311646,2.241127,2.6510892,2.3075018,1.9639144,1.6242313,1.2806439,0.93705654,1.2064602,1.475864,1.7491722,2.018576,2.2879796,2.3231194,2.3621633,2.4012074,2.436347,2.475391,2.1669433,1.8584955,1.5539521,1.2455044,0.93705654,0.9097257,0.8823949,0.8550641,0.8277333,0.80040246,0.9019169,1.0034313,1.1088502,1.2103647,1.3118792,1.1713207,1.0268579,0.8862993,0.7418364,0.60127795,0.94486535,1.2884527,1.6359446,1.979532,2.3231194,2.5573835,2.7916477,3.0220075,3.2562714,3.4866312,3.3187418,3.1508527,2.9868677,2.8189783,2.6510892,2.8385005,3.0259118,3.213323,3.4007344,3.5881457,3.2875066,2.9868677,2.6862288,2.3855898,2.0888553,1.737459,1.3860629,1.038571,0.6871748,0.3357786,0.40996224,0.48414588,0.5544251,0.62860876,0.698888,0.74574083,0.78868926,0.8355421,0.8784905,0.92534333,1.0307622,1.1361811,1.2415999,1.3431144,1.4485333,1.261122,1.0737107,0.8862993,0.698888,0.5114767,0.40996224,0.30844778,0.20693332,0.10151446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05466163,0.058566034,0.058566034,0.062470436,0.08589685,0.10932326,0.12884527,0.15227169,0.1756981,0.1835069,0.19131571,0.19912452,0.20693332,0.21083772,0.30063897,0.39434463,0.48414588,0.57394713,0.6637484,0.7262188,0.79259366,0.8589685,0.92143893,0.9878138,0.8706817,0.75745404,0.6442264,0.5270943,0.41386664,0.40605783,0.39824903,0.39044023,0.38263142,0.37482262,0.32016098,0.26549935,0.21083772,0.15617609,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.5309987,0.8589685,1.1908426,1.5188124,1.8506867,2.1278992,2.4051118,2.6823244,2.959537,3.2367494,3.1000953,2.9634414,2.8267872,2.6862288,2.5495746,3.2445583,3.9395418,4.6345253,5.3295093,6.0244927,5.8292727,5.6340523,5.4388323,5.2436123,5.0483923,4.7907014,4.5369153,4.279225,4.0215344,3.7638438,4.4861584,5.2084727,5.930787,6.6531014,7.375416,7.0630636,6.754616,6.446168,6.133816,5.825368,9.866425,13.911386,17.952442,21.993498,26.038458,21.626484,17.218414,12.806439,8.398369,3.9863946,3.853645,3.7208953,3.5881457,3.4593005,3.3265507,3.6857557,4.0488653,4.4119744,4.775084,5.138193,6.0205884,6.9068875,7.793187,8.675582,9.561881,8.843472,8.128965,7.4105554,6.6921453,5.9737353,7.7111945,9.448653,11.186112,12.923572,14.661031,14.286208,13.907481,13.528754,13.153932,12.775204,12.431617,12.091934,11.748346,11.404759,11.061172,11.272009,11.482847,11.693685,11.900618,12.111456,10.741011,9.370565,8.0040245,6.6335793,5.263134,4.3534083,3.4436827,2.533957,1.6242313,0.7106012,0.5700427,0.42557985,0.28502136,0.14446288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.98390937,1.9639144,2.9478238,3.9317331,4.911738,3.9434462,2.979059,2.0107672,1.0424755,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.3513962,0.6676528,0.98390937,1.2962615,1.6125181,1.6710842,1.7335546,1.7921207,1.8506867,1.9131571,2.233318,2.5573835,2.8814487,3.2016098,3.5256753,4.185519,4.845363,5.505207,6.165051,6.824895,6.899079,6.9732623,7.0513506,7.125534,7.1997175,8.52331,9.846903,11.166591,12.490183,13.813775,14.34087,14.871868,15.402867,15.933866,16.46096,14.294017,12.127073,9.96013,7.793187,5.6262436,5.181142,4.7399445,4.298747,3.853645,3.4124475,3.5842414,3.7560349,3.9317331,4.1035266,4.2753205,4.5447245,4.814128,5.083532,5.35684,5.6262436,5.2436123,4.8648853,4.4861584,4.1035266,3.7247996,4.283129,4.841459,5.395884,5.9542136,6.5125427,9.148014,11.783486,14.418958,17.054428,19.685997,23.078922,26.467943,29.856964,33.245987,36.638912,34.69842,32.76184,30.825256,28.888672,26.948185,23.51231,20.076437,16.636658,13.200784,9.761005,10.198298,10.631687,11.06898,11.502369,11.935758,12.728352,13.520945,14.313539,15.1061325,15.8987255,15.820638,15.738646,15.660558,15.578565,15.500477,15.469242,15.441911,15.410676,15.37944,15.348206,15.14908,14.949956,14.750832,14.551707,14.348679,13.813775,13.2788725,12.743969,12.209065,11.674163,10.604357,9.534551,8.464745,7.394938,6.3251314,5.7316628,5.134289,4.5408196,3.9434462,3.349977,2.7565079,2.1591344,1.5656652,0.96829176,0.37482262,0.3240654,0.27330816,0.22645533,0.1756981,0.12494087,0.12103647,0.113227665,0.10932326,0.10541886,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.093705654,0.113227665,0.13665408,0.15617609,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.08980125,0.1796025,0.26940376,0.359205,0.44900626,0.76916724,1.0893283,1.4094892,1.7296503,2.0498111,1.8389735,1.6281357,1.4212024,1.2103647,0.999527,1.1517987,1.3040704,1.456342,1.6086137,1.7608855,1.8623998,1.9639144,2.0615244,2.1630387,2.260649,2.1864653,2.1083772,2.0302892,1.9522011,1.8741131,1.8194515,1.7647898,1.7101282,1.6554666,1.6008049,1.6671798,1.7335546,1.8038338,1.8702087,1.9365835,1.7882162,1.6437533,1.4953861,1.3470187,1.1986516,1.5266213,1.8545911,2.182561,2.5105307,2.8385005,2.9907722,3.1430438,3.2953155,3.4475873,3.5998588,3.4788225,3.3538816,3.232845,3.1118085,2.9868677,3.0141985,3.0376248,3.0610514,3.0883822,3.1118085,3.0141985,2.912684,2.8111696,2.7135596,2.612045,2.2255092,1.8389735,1.4485333,1.0619974,0.6754616,0.8199245,0.96438736,1.1088502,1.2533131,1.4016805,1.4914817,1.5812829,1.6710842,1.7608855,1.8506867,2.0459068,2.2450314,2.4441557,2.639376,2.8385005,2.475391,2.1122816,1.7491722,1.3860629,1.0268579,0.8199245,0.61689556,0.40996224,0.20693332,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.042948425,0.046852827,0.05075723,0.058566034,0.062470436,0.08199245,0.10151446,0.12103647,0.14055848,0.1639849,0.1639849,0.1678893,0.1717937,0.1717937,0.1756981,0.26940376,0.359205,0.45291066,0.5466163,0.63641757,0.6676528,0.698888,0.7262188,0.75745404,0.78868926,0.6949836,0.60127795,0.5114767,0.41777104,0.3240654,0.3240654,0.32016098,0.31625658,0.31625658,0.31235218,0.26549935,0.21864653,0.1717937,0.12103647,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.39824903,0.6442264,0.8941081,1.1400855,1.3860629,1.6047094,1.8233559,2.0380979,2.2567444,2.475391,2.3855898,2.2996929,2.2137961,2.1239948,2.0380979,2.639376,3.240654,3.8458362,4.447114,5.0483923,5.009348,4.970304,4.93126,4.8883114,4.8492675,4.661856,4.4705405,4.279225,4.0918136,3.900498,4.369026,4.841459,5.309987,5.7785153,6.250948,6.180669,6.1103897,6.04011,5.969831,5.899552,9.2221985,12.544845,15.867491,19.190138,22.512783,19.229181,15.949483,12.665881,9.382278,6.098676,5.735567,5.368553,5.0054436,4.6384296,4.2753205,4.2011366,4.126953,4.0488653,3.9746814,3.900498,4.7711797,5.6418614,6.5086384,7.37932,8.250002,7.6135845,6.9810715,6.3446536,5.708236,5.0757227,6.8756523,8.675582,10.475512,12.27544,14.07537,14.356487,14.641508,14.922626,15.203742,15.488764,15.039758,14.590752,14.145649,13.696643,13.251541,13.544372,13.841106,14.133936,14.430671,14.723501,13.173453,11.619501,10.065549,8.515501,6.9615493,5.8566036,4.747753,3.638903,2.533957,1.4251068,1.1400855,0.8550641,0.5700427,0.28502136,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6559396,1.3118792,1.9639144,2.619854,3.2757936,2.631567,1.9834363,1.33921,0.6949836,0.05075723,0.046852827,0.039044023,0.03513962,0.031235218,0.023426414,0.4958591,0.96829176,1.4407244,1.9131571,2.3855898,2.366068,2.3426414,2.3192148,2.2957885,2.2762666,2.8775444,3.4788225,4.084005,4.6852827,5.2865605,6.278279,7.266093,8.257811,9.245625,10.237343,10.323239,10.413041,10.498938,10.588739,10.674636,10.452085,10.229534,10.006983,9.784432,9.561881,9.846903,10.128019,10.409137,10.694158,10.975275,9.530646,8.086017,6.6413884,5.196759,3.7482262,3.455396,3.1586614,2.8658314,2.5690966,2.2762666,2.3894942,2.5066261,2.619854,2.7330816,2.8502135,3.0298162,3.2094188,3.3890212,3.5686235,3.7482262,3.7794614,3.8106966,3.8419318,3.8692627,3.900498,4.466636,5.036679,5.602817,6.168956,6.7389984,8.265619,9.792241,11.318862,12.849388,14.376009,17.023193,19.670378,22.317564,24.964748,27.611933,26.424995,25.238056,24.051117,22.86418,21.673336,19.623526,17.573715,15.523903,13.4740925,11.424281,12.365242,13.306203,14.243259,15.18422,16.125181,17.358973,18.58886,19.82265,21.056442,22.286327,22.294136,22.29804,22.301945,22.305851,22.31366,22.454218,22.59868,22.739239,22.883701,23.02426,22.723621,22.426888,22.126247,21.82561,21.52497,20.720663,19.92026,19.115953,18.315552,17.511244,15.906535,14.301826,12.697116,11.092407,9.487698,8.59359,7.703386,6.8092775,5.919074,5.024966,4.1308575,3.240654,2.3465457,1.456342,0.5622339,0.48805028,0.41386664,0.3357786,0.26159495,0.18741131,0.1796025,0.1717937,0.1639849,0.15617609,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.093705654,0.13665408,0.1756981,0.21864653,0.26159495,0.21083772,0.15617609,0.10541886,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.5309987,0.76135844,0.9917182,1.2181735,1.4485333,1.3743496,1.2962615,1.2181735,1.1400855,1.0619974,1.097137,1.1322767,1.1674163,1.2025559,1.2376955,1.4016805,1.5617609,1.7257458,1.8858263,2.0498111,2.2020829,2.3543546,2.5066261,2.6588979,2.8111696,2.7291772,2.6471848,2.5651922,2.4831998,2.4012074,2.4324427,2.463678,2.4988174,2.5300527,2.5612879,2.4090161,2.2567444,2.1044729,1.9522011,1.7999294,2.1083772,2.4207294,2.7291772,3.0415294,3.349977,3.4241607,3.49444,3.5686235,3.638903,3.7130866,3.6349986,3.5569105,3.4788225,3.4007344,3.3265507,3.1859922,3.049338,2.912684,2.77603,2.639376,2.736986,2.8385005,2.9361105,3.0376248,3.1391394,2.7135596,2.2879796,1.8623998,1.43682,1.0112402,1.2298868,1.4485333,1.6632754,1.8819219,2.1005683,2.233318,2.3699722,2.5066261,2.639376,2.77603,3.0649557,3.3538816,3.6467118,3.9356375,4.224563,3.6857557,3.1508527,2.612045,2.0732377,1.5383345,1.2298868,0.92143893,0.61689556,0.30844778,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.031235218,0.039044023,0.046852827,0.05466163,0.062470436,0.078088045,0.09761006,0.113227665,0.13274968,0.14836729,0.14836729,0.14446288,0.14055848,0.14055848,0.13665408,0.23426414,0.3279698,0.42167544,0.5192855,0.61299115,0.60908675,0.60127795,0.59737355,0.59346914,0.58566034,0.5192855,0.44900626,0.37872702,0.30844778,0.23816854,0.23816854,0.24207294,0.24597734,0.24597734,0.24988174,0.21083772,0.1717937,0.12884527,0.08980125,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.26549935,0.42948425,0.59346914,0.76135844,0.92534333,1.0815194,1.2415999,1.397776,1.5539521,1.7140326,1.6749885,1.6359446,1.6008049,1.5617609,1.5266213,2.0341935,2.5456703,3.0532427,3.5647192,4.0761957,4.1894236,4.3065557,4.4197836,4.5369153,4.650143,4.5291066,4.4041657,4.283129,4.1581883,4.037152,4.2557983,4.474445,4.689187,4.9078336,5.12648,5.2943697,5.466163,5.6340523,5.805846,5.9737353,8.577971,11.178304,13.78254,16.386776,18.987108,16.831879,14.676648,12.521418,10.366188,8.210958,7.6135845,7.016211,6.4188375,5.8214636,5.22409,4.7126136,4.2011366,3.6857557,3.174279,2.6628022,3.5178664,4.3729305,5.2279944,6.083059,6.9381227,6.3836975,5.833177,5.278752,4.728231,4.173806,6.036206,7.898606,9.761005,11.623405,13.4858055,14.430671,15.371632,16.316498,17.257458,18.19842,17.647898,17.093473,16.542952,15.988527,15.438006,15.816733,16.199366,16.578093,16.95682,17.335546,15.601992,13.868437,12.130978,10.397423,8.663869,7.355894,6.0518236,4.747753,3.4436827,2.135708,1.7101282,1.2806439,0.8550641,0.42557985,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3279698,0.6559396,0.98390937,1.3118792,1.6359446,1.3157835,0.9917182,0.6715572,0.3474918,0.023426414,0.023426414,0.019522011,0.015617609,0.015617609,0.011713207,0.6442264,1.2728351,1.901444,2.533957,3.1625657,3.057147,2.951728,2.8463092,2.7408905,2.639376,3.521771,4.4041657,5.2865605,6.168956,7.0513506,8.371038,9.690726,11.010414,12.330102,13.64979,13.751305,13.848915,13.950429,14.051944,14.149553,12.380859,10.61607,8.847376,7.0786815,5.3138914,5.349031,5.3841705,5.4193106,5.4505453,5.4856853,4.7633705,4.041056,3.3187418,2.5964274,1.8741131,1.7257458,1.5812829,1.4329157,1.2845483,1.1361811,1.1947471,1.2533131,1.3118792,1.3665408,1.4251068,1.5149081,1.6047094,1.6945106,1.7843118,1.8741131,2.3153105,2.7565079,3.193801,3.6349986,4.0761957,4.6540475,5.2318993,5.805846,6.3836975,6.9615493,7.3832245,7.800996,8.2226715,8.644346,9.062118,10.967466,12.872814,14.778163,16.683512,18.58886,18.151566,17.714273,17.273075,16.835783,16.398489,15.738646,15.074897,14.411149,13.751305,13.087557,14.532186,15.976814,17.421442,18.866072,20.310701,21.98569,23.656773,25.331762,27.002846,28.673931,28.763731,28.853533,28.943335,29.037039,29.12684,29.439194,29.75545,30.071707,30.384058,30.700315,30.302067,29.899912,29.501663,29.09951,28.701262,27.631454,26.56165,25.491842,24.41813,23.348326,21.208714,19.069101,16.92949,14.789876,12.650263,11.45942,10.268578,9.081639,7.890797,6.699954,5.5091114,4.318269,3.1313305,1.9404879,0.74964523,0.6481308,0.5505207,0.44900626,0.3513962,0.24988174,0.23816854,0.23035973,0.21864653,0.21083772,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.08980125,0.15617609,0.21864653,0.28502136,0.3513962,0.28111696,0.21083772,0.14055848,0.07027924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.28892577,0.42948425,0.5700427,0.7106012,0.8511597,0.9058213,0.96048295,1.0151446,1.0698062,1.1244678,1.0424755,0.96048295,0.8784905,0.79649806,0.7106012,0.93705654,1.1635119,1.3860629,1.6125181,1.8389735,2.2216048,2.6042364,2.9868677,3.3655949,3.7482262,3.638903,3.5295796,3.4202564,3.310933,3.2016098,3.1977055,3.193801,3.193801,3.1898966,3.1859922,3.0298162,2.87364,2.7135596,2.5573835,2.4012074,2.6940374,2.9868677,3.2757936,3.5686235,3.8614538,3.853645,3.8458362,3.8419318,3.8341231,3.8263142,3.7911747,3.7599394,3.7287042,3.6935644,3.6623292,3.3616903,3.0610514,2.7643168,2.463678,2.1630387,2.463678,2.7643168,3.0610514,3.3616903,3.6623292,3.2016098,2.736986,2.2762666,1.8116426,1.3509232,1.639849,1.9287747,2.2216048,2.5105307,2.7994564,2.979059,3.1586614,3.338264,3.521771,3.7013733,4.084005,4.466636,4.8492675,5.2318993,5.610626,4.900025,4.1894236,3.474918,2.7643168,2.0498111,1.639849,1.2298868,0.8199245,0.40996224,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.023426414,0.031235218,0.042948425,0.05075723,0.062470436,0.078088045,0.093705654,0.10932326,0.12103647,0.13665408,0.12884527,0.12103647,0.113227665,0.10932326,0.10151446,0.19912452,0.29673457,0.39434463,0.48805028,0.58566034,0.5466163,0.5075723,0.46852827,0.42557985,0.38653582,0.339683,0.29283017,0.24597734,0.19912452,0.14836729,0.15617609,0.1639849,0.1717937,0.1796025,0.18741131,0.15617609,0.12103647,0.08980125,0.058566034,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.13274968,0.21474212,0.29673457,0.37872702,0.46071947,0.5583295,0.6559396,0.75354964,0.8511597,0.94876975,0.96438736,0.97610056,0.9878138,0.999527,1.0112402,1.4290112,1.8467822,2.2645533,2.6823244,3.1000953,3.3694992,3.638903,3.9083066,4.181615,4.4510183,4.396357,4.3416953,4.283129,4.2284675,4.173806,4.138666,4.1035266,4.068387,4.0332475,3.998108,4.40807,4.8180323,5.2318993,5.6418614,6.0518236,7.9337454,9.815667,11.697589,13.579511,15.461433,14.434575,13.407718,12.380859,11.354002,10.323239,9.495506,8.663869,7.8361354,7.0044975,6.1767645,5.22409,4.2753205,3.3265507,2.3738766,1.4251068,2.2645533,3.1039999,3.9434462,4.786797,5.6262436,5.153811,4.6852827,4.2167544,3.7443218,3.2757936,5.2006636,7.125534,9.050405,10.975275,12.900145,14.50095,16.10566,17.706465,19.311174,20.911978,20.256039,19.596195,18.940256,18.284315,17.624472,18.089096,18.553719,19.018343,19.486872,19.951496,18.030529,16.113468,14.196406,12.2793455,10.362284,8.859089,7.355894,5.8566036,4.3534083,2.8502135,2.280171,1.7101282,1.1400855,0.5700427,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.78868926,1.5734742,2.3621633,3.1508527,3.9356375,3.7482262,3.5608149,3.3734035,3.1859922,2.998581,4.1620927,5.3256044,6.4891167,7.648724,8.812236,10.4637985,12.111456,13.763018,15.410676,17.062239,17.175465,17.288692,17.40192,17.511244,17.624472,14.313539,10.998701,7.687768,4.376835,1.0619974,0.8511597,0.63641757,0.42557985,0.21083772,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.8511597,1.698415,2.5495746,3.4007344,4.251894,4.8375545,5.423215,6.012779,6.5984397,7.1880045,6.5008297,5.813655,5.12648,4.4393053,3.7482262,4.911738,6.0752497,7.238762,8.398369,9.561881,9.874233,10.186585,10.498938,10.81129,11.123642,11.849861,12.576079,13.298394,14.024612,14.750832,16.69913,18.651329,20.599627,22.551826,24.500124,26.612406,28.724688,30.83697,32.94925,35.06153,35.237232,35.41293,35.588627,35.764324,35.93612,36.424168,36.91222,37.40027,37.88832,38.37637,37.876606,37.376842,36.873177,36.373413,35.87365,34.53834,33.19913,31.863827,30.524616,29.189312,26.510891,23.836376,21.16186,18.487345,15.812829,14.325252,12.837675,11.350098,9.86252,8.374943,6.8873653,5.3997884,3.912211,2.4246337,0.93705654,0.81211567,0.6871748,0.5622339,0.43729305,0.31235218,0.30063897,0.28892577,0.27330816,0.26159495,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.3513962,0.26159495,0.1756981,0.08589685,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.43729305,0.62470436,0.81211567,0.999527,1.1869383,0.9878138,0.78868926,0.58566034,0.38653582,0.18741131,0.47633708,0.76135844,1.0502841,1.33921,1.6242313,2.2372224,2.8502135,3.4632049,4.0761957,4.689187,4.548629,4.4119744,4.2753205,4.138666,3.998108,3.9629683,3.9239242,3.8887846,3.8497405,3.8106966,3.6506162,3.4866312,3.3265507,3.1625657,2.998581,3.2757936,3.5491016,3.8263142,4.0996222,4.376835,4.2870336,4.2011366,4.1113358,4.025439,3.9356375,3.951255,3.9629683,3.9746814,3.9863946,3.998108,3.5373883,3.076669,2.612045,2.1513257,1.6867018,2.1864653,2.6862288,3.1859922,3.6857557,4.1894236,3.6857557,3.1859922,2.6862288,2.1864653,1.6867018,2.0498111,2.4129205,2.77603,3.1391394,3.4983444,3.7247996,3.951255,4.173806,4.4002614,4.6267166,5.099149,5.575486,6.0518236,6.524256,7.000593,6.114294,5.22409,4.337791,3.4514916,2.5612879,2.0498111,1.5383345,1.0268579,0.5114767,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.1639849,0.26159495,0.3631094,0.46071947,0.5622339,0.48805028,0.41386664,0.3357786,0.26159495,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.24988174,0.31235218,0.37482262,0.43729305,0.4997635,0.8238289,1.1517987,1.475864,1.7999294,2.1239948,2.5495746,2.9751544,3.4007344,3.8263142,4.251894,4.263607,4.2753205,4.2870336,4.298747,4.3143644,4.025439,3.736513,3.4514916,3.1625657,2.87364,3.5256753,4.173806,4.825841,5.473972,6.126007,7.289519,8.449126,9.612638,10.77615,11.935758,12.037272,12.138786,12.236397,12.337912,12.439425,11.373524,10.311526,9.249529,8.187531,7.125534,5.735567,4.349504,2.9634414,1.5734742,0.18741131,1.0112402,1.8389735,2.6628022,3.4866312,4.3143644,3.9239242,3.5373883,3.1508527,2.7643168,2.3738766,4.3612175,6.348558,8.335898,10.323239,12.31058,14.575133,16.835783,19.100336,21.360985,23.625538,22.86418,22.098917,21.337559,20.5762,19.810938,20.361458,20.911978,21.4625,22.01302,22.563541,20.462973,18.362404,16.261835,14.161267,12.0606985,10.362284,8.663869,6.9615493,5.263134,3.5608149,2.8502135,2.135708,1.4251068,0.7106012,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.62860876,1.261122,1.8897307,2.5183394,3.1508527,2.998581,2.8502135,2.7018464,2.5495746,2.4012074,3.330455,4.2597027,5.1889505,6.1181984,7.0513506,8.371038,9.690726,11.010414,12.330102,13.64979,13.739592,13.829392,13.919194,14.008995,14.098797,11.4516115,8.800523,6.1494336,3.4983444,0.8511597,0.6910792,0.5309987,0.3709182,0.21083772,0.05075723,0.23426414,0.41386664,0.59737355,0.78088045,0.96438736,1.5969005,2.233318,2.8658314,3.5022488,4.138666,3.8575494,3.5764325,3.2992198,3.018103,2.736986,2.2957885,1.8584955,1.4172981,0.97610056,0.5388075,1.1088502,1.6827974,2.2567444,2.8267872,3.4007344,3.873167,4.349504,4.825841,5.298274,5.774611,5.22409,4.6735697,4.123049,3.5764325,3.0259118,3.959064,4.8883114,5.8214636,6.754616,7.687768,7.929841,8.171914,8.413987,8.65606,8.898132,9.479889,10.061645,10.639496,11.221252,11.799104,13.360865,14.92653,16.48829,18.05005,19.611813,21.396124,23.176533,24.960844,26.741251,28.525562,28.763731,28.997995,29.236164,29.474333,29.712502,30.263021,30.813543,31.364063,31.910679,32.4612,32.004387,31.54757,31.090755,30.63394,30.173222,29.119032,28.06094,27.002846,25.944754,24.88666,22.645533,20.404406,18.159374,15.918248,13.673217,12.419904,11.166591,9.909373,8.65606,7.3988423,6.36808,5.3412223,4.31046,3.279698,2.2489357,1.9912452,1.7296503,1.4719596,1.2103647,0.94876975,1.0112402,1.0698062,1.1283722,1.1908426,1.2494087,1.0190489,0.78478485,0.5544251,0.32016098,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.093705654,0.14055848,0.19131571,0.23816854,0.19131571,0.14055848,0.093705654,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14446288,0.21864653,0.28892577,0.3631094,0.28892577,0.21864653,0.14446288,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.05075723,0.093705654,0.13274968,0.1717937,0.21083772,0.38263142,0.5544251,0.7223144,0.8941081,1.0619974,0.96438736,0.8628729,0.76135844,0.6637484,0.5622339,0.8433509,1.1283722,1.4094892,1.6906061,1.9756275,2.5612879,3.1430438,3.7287042,4.3143644,4.900025,4.9468775,4.989826,5.036679,5.0796275,5.12648,4.927356,4.728231,4.533011,4.3338866,4.138666,3.8965936,3.6506162,3.408543,3.1664703,2.9243972,3.4046388,3.8848803,4.365122,4.845363,5.3256044,4.985922,4.650143,4.3143644,3.9746814,3.638903,3.795079,3.951255,4.1113358,4.267512,4.423688,3.998108,3.5764325,3.1508527,2.7252727,2.2996929,2.6042364,2.9087796,3.213323,3.521771,3.8263142,3.3655949,2.9048753,2.4441557,1.9834363,1.5266213,1.796025,2.069333,2.3426414,2.6159496,2.8892577,3.076669,3.2640803,3.4514916,3.638903,3.8263142,4.1972322,4.5681505,4.942973,5.3138914,5.688714,5.165524,4.646239,4.126953,3.6076677,3.0883822,2.7018464,2.3192148,1.9326792,1.5461433,1.1635119,1.0659018,0.97219616,0.8784905,0.78088045,0.6871748,0.5505207,0.41386664,0.27330816,0.13665408,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.10541886,0.09761006,0.08980125,0.08199245,0.07418364,0.15617609,0.23426414,0.31625658,0.39434463,0.47633708,0.41386664,0.3553006,0.29673457,0.23426414,0.1756981,0.14836729,0.12494087,0.10151446,0.07418364,0.05075723,0.058566034,0.07027924,0.078088045,0.08980125,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.015617609,0.023426414,0.027330816,0.031235218,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.042948425,0.046852827,0.046852827,0.05075723,0.08199245,0.113227665,0.14836729,0.1796025,0.21083772,0.25769055,0.30063897,0.3474918,0.39434463,0.43729305,0.6949836,0.95267415,1.2103647,1.4680552,1.7257458,2.0615244,2.4012074,2.736986,3.076669,3.4124475,3.4241607,3.4319696,3.4436827,3.4514916,3.4632049,3.240654,3.0220075,2.803361,2.5808098,2.3621633,2.87364,3.3812122,3.892689,4.4041657,4.911738,5.840986,6.7663293,7.6955767,8.62092,9.550168,9.628256,9.710248,9.788337,9.870329,9.948417,9.101162,8.250002,7.3988423,6.551587,5.700427,4.630621,3.5647192,2.4988174,1.4290112,0.3631094,0.9917182,1.6242313,2.25284,2.8814487,3.513962,3.2836022,3.0532427,2.822883,2.592523,2.3621633,3.9356375,5.5091114,7.0786815,8.652155,10.22563,12.138786,14.055848,15.969006,17.886066,19.799223,19.865599,19.935879,20.002253,20.068628,20.138906,20.517633,20.89636,21.278992,21.657719,22.036446,20.053009,18.073479,16.090042,14.106606,12.123169,10.639496,9.155824,7.6682463,6.184573,4.7009,3.775557,2.8502135,1.9248703,0.999527,0.07418364,0.06637484,0.05466163,0.046852827,0.03513962,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.47243267,0.94486535,1.4172981,1.8897307,2.3621633,2.2489357,2.135708,2.0263848,1.9131571,1.7999294,2.4988174,3.193801,3.892689,4.591577,5.2865605,6.278279,7.266093,8.257811,9.245625,10.237343,10.303718,10.373997,10.4403715,10.506746,10.573121,8.58578,6.5984397,4.6110992,2.6237583,0.63641757,0.5309987,0.42167544,0.31625658,0.20693332,0.10151446,0.46462387,0.8316377,1.1947471,1.5617609,1.9248703,3.193801,4.466636,5.735567,7.0044975,8.273428,7.715099,7.1567693,6.5945354,6.036206,5.473972,4.5954814,3.716991,2.8345962,1.9561055,1.0737107,1.3704453,1.6632754,1.9600099,2.2567444,2.5495746,2.912684,3.2757936,3.638903,3.998108,4.3612175,3.951255,3.5373883,3.1235218,2.7135596,2.2996929,3.0024853,3.7052777,4.40807,5.1108627,5.813655,5.985449,6.1572423,6.329036,6.5008297,6.676528,7.1099167,7.5433054,7.9805984,8.413987,8.85128,10.0265045,11.20173,12.376955,13.548276,14.723501,16.175938,17.628376,19.080814,20.53325,21.98569,22.286327,22.586967,22.887606,23.188246,23.488884,24.101875,24.710962,25.323954,25.936945,26.549934,26.136068,25.718298,25.304432,24.890564,24.476698,23.695818,22.91884,22.141865,21.36489,20.587914,18.77627,16.968533,15.15689,13.349152,11.537509,10.514555,9.491602,8.468649,7.445695,6.426646,5.852699,5.278752,4.7087092,4.134762,3.5608149,3.1664703,2.7721257,2.377781,1.9834363,1.5890918,1.7218413,1.8506867,1.9834363,2.1161861,2.2489357,1.8350691,1.4212024,1.0034313,0.58956474,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.093705654,0.19131571,0.28502136,0.37872702,0.47633708,0.37872702,0.28502136,0.19131571,0.093705654,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.113227665,0.1717937,0.23035973,0.28892577,0.23035973,0.1717937,0.113227665,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.05466163,0.08589685,0.113227665,0.14446288,0.1756981,0.3279698,0.48024148,0.63251317,0.78478485,0.93705654,0.93705654,0.93705654,0.93705654,0.93705654,0.93705654,1.2142692,1.4914817,1.7686942,2.0459068,2.3231194,2.8814487,3.4397783,3.998108,4.5564375,5.1108627,5.3412223,5.5676775,5.794133,6.0205884,6.250948,5.891743,5.5364423,5.1772375,4.8219366,4.462732,4.138666,3.8185053,3.49444,3.174279,2.8502135,3.533484,4.220659,4.903929,5.591104,6.2743745,5.688714,5.099149,4.513489,3.9239242,3.338264,3.638903,3.9434462,4.2440853,4.548629,4.8492675,4.462732,4.0761957,3.6857557,3.2992198,2.912684,3.0220075,3.1313305,3.240654,3.3538816,3.4632049,3.0415294,2.6237583,2.2020829,1.7843118,1.3626363,1.5461433,1.7257458,1.9092526,2.0927596,2.2762666,2.4246337,2.5769055,2.7252727,2.87364,3.0259118,3.2953155,3.5647192,3.8341231,4.1035266,4.376835,4.220659,4.068387,3.9161155,3.7638438,3.611572,3.3538816,3.096191,2.8385005,2.5808098,2.3231194,2.135708,1.9443923,1.7530766,1.5656652,1.3743496,1.1010414,0.8238289,0.5505207,0.27330816,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.09761006,0.093705654,0.093705654,0.08980125,0.08589685,0.14836729,0.20693332,0.26940376,0.3279698,0.38653582,0.3435874,0.29673457,0.25378615,0.20693332,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.039044023,0.046852827,0.05075723,0.058566034,0.06637484,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.03513962,0.046852827,0.05466163,0.06637484,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.078088045,0.08589685,0.08980125,0.093705654,0.10151446,0.12884527,0.15617609,0.1835069,0.21083772,0.23816854,0.26549935,0.29283017,0.32016098,0.3474918,0.37482262,0.5661383,0.75354964,0.94486535,1.1361811,1.3235924,1.5734742,1.8233559,2.0732377,2.3231194,2.5769055,2.5808098,2.5886188,2.5964274,2.6042364,2.612045,2.4597735,2.3075018,2.15523,2.0029583,1.8506867,2.2216048,2.5886188,2.959537,3.330455,3.7013733,4.3924527,5.083532,5.7785153,6.4695945,7.1606736,7.223144,7.28171,7.3441806,7.4027467,7.461313,6.824895,6.1884775,5.548156,4.911738,4.2753205,3.5256753,2.7799344,2.0341935,1.2845483,0.5388075,0.97219616,1.4055848,1.8428779,2.2762666,2.7135596,2.639376,2.5690966,2.494913,2.4207294,2.35045,3.506153,4.6657605,5.8214636,6.9810715,8.136774,9.706344,11.272009,12.841579,14.407245,15.976814,16.870922,17.768934,18.666946,19.56496,20.462973,20.67381,20.880743,21.091581,21.302418,21.513256,19.646952,17.780647,15.918248,14.051944,12.185639,10.916709,9.647778,8.378847,7.1060123,5.8370814,4.7009,3.5608149,2.4246337,1.2884527,0.14836729,0.12884527,0.10932326,0.08980125,0.07027924,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.31625658,0.62860876,0.94486535,1.261122,1.5734742,1.4992905,1.4251068,1.3509232,1.2767396,1.1986516,1.6632754,2.1318035,2.5964274,3.0610514,3.5256753,4.185519,4.845363,5.505207,6.165051,6.824895,6.871748,6.914696,6.9615493,7.0044975,7.0513506,5.7238536,4.4002614,3.076669,1.7491722,0.42557985,0.3709182,0.31625658,0.26159495,0.20693332,0.14836729,0.698888,1.2455044,1.7921207,2.338737,2.8892577,4.7907014,6.6960497,8.601398,10.506746,12.412095,11.572648,10.733202,9.893755,9.054309,8.210958,6.89127,5.571582,4.251894,2.9322062,1.6125181,1.6281357,1.6476578,1.6632754,1.6827974,1.698415,1.9482968,2.1981785,2.4519646,2.7018464,2.951728,2.6745155,2.4012074,2.1239948,1.8506867,1.5734742,2.0459068,2.5183394,2.9907722,3.4632049,3.9356375,4.041056,4.142571,4.2440853,4.3455997,4.4510183,4.7399445,5.02887,5.3217,5.610626,5.899552,6.688241,7.47693,8.261715,9.050405,9.839094,10.959657,12.084125,13.204688,14.329156,15.449719,15.812829,16.175938,16.539047,16.898252,17.261362,17.936825,18.612286,19.287746,19.96321,20.63867,20.263847,19.89293,19.518106,19.147188,18.77627,18.276506,17.780647,17.280884,16.785025,16.289165,14.9109125,13.532659,12.154405,10.77615,9.4018,8.609207,7.8205175,7.0318284,6.239235,5.4505453,5.3334136,5.2201858,5.1030536,4.989826,4.8765984,4.3455997,3.814601,3.2836022,2.7565079,2.2255092,2.4285383,2.6354716,2.8385005,3.0454338,3.2484627,2.6510892,2.0537157,1.456342,0.8589685,0.26159495,0.21083772,0.15617609,0.10541886,0.05075723,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14055848,0.28502136,0.42557985,0.5700427,0.7106012,0.5700427,0.42557985,0.28502136,0.14055848,0.0,0.0,0.0,0.0,0.0,0.0,0.042948425,0.08589685,0.12884527,0.1717937,0.21083772,0.1717937,0.12884527,0.08589685,0.042948425,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.058566034,0.078088045,0.09761006,0.11713207,0.13665408,0.27330816,0.40605783,0.5427119,0.679366,0.81211567,0.9136301,1.0112402,1.1127546,1.2142692,1.3118792,1.5851873,1.8584955,2.1318035,2.4012074,2.6745155,3.2055142,3.736513,4.263607,4.794606,5.3256044,5.735567,6.1455293,6.5554914,6.9654536,7.375416,6.8561306,6.3407493,5.8214636,5.3060827,4.786797,4.3846436,3.9824903,3.5803368,3.1781836,2.77603,3.6662338,4.5564375,5.446641,6.336845,7.223144,6.387602,5.548156,4.7126136,3.873167,3.0376248,3.4866312,3.9317331,4.380739,4.825841,5.2748475,4.9234514,4.575959,4.224563,3.873167,3.5256753,3.4397783,3.3538816,3.2718892,3.1859922,3.1000953,2.7213683,2.338737,1.9600099,1.5812829,1.1986516,1.2923572,1.3860629,1.475864,1.5695697,1.6632754,1.7765031,1.8858263,1.999054,2.1122816,2.2255092,2.3933985,2.5612879,2.7291772,2.893162,3.0610514,3.2757936,3.49444,3.7091823,3.9239242,4.138666,4.0059166,3.8770714,3.7482262,3.619381,3.4866312,3.2016098,2.9165885,2.631567,2.3465457,2.0615244,1.6515622,1.2376955,0.8238289,0.41386664,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.08980125,0.093705654,0.093705654,0.09761006,0.10151446,0.14055848,0.1796025,0.21864653,0.26159495,0.30063897,0.26940376,0.23816854,0.21083772,0.1796025,0.14836729,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.031235218,0.03513962,0.039044023,0.046852827,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.05075723,0.06637484,0.08199245,0.09761006,0.113227665,0.113227665,0.113227665,0.113227665,0.113227665,0.113227665,0.12103647,0.12884527,0.13665408,0.14055848,0.14836729,0.1717937,0.19522011,0.21864653,0.23816854,0.26159495,0.27330816,0.28111696,0.29283017,0.30063897,0.31235218,0.43338865,0.5583295,0.679366,0.80430686,0.92534333,1.0893283,1.2494087,1.4133936,1.5734742,1.737459,1.7413634,1.7491722,1.7530766,1.756981,1.7608855,1.678893,1.5929961,1.5070993,1.4212024,1.33921,1.5656652,1.796025,2.0263848,2.2567444,2.4871042,2.9439192,3.4007344,3.8614538,4.318269,4.775084,4.814128,4.853172,4.8961205,4.9351645,4.9742084,4.548629,4.126953,3.7013733,3.2757936,2.8502135,2.4207294,1.9951496,1.5656652,1.1400855,0.7106012,0.95267415,1.1908426,1.4329157,1.6710842,1.9131571,1.999054,2.0810463,2.1669433,2.25284,2.338737,3.0805733,3.8224099,4.564246,5.3060827,6.0518236,7.269997,8.488171,9.710248,10.928422,12.150499,13.8762455,15.605896,17.331642,19.061293,20.787037,20.826082,20.86903,20.908073,20.947119,20.986162,19.240894,17.491722,15.746454,13.997282,12.24811,11.193921,10.139732,9.085544,8.031356,6.9732623,5.6262436,4.2753205,2.9243972,1.5734742,0.22645533,0.19522011,0.1639849,0.13665408,0.10541886,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15617609,0.31625658,0.47243267,0.62860876,0.78868926,0.74964523,0.7106012,0.6754616,0.63641757,0.60127795,0.8316377,1.0659018,1.2962615,1.5305257,1.7608855,2.0927596,2.4207294,2.7526035,3.0805733,3.4124475,3.435874,3.4593005,3.4788225,3.5022488,3.5256753,2.8619268,2.1981785,1.5383345,0.8745861,0.21083772,0.21083772,0.20693332,0.20693332,0.20302892,0.19912452,0.92924774,1.6593709,2.3894942,3.1196175,3.8497405,6.3915067,8.929368,11.471134,14.008995,16.55076,15.430198,14.309634,13.189071,12.068507,10.951848,9.190963,7.4300776,5.6691923,3.9083066,2.1513257,1.8897307,1.6281357,1.3704453,1.1088502,0.8511597,0.9878138,1.1244678,1.261122,1.4016805,1.5383345,1.4016805,1.261122,1.1244678,0.9878138,0.8511597,1.0932326,1.3353056,1.5773785,1.8194515,2.0615244,2.096664,2.1278992,2.1591344,2.194274,2.2255092,2.3699722,2.514435,2.6588979,2.803361,2.951728,3.349977,3.7482262,4.1503797,4.548629,4.950782,5.743376,6.5359693,7.328563,8.121157,8.913751,9.339331,9.761005,10.186585,10.612165,11.037745,11.775677,12.513609,13.251541,13.985569,14.723501,14.395531,14.063657,13.735687,13.403813,13.075843,12.857197,12.63855,12.423808,12.205161,11.986515,11.04165,10.096785,9.151918,8.207053,7.262188,6.703859,6.1494336,5.591104,5.0327744,4.474445,4.8180323,5.1616197,5.5013027,5.84489,6.1884775,5.520825,4.8570766,4.193328,3.5256753,2.8619268,3.1391394,3.416352,3.6935644,3.970777,4.251894,3.4710135,2.690133,1.9092526,1.1283722,0.3513962,0.28111696,0.21083772,0.14055848,0.07027924,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19131571,0.37872702,0.5700427,0.76135844,0.94876975,0.76135844,0.5700427,0.37872702,0.19131571,0.0,0.0,0.0,0.0,0.0,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.10932326,0.08199245,0.05466163,0.027330816,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.058566034,0.07027924,0.078088045,0.08980125,0.10151446,0.21864653,0.3357786,0.45291066,0.5700427,0.6871748,0.8862993,1.0893283,1.2884527,1.4875772,1.6867018,1.9561055,2.2216048,2.4910088,2.7565079,3.0259118,3.5256753,4.029343,4.533011,5.036679,5.5364423,6.1299114,6.7233806,7.3168497,7.9064145,8.499884,7.824422,7.1450562,6.46569,5.7902284,5.1108627,4.630621,4.1464753,3.6662338,3.182088,2.7018464,3.795079,4.8883114,5.985449,7.0786815,8.175818,7.08649,6.001066,4.911738,3.8263142,2.736986,3.330455,3.9239242,4.513489,5.1069584,5.700427,5.388075,5.0757227,4.7633705,4.4510183,4.138666,3.8575494,3.5764325,3.2992198,3.018103,2.736986,2.397303,2.05762,1.717937,1.3782539,1.038571,1.038571,1.0424755,1.0463798,1.0463798,1.0502841,1.1244678,1.1986516,1.2767396,1.3509232,1.4251068,1.4914817,1.5539521,1.620327,1.6867018,1.7491722,2.330928,2.9165885,3.4983444,4.0801005,4.661856,4.661856,4.657952,4.6540475,4.6540475,4.650143,4.271416,3.8887846,3.5100577,3.1313305,2.7486992,2.1981785,1.6515622,1.1010414,0.5505207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.08199245,0.08980125,0.09761006,0.10541886,0.113227665,0.13274968,0.15227169,0.1717937,0.19131571,0.21083772,0.19912452,0.1835069,0.1678893,0.15227169,0.13665408,0.113227665,0.08589685,0.062470436,0.039044023,0.011713207,0.015617609,0.015617609,0.019522011,0.023426414,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.07027924,0.08980125,0.10932326,0.12884527,0.14836729,0.14836729,0.14836729,0.14836729,0.14836729,0.14836729,0.16008049,0.1717937,0.1796025,0.19131571,0.19912452,0.21864653,0.23426414,0.25378615,0.26940376,0.28892577,0.28111696,0.27330816,0.26549935,0.25769055,0.24988174,0.30454338,0.359205,0.41386664,0.46852827,0.5231899,0.60127795,0.6754616,0.74964523,0.8238289,0.9019169,0.9019169,0.9058213,0.9058213,0.9097257,0.9136301,0.8941081,0.8784905,0.8589685,0.8433509,0.8238289,0.9136301,1.0034313,1.0932326,1.183034,1.2767396,1.4992905,1.7218413,1.9443923,2.1630387,2.3855898,2.4090161,2.4285383,2.4480603,2.4675822,2.4871042,2.2762666,2.0615244,1.8506867,1.6359446,1.4251068,1.3157835,1.2103647,1.1010414,0.9956226,0.8862993,0.93315214,0.97610056,1.0229534,1.0659018,1.1127546,1.3548276,1.5969005,1.8389735,2.0810463,2.3231194,2.6510892,2.979059,3.3070288,3.6349986,3.9629683,4.83365,5.708236,6.578918,7.453504,8.324185,10.881569,13.438952,15.996336,18.553719,21.111103,20.982258,20.853413,20.720663,20.591818,20.462973,18.830933,17.202797,15.570756,13.94262,12.31058,11.471134,10.631687,9.792241,8.952794,8.113348,6.551587,4.985922,3.4241607,1.8623998,0.30063897,0.26159495,0.21864653,0.1796025,0.14055848,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,1.1635119,2.0732377,2.9868677,3.900498,4.814128,7.988407,11.162686,14.336966,17.511244,20.689428,19.287746,17.886066,16.48829,15.086611,13.688834,11.486752,9.288573,7.08649,4.8883114,2.6862288,2.1513257,1.6125181,1.0737107,0.5388075,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.5231899,0.9878138,1.4485333,1.9131571,2.3738766,2.8619268,3.349977,3.8380275,4.3260775,4.814128,5.610626,6.4110284,7.211431,8.011833,8.812236,8.52331,8.238289,7.9493628,7.6643414,7.375416,7.437886,7.5003567,7.562827,7.6252975,7.687768,7.1762915,6.66091,6.1494336,5.6379566,5.12648,4.7985106,4.474445,4.1503797,3.8263142,3.4983444,4.298747,5.099149,5.899552,6.699954,7.5003567,6.699954,5.899552,5.099149,4.298747,3.4983444,3.8497405,4.2011366,4.548629,4.900025,5.251421,4.2870336,3.3265507,2.3621633,1.4016805,0.43729305,0.3513962,0.26159495,0.1756981,0.08589685,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23816854,0.47633708,0.7106012,0.94876975,1.1869383,0.94876975,0.7106012,0.47633708,0.23816854,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.1639849,0.26159495,0.3631094,0.46071947,0.5622339,0.8628729,1.1635119,1.4641509,1.7608855,2.0615244,2.3231194,2.5886188,2.8502135,3.1118085,3.3734035,3.8497405,4.3260775,4.7985106,5.2748475,5.7511845,6.524256,7.3012323,8.074304,8.85128,9.6243515,8.78881,7.9493628,7.113821,6.2743745,5.4388323,4.8765984,4.3143644,3.7482262,3.1859922,2.6237583,3.9239242,5.22409,6.524256,7.824422,9.124588,7.7892823,6.4500723,5.1108627,3.775557,2.436347,3.174279,3.912211,4.650143,5.388075,6.126007,5.8487945,5.575486,5.298274,5.024966,4.7516575,4.2753205,3.7989833,3.3265507,2.8502135,2.3738766,2.0732377,1.7765031,1.475864,1.175225,0.8745861,0.78868926,0.698888,0.61299115,0.5231899,0.43729305,0.47633708,0.5114767,0.5505207,0.58566034,0.62470436,0.58566034,0.5505207,0.5114767,0.47633708,0.43729305,1.3860629,2.338737,3.2875066,4.2362766,5.1889505,5.3138914,5.4388323,5.563773,5.688714,5.813655,5.337318,4.860981,4.388548,3.912211,3.435874,2.7486992,2.0615244,1.3743496,0.6871748,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,0.26159495,0.27330816,0.28892577,0.30063897,0.31235218,0.28892577,0.26159495,0.23816854,0.21083772,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.113227665,0.1639849,0.21083772,0.26159495,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21083772,0.42557985,0.63641757,0.8511597,1.0619974,0.9136301,0.76135844,0.61299115,0.46071947,0.31235218,0.7106012,1.1127546,1.5110037,1.9131571,2.3114061,2.2255092,2.135708,2.0498111,1.9639144,1.8741131,2.4012074,2.9243972,3.4514916,3.9746814,4.5017757,7.8868923,11.275913,14.661031,18.05005,21.439074,21.138433,20.837795,20.537155,20.236517,19.935879,18.424873,16.91387,15.398962,13.887959,12.373051,11.748346,11.123642,10.498938,9.874233,9.249529,7.473026,5.700427,3.9239242,2.1513257,0.37482262,0.3240654,0.27330816,0.22645533,0.1756981,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.92924774,1.6593709,2.3894942,3.1196175,3.8497405,6.3915067,8.929368,11.471134,14.008995,16.55076,15.430198,14.309634,13.189071,12.068507,10.951848,9.190963,7.4300776,5.6691923,3.9083066,2.1513257,1.7218413,1.2884527,0.8589685,0.42948425,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10932326,0.12103647,0.12884527,0.14055848,0.14836729,0.12103647,0.093705654,0.06637484,0.039044023,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.019522011,0.027330816,0.03513962,0.042948425,0.05075723,0.42167544,0.78868926,1.1596074,1.5305257,1.901444,2.2918842,2.67842,3.06886,3.4593005,3.8497405,4.4900627,5.1303844,5.7707067,6.4110284,7.0513506,6.8209906,6.590631,6.3602715,6.1299114,5.899552,5.9542136,6.008875,6.0635366,6.1181984,6.1767645,5.794133,5.4154058,5.036679,4.6540475,4.2753205,4.1308575,3.9863946,3.8419318,3.6935644,3.5491016,4.4588275,5.364649,6.2743745,7.180196,8.086017,7.230953,6.3719845,5.5169206,4.657952,3.7989833,4.01763,4.2362766,4.4510183,4.6696653,4.8883114,4.025439,3.1625657,2.2996929,1.43682,0.57394713,0.46071947,0.3435874,0.23035973,0.113227665,0.0,0.0,0.0,0.0,0.0,0.0,0.15617609,0.30844778,0.46462387,0.62079996,0.77307165,0.8160201,0.8589685,0.9019169,0.94486535,0.9878138,1.0268579,1.0659018,1.1088502,1.1478943,1.1869383,1.4992905,1.8077383,2.1161861,2.4285383,2.736986,2.397303,2.05762,1.717937,1.3782539,1.038571,0.8316377,0.62860876,0.42167544,0.21864653,0.011713207,0.015617609,0.023426414,0.027330816,0.031235218,0.039044023,0.046852827,0.058566034,0.06637484,0.078088045,0.08589685,0.093705654,0.09761006,0.10151446,0.10932326,0.113227665,0.093705654,0.07418364,0.05075723,0.031235218,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.19131571,0.37872702,0.5700427,0.76135844,0.94876975,0.76916724,0.58566034,0.40215343,0.21864653,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.078088045,0.12103647,0.1639849,0.20693332,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.031235218,0.03513962,0.039044023,0.046852827,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.12884527,0.21083772,0.28892577,0.3709182,0.44900626,0.75745404,1.0659018,1.3743496,1.678893,1.9873407,2.182561,2.377781,2.5730011,2.7682211,2.9634414,3.2914112,3.6232853,3.951255,4.283129,4.6110992,5.298274,5.989353,6.676528,7.363703,8.050878,7.3597984,6.6687193,5.9815445,5.290465,4.5993857,4.154284,3.7052777,3.2562714,2.8111696,2.3621633,3.349977,4.337791,5.3256044,6.3134184,7.3012323,6.902983,6.504734,6.1064854,5.708236,5.3138914,5.4115014,5.5091114,5.606722,5.704332,5.801942,5.434928,5.0718184,4.704805,4.3416953,3.9746814,3.611572,3.2445583,2.8814487,2.514435,2.1513257,1.8702087,1.5890918,1.3118792,1.0307622,0.74964523,0.6715572,0.58956474,0.5114767,0.42948425,0.3513962,0.37872702,0.40996224,0.44119745,0.46852827,0.4997635,0.48805028,0.48024148,0.46852827,0.46071947,0.44900626,1.2064602,1.9639144,2.7213683,3.4788225,4.2362766,4.3260775,4.4119744,4.5017757,4.5876727,4.6735697,4.298747,3.9239242,3.5491016,3.174279,2.7994564,2.241127,1.678893,1.1205635,0.5583295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.058566034,0.07027924,0.078088045,0.08980125,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.08980125,0.11713207,0.14446288,0.1717937,0.19912452,0.21083772,0.21864653,0.23035973,0.23816854,0.24988174,0.25769055,0.26549935,0.27330816,0.28111696,0.28892577,0.30063897,0.31625658,0.3318742,0.3474918,0.3631094,0.3513962,0.3357786,0.3240654,0.31235218,0.30063897,0.29283017,0.28502136,0.27721256,0.26940376,0.26159495,0.22645533,0.19131571,0.15617609,0.12103647,0.08589685,0.078088045,0.07418364,0.06637484,0.058566034,0.05075723,0.093705654,0.13665408,0.1756981,0.21864653,0.26159495,0.22645533,0.19131571,0.15617609,0.12103647,0.08589685,0.07418364,0.058566034,0.042948425,0.027330816,0.011713207,0.019522011,0.027330816,0.03513962,0.042948425,0.05075723,0.07418364,0.093705654,0.11713207,0.14055848,0.1639849,0.3709182,0.57785153,0.78478485,0.9917182,1.1986516,1.0854238,0.96829176,0.8550641,0.7418364,0.62470436,0.8784905,1.1361811,1.3899672,1.6437533,1.901444,1.8428779,1.7843118,1.7257458,1.6710842,1.6125181,2.2098918,2.8072653,3.4046388,4.0020123,4.5993857,7.125534,9.651682,12.173926,14.700074,17.226223,16.968533,16.714746,16.46096,16.20327,15.949483,14.774258,13.599033,12.423808,11.248583,10.073358,9.554072,9.034787,8.515501,7.996216,7.473026,6.0479193,4.618908,3.193801,1.7647898,0.3357786,0.29283017,0.24597734,0.20302892,0.15617609,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.698888,1.2455044,1.7921207,2.338737,2.8892577,4.7907014,6.6960497,8.601398,10.506746,12.412095,11.572648,10.733202,9.893755,9.054309,8.210958,6.89127,5.571582,4.251894,2.9322062,1.6125181,1.2884527,0.96829176,0.6442264,0.3240654,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.08199245,0.08980125,0.09761006,0.10541886,0.113227665,0.093705654,0.078088045,0.058566034,0.042948425,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.027330816,0.031235218,0.031235218,0.03513962,0.039044023,0.31625658,0.59346914,0.8706817,1.1478943,1.4251068,1.717937,2.0107672,2.3035975,2.5964274,2.8892577,3.3655949,3.8458362,4.3260775,4.806319,5.2865605,5.114767,4.942973,4.7711797,4.5993857,4.423688,4.4705405,4.521298,4.5681505,4.6150036,4.661856,4.415879,4.165997,3.9200199,3.6740425,3.4241607,3.4593005,3.49444,3.5295796,3.5647192,3.5998588,4.6150036,5.630148,6.6452928,7.660437,8.675582,7.7619514,6.844417,5.930787,5.0132523,4.0996222,4.185519,4.271416,4.3534083,4.4393053,4.5252023,3.7638438,2.998581,2.2372224,1.475864,0.7106012,0.5700427,0.42557985,0.28502136,0.14055848,0.0,0.0,0.0,0.0,0.0,0.0,0.30844778,0.62079996,0.92924774,1.2415999,1.5500476,1.6359446,1.7218413,1.8038338,1.8897307,1.9756275,2.0537157,2.135708,2.2137961,2.2957885,2.3738766,2.9946766,3.6154766,4.2362766,4.853172,5.473972,4.794606,4.11524,3.435874,2.7565079,2.0732377,1.6632754,1.2533131,0.8433509,0.43338865,0.023426414,0.03513962,0.046852827,0.05466163,0.06637484,0.07418364,0.093705654,0.113227665,0.13665408,0.15617609,0.1756981,0.1835069,0.19522011,0.20693332,0.21474212,0.22645533,0.1835069,0.14446288,0.10541886,0.06637484,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.14055848,0.28502136,0.42557985,0.5700427,0.7106012,0.58566034,0.45681506,0.3318742,0.20302892,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.14836729,0.21864653,0.29283017,0.3631094,0.43729305,0.3513962,0.26159495,0.1756981,0.08589685,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.046852827,0.046852827,0.042948425,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.09761006,0.15617609,0.21864653,0.27721256,0.3357786,0.6520352,0.96829176,1.2806439,1.5969005,1.9131571,2.0380979,2.1669433,2.2957885,2.4207294,2.5495746,2.7330816,2.920493,3.1039999,3.2914112,3.474918,4.0761957,4.6735697,5.2748475,5.8761253,6.473499,5.930787,5.388075,4.8492675,4.3065557,3.7638438,3.4280653,3.096191,2.7643168,2.4324427,2.1005683,2.77603,3.4514916,4.126953,4.7985106,5.473972,6.016684,6.559396,7.1021075,7.6448197,8.187531,7.6448197,7.1021075,6.559396,6.016684,5.473972,5.0210614,4.564246,4.1113358,3.6545205,3.2016098,2.9439192,2.690133,2.436347,2.1786566,1.9248703,1.6632754,1.4055848,1.1439898,0.8862993,0.62470436,0.5544251,0.48024148,0.40605783,0.3357786,0.26159495,0.28502136,0.30844778,0.3318742,0.3513962,0.37482262,0.39434463,0.40996224,0.42557985,0.44510186,0.46071947,1.0268579,1.5929961,2.1591344,2.7213683,3.2875066,3.338264,3.3890212,3.435874,3.4866312,3.5373883,3.2640803,2.9868677,2.7135596,2.436347,2.1630387,1.7296503,1.2962615,0.8667773,0.43338865,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.046852827,0.05075723,0.058566034,0.06637484,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.093705654,0.12103647,0.15227169,0.1835069,0.21083772,0.23426414,0.25378615,0.27330816,0.29283017,0.31235218,0.31625658,0.31625658,0.32016098,0.3240654,0.3240654,0.3435874,0.359205,0.37872702,0.39434463,0.41386664,0.41386664,0.41386664,0.41386664,0.41386664,0.41386664,0.40996224,0.40605783,0.40605783,0.40215343,0.39824903,0.3435874,0.28502136,0.22645533,0.1717937,0.113227665,0.09761006,0.08199245,0.06637484,0.05075723,0.039044023,0.07418364,0.10932326,0.14055848,0.1756981,0.21083772,0.19131571,0.1717937,0.15227169,0.13274968,0.113227665,0.093705654,0.078088045,0.058566034,0.042948425,0.023426414,0.039044023,0.05466163,0.07027924,0.08589685,0.10151446,0.14446288,0.19131571,0.23426414,0.28111696,0.3240654,0.5270943,0.7301232,0.93315214,1.1361811,1.33921,1.2572175,1.1791295,1.097137,1.0190489,0.93705654,1.0463798,1.1557031,1.2689307,1.3782539,1.4875772,1.4602464,1.4329157,1.4055848,1.3782539,1.3509232,2.018576,2.690133,3.3616903,4.029343,4.7009,6.364176,8.023546,9.686822,11.350098,13.013372,12.802535,12.591698,12.380859,12.173926,11.963089,11.123642,10.2881,9.448653,8.6131115,7.773665,7.3597984,6.9459314,6.5281606,6.114294,5.700427,4.618908,3.541293,2.4597735,1.3782539,0.30063897,0.26159495,0.21864653,0.1796025,0.14055848,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.46462387,0.8316377,1.1947471,1.5617609,1.9248703,3.193801,4.466636,5.735567,7.0044975,8.273428,7.715099,7.1567693,6.5945354,6.036206,5.473972,4.5954814,3.716991,2.8345962,1.9561055,1.0737107,0.8589685,0.6442264,0.42948425,0.21474212,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05466163,0.058566034,0.06637484,0.07027924,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.03513962,0.031235218,0.031235218,0.027330816,0.023426414,0.21083772,0.39434463,0.58175594,0.76526284,0.94876975,1.1439898,1.33921,1.53443,1.7296503,1.9248703,2.2450314,2.5651922,2.8853533,3.2055142,3.5256753,3.408543,3.2953155,3.1781836,3.0649557,2.951728,2.9907722,3.0298162,3.06886,3.1118085,3.1508527,3.0337205,2.920493,2.803361,2.690133,2.5769055,2.7916477,3.0063896,3.2211318,3.435874,3.6506162,4.7711797,5.8956475,7.016211,8.140678,9.261242,8.289046,7.3168497,6.3446536,5.3724575,4.4002614,4.3534083,4.3065557,4.2557983,4.2089458,4.1620927,3.4983444,2.8385005,2.174752,1.5110037,0.8511597,0.679366,0.5114767,0.339683,0.1717937,0.0,0.0,0.0,0.0,0.0,0.0,0.46462387,0.92924774,1.3938715,1.8584955,2.3231194,2.4519646,2.5808098,2.7057507,2.8345962,2.9634414,3.0805733,3.2016098,3.3226464,3.4436827,3.5608149,4.493967,5.423215,6.3524623,7.28171,8.210958,7.191909,6.17286,5.153811,4.1308575,3.1118085,2.4988174,1.8819219,1.2689307,0.6520352,0.039044023,0.05075723,0.06637484,0.08199245,0.09761006,0.113227665,0.14055848,0.1717937,0.20302892,0.23426414,0.26159495,0.27721256,0.29283017,0.30844778,0.3240654,0.3357786,0.27721256,0.21864653,0.15617609,0.09761006,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.093705654,0.19131571,0.28502136,0.37872702,0.47633708,0.40215343,0.3318742,0.25769055,0.1835069,0.113227665,0.113227665,0.113227665,0.113227665,0.113227665,0.113227665,0.21474212,0.31625658,0.42167544,0.5231899,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.06637484,0.05466163,0.046852827,0.03513962,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.06637484,0.10541886,0.14446288,0.1835069,0.22645533,0.5466163,0.8706817,1.1908426,1.5149081,1.8389735,1.8975395,1.9561055,2.018576,2.077142,2.135708,2.1786566,2.2177005,2.2567444,2.2957885,2.338737,2.8502135,3.3616903,3.873167,4.388548,4.900025,4.50568,4.1113358,3.7130866,3.3187418,2.9243972,2.7057507,2.4910088,2.2723622,2.0537157,1.8389735,2.1981785,2.5612879,2.9243972,3.2875066,3.6506162,5.134289,6.6140575,8.097731,9.581403,11.061172,9.878138,8.699008,7.5159745,6.3329406,5.1499066,4.60329,4.0605783,3.513962,2.97125,2.4246337,2.280171,2.135708,1.9912452,1.8467822,1.698415,1.4602464,1.2181735,0.98000497,0.7418364,0.4997635,0.43338865,0.3709182,0.30454338,0.23816854,0.1756981,0.19131571,0.20693332,0.21864653,0.23426414,0.24988174,0.29673457,0.339683,0.38653582,0.42948425,0.47633708,0.8472553,1.2181735,1.5929961,1.9639144,2.338737,2.35045,2.3621633,2.3738766,2.3855898,2.4012074,2.2255092,2.0498111,1.8741131,1.698415,1.5266213,1.2181735,0.9136301,0.60908675,0.30454338,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.031235218,0.03513962,0.039044023,0.046852827,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.093705654,0.12884527,0.16008049,0.19131571,0.22645533,0.25378615,0.28502136,0.31625658,0.3435874,0.37482262,0.3709182,0.3709182,0.3670138,0.3631094,0.3631094,0.38263142,0.40215343,0.42167544,0.44119745,0.46071947,0.47633708,0.48805028,0.4997635,0.5114767,0.5231899,0.5270943,0.5309987,0.5309987,0.5349031,0.5388075,0.45681506,0.37872702,0.29673457,0.21864653,0.13665408,0.113227665,0.093705654,0.07027924,0.046852827,0.023426414,0.05075723,0.078088045,0.10932326,0.13665408,0.1639849,0.15617609,0.15227169,0.14836729,0.14055848,0.13665408,0.11713207,0.09761006,0.078088045,0.058566034,0.039044023,0.058566034,0.08199245,0.10541886,0.12884527,0.14836729,0.21864653,0.28502136,0.3513962,0.42167544,0.48805028,0.6832704,0.8823949,1.0815194,1.2767396,1.475864,1.4290112,1.3860629,1.33921,1.2962615,1.2494087,1.2142692,1.1791295,1.1439898,1.1088502,1.0737107,1.077615,1.0815194,1.0815194,1.0854238,1.0893283,1.8311646,2.5730011,3.3148375,4.056674,4.7985106,5.5989127,6.3993154,7.1997175,8.00012,8.800523,8.636538,8.468649,8.304664,8.140678,7.9766936,7.47693,6.9732623,6.473499,5.9737353,5.473972,5.165524,4.853172,4.5447245,4.2362766,3.9239242,3.193801,2.4597735,1.7257458,0.9956226,0.26159495,0.22645533,0.19131571,0.15617609,0.12103647,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.23426414,0.41386664,0.59737355,0.78088045,0.96438736,1.5969005,2.233318,2.8658314,3.5022488,4.138666,3.8575494,3.5764325,3.2992198,3.018103,2.736986,2.2957885,1.8584955,1.4172981,0.97610056,0.5388075,0.42948425,0.3240654,0.21474212,0.10932326,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.027330816,0.031235218,0.031235218,0.03513962,0.039044023,0.039044023,0.042948425,0.046852827,0.046852827,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.042948425,0.03513962,0.027330816,0.019522011,0.011713207,0.10541886,0.19912452,0.28892577,0.38263142,0.47633708,0.57394713,0.6715572,0.76916724,0.8667773,0.96438736,1.1205635,1.2806439,1.4407244,1.6008049,1.7608855,1.7062237,1.6476578,1.5890918,1.5305257,1.475864,1.5070993,1.5383345,1.5734742,1.6047094,1.6359446,1.6554666,1.6710842,1.6906061,1.7062237,1.7257458,2.1200905,2.514435,2.9087796,3.3031244,3.7013733,4.93126,6.1611466,7.3910336,8.62092,9.850807,8.8200445,7.7892823,6.75852,5.7316628,4.7009,4.521298,4.3416953,4.1581883,3.978586,3.7989833,3.2367494,2.6745155,2.1122816,1.5500476,0.9878138,0.78868926,0.59346914,0.39434463,0.19912452,0.0,0.0,0.0,0.0,0.0,0.0,0.62079996,1.2415999,1.8584955,2.4792955,3.1000953,3.2718892,3.4397783,3.611572,3.7794614,3.951255,4.1113358,4.271416,4.4314966,4.591577,4.7516575,5.989353,7.230953,8.468649,9.710248,10.951848,9.589212,8.23048,6.871748,5.5091114,4.1503797,3.330455,2.5105307,1.6906061,0.8706817,0.05075723,0.07027924,0.08980125,0.10932326,0.12884527,0.14836729,0.19131571,0.23035973,0.26940376,0.30844778,0.3513962,0.3709182,0.39044023,0.40996224,0.42948425,0.44900626,0.3709182,0.28892577,0.21083772,0.12884527,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.046852827,0.093705654,0.14055848,0.19131571,0.23816854,0.21864653,0.20302892,0.1835069,0.1678893,0.14836729,0.14836729,0.14836729,0.14836729,0.14836729,0.14836729,0.28111696,0.41386664,0.5466163,0.679366,0.81211567,0.6481308,0.48805028,0.3240654,0.1639849,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.08199245,0.06637484,0.046852827,0.031235218,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.031235218,0.05075723,0.07418364,0.093705654,0.113227665,0.44119745,0.77307165,1.1010414,1.4329157,1.7608855,1.7530766,1.7491722,1.7413634,1.7335546,1.7257458,1.620327,1.5149081,1.4094892,1.3040704,1.1986516,1.6242313,2.0498111,2.475391,2.900971,3.3265507,3.076669,2.8306916,2.5808098,2.3348327,2.0888553,1.9834363,1.8819219,1.7804074,1.678893,1.5734742,1.6242313,1.6749885,1.7257458,1.7765031,1.8233559,4.2479897,6.6687193,9.093353,11.514082,13.938716,12.11536,10.292005,8.468649,6.649197,4.825841,4.1894236,3.5569105,2.920493,2.2840753,1.6515622,1.6164225,1.5812829,1.5461433,1.5110037,1.475864,1.2533131,1.0346665,0.8160201,0.59346914,0.37482262,0.31625658,0.26159495,0.20302892,0.14446288,0.08589685,0.093705654,0.10151446,0.10932326,0.11713207,0.12494087,0.19912452,0.26940376,0.3435874,0.41386664,0.48805028,0.6676528,0.8472553,1.0268579,1.2064602,1.3860629,1.3626363,1.33921,1.3118792,1.2884527,1.261122,1.1869383,1.1127546,1.038571,0.96438736,0.8862993,0.7106012,0.5309987,0.3553006,0.1756981,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.015617609,0.015617609,0.019522011,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.09761006,0.13274968,0.1678893,0.20302892,0.23816854,0.27721256,0.31625658,0.359205,0.39824903,0.43729305,0.42948425,0.42167544,0.41386664,0.40605783,0.39824903,0.42167544,0.44510186,0.46852827,0.48805028,0.5114767,0.5388075,0.5622339,0.58566034,0.61299115,0.63641757,0.6442264,0.6520352,0.659844,0.6676528,0.6754616,0.57394713,0.46852827,0.3670138,0.26549935,0.1639849,0.13274968,0.10151446,0.07418364,0.042948425,0.011713207,0.031235218,0.05075723,0.07418364,0.093705654,0.113227665,0.12103647,0.13274968,0.14055848,0.15227169,0.1639849,0.14055848,0.11713207,0.093705654,0.07418364,0.05075723,0.078088045,0.10932326,0.14055848,0.1717937,0.19912452,0.28892577,0.37872702,0.46852827,0.5583295,0.6481308,0.8433509,1.0346665,1.2259823,1.4212024,1.6125181,1.6008049,1.5929961,1.5812829,1.5734742,1.5617609,1.3821584,1.2025559,1.0229534,0.8433509,0.6637484,0.6949836,0.7262188,0.76135844,0.79259366,0.8238289,1.639849,2.455869,3.2718892,4.084005,4.900025,4.8375545,4.775084,4.7126136,4.650143,4.5876727,4.466636,4.3455997,4.2284675,4.1074314,3.9863946,3.8263142,3.6623292,3.4983444,3.338264,3.174279,2.97125,2.7643168,2.5612879,2.3543546,2.1513257,1.7647898,1.3782539,0.9956226,0.60908675,0.22645533,0.19522011,0.1639849,0.13665408,0.10541886,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.27330816,0.42557985,0.57394713,0.7262188,0.8745861,1.4485333,2.0263848,2.6003318,3.174279,3.7482262,5.087436,6.426646,7.7619514,9.101162,10.436467,9.351044,8.261715,7.1762915,6.086963,5.001539,4.689187,4.376835,4.0605783,3.7482262,3.435874,2.9751544,2.514435,2.0498111,1.5890918,1.1244678,0.9019169,0.6754616,0.44900626,0.22645533,0.0,0.0,0.0,0.0,0.0,0.0,0.77307165,1.5500476,2.3231194,3.1000953,3.873167,4.087909,4.298747,4.513489,4.7243266,4.939069,5.138193,5.337318,5.5364423,5.735567,5.938596,7.4886436,9.0386915,10.588739,12.138786,13.688834,11.986515,10.2881,8.58578,6.8873653,5.1889505,4.1620927,3.1391394,2.1122816,1.0893283,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.23816854,0.28892577,0.3357786,0.38653582,0.43729305,0.46071947,0.48805028,0.5114767,0.5388075,0.5622339,0.46071947,0.3631094,0.26159495,0.1639849,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.3513962,0.5114767,0.6754616,0.8394465,0.999527,0.80040246,0.60127795,0.39824903,0.19912452,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3357786,0.6754616,1.0112402,1.3509232,1.6867018,1.6125181,1.5383345,1.4641509,1.3860629,1.3118792,1.0619974,0.81211567,0.5622339,0.31235218,0.062470436,0.39824903,0.737932,1.0737107,1.4133936,1.7491722,1.6515622,1.5500476,1.4485333,1.3509232,1.2494087,1.261122,1.2767396,1.2884527,1.3001659,1.3118792,1.0502841,0.78868926,0.5231899,0.26159495,0.0,3.3616903,6.7233806,10.088976,13.450665,16.812357,14.348679,11.888905,9.425227,6.9615493,4.5017757,3.775557,3.049338,2.3231194,1.6008049,0.8745861,0.94876975,1.0268579,1.1010414,1.175225,1.2494087,1.0502841,0.8511597,0.6481308,0.44900626,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.48805028,0.47633708,0.46071947,0.44900626,0.43729305,0.37482262,0.31235218,0.24988174,0.18741131,0.12494087,0.14836729,0.1756981,0.19912452,0.22645533,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.10151446,0.13665408,0.1756981,0.21083772,0.24988174,0.30063897,0.3513962,0.39824903,0.44900626,0.4997635,0.48805028,0.47633708,0.46071947,0.44900626,0.43729305,0.46071947,0.48805028,0.5114767,0.5388075,0.5622339,0.60127795,0.63641757,0.6754616,0.7106012,0.74964523,0.76135844,0.77307165,0.78868926,0.80040246,0.81211567,0.6871748,0.5622339,0.43729305,0.31235218,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.10151446,0.13665408,0.1756981,0.21083772,0.24988174,0.3631094,0.47633708,0.58566034,0.698888,0.81211567,0.999527,1.1869383,1.3743496,1.5617609,1.7491722,1.7765031,1.7999294,1.8233559,1.8506867,1.8741131,1.5500476,1.2259823,0.9019169,0.57394713,0.24988174,0.31235218,0.37482262,0.43729305,0.4997635,0.5622339,1.4485333,2.338737,3.2250361,4.1113358,5.001539,4.0761957,3.1508527,2.2255092,1.3001659,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.1756981,0.3513962,0.5231899,0.698888,0.8745861,0.77307165,0.6754616,0.57394713,0.47633708,0.37482262,0.3357786,0.30063897,0.26159495,0.22645533,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.031235218,0.046852827,0.06637484,0.08199245,0.10151446,0.21864653,0.339683,0.46071947,0.58175594,0.698888,1.1596074,1.620327,2.0810463,2.541766,2.998581,4.068387,5.138193,6.211904,7.28171,8.351517,7.480835,6.610153,5.7394714,4.8687897,3.998108,3.7482262,3.4983444,3.2484627,2.998581,2.7486992,2.3816853,2.0107672,1.639849,1.2689307,0.9019169,0.71841,0.5388075,0.359205,0.1796025,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.62860876,1.2494087,1.8663043,2.4831998,3.1000953,3.2718892,3.4397783,3.611572,3.7794614,3.951255,4.1113358,4.271416,4.4314966,4.591577,4.7516575,5.989353,7.230953,8.468649,9.710248,10.951848,9.600925,8.253906,6.9068875,5.559869,4.21285,3.5373883,2.8619268,2.1864653,1.5110037,0.8394465,0.80430686,0.77307165,0.7418364,0.7066968,0.6754616,0.71841,0.76135844,0.80430686,0.8433509,0.8862993,0.8316377,0.77307165,0.7145056,0.6559396,0.60127795,0.48805028,0.37872702,0.26940376,0.16008049,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.14836729,0.14836729,0.14836729,0.14836729,0.14836729,0.28111696,0.40996224,0.5388075,0.6715572,0.80040246,0.6481308,0.4958591,0.3435874,0.19131571,0.039044023,0.1835069,0.3318742,0.48024148,0.62860876,0.77307165,0.62079996,0.46462387,0.30844778,0.15617609,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.1796025,0.16008049,0.14055848,0.12103647,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.27721256,0.5544251,0.8316377,1.1088502,1.3860629,1.4133936,1.4407244,1.4680552,1.4992905,1.5266213,1.3314011,1.1400855,0.94876975,0.75354964,0.5622339,0.8160201,1.0737107,1.3274968,1.5812829,1.8389735,1.7101282,1.5812829,1.456342,1.3274968,1.1986516,1.1713207,1.1400855,1.1088502,1.0815194,1.0502841,0.8550641,0.659844,0.46462387,0.26940376,0.07418364,2.8111696,5.5442514,8.281238,11.014318,13.751305,12.216875,10.686349,9.151918,7.621393,6.086963,5.2318993,4.376835,3.521771,2.6667068,1.8116426,1.6632754,1.5110037,1.3626363,1.2142692,1.0619974,0.8902037,0.71841,0.5466163,0.3709182,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.24597734,0.28892577,0.3357786,0.37872702,0.42557985,0.40996224,0.39434463,0.37872702,0.3631094,0.3513962,0.30063897,0.24988174,0.19912452,0.14836729,0.10151446,0.12103647,0.14055848,0.16008049,0.1796025,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.10932326,0.14446288,0.1796025,0.21474212,0.24988174,0.29283017,0.3357786,0.37872702,0.42167544,0.46071947,0.45681506,0.45291066,0.44900626,0.44119745,0.43729305,0.46852827,0.5036679,0.5349031,0.5661383,0.60127795,0.62860876,0.659844,0.6910792,0.71841,0.74964523,0.78088045,0.8160201,0.8472553,0.8784905,0.9136301,0.8394465,0.76135844,0.6871748,0.61299115,0.5388075,0.48414588,0.43338865,0.37872702,0.3279698,0.27330816,0.29673457,0.31625658,0.3357786,0.3553006,0.37482262,0.38263142,0.39044023,0.39824903,0.40605783,0.41386664,0.44119745,0.46852827,0.4958591,0.5231899,0.5505207,0.60518235,0.659844,0.7145056,0.76916724,0.8238289,1.1869383,1.5500476,1.9131571,2.2762666,2.639376,2.455869,2.2723622,2.0888553,1.9092526,1.7257458,1.7218413,1.7218413,1.717937,1.7140326,1.7140326,1.4485333,1.1869383,0.92534333,0.6637484,0.39824903,0.42948425,0.46071947,0.48805028,0.5192855,0.5505207,1.2415999,1.9365835,2.6276627,3.3187418,4.0137253,3.2992198,2.5886188,1.8741131,1.1635119,0.44900626,0.3631094,0.27330816,0.18741131,0.10151446,0.011713207,0.14836729,0.28892577,0.42557985,0.5622339,0.698888,0.62079996,0.5388075,0.46071947,0.37872702,0.30063897,0.26940376,0.23816854,0.21083772,0.1796025,0.14836729,0.13665408,0.12494087,0.113227665,0.10151446,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.015617609,0.015617609,0.019522011,0.023426414,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.03513962,0.046852827,0.05466163,0.06637484,0.07418364,0.1639849,0.25378615,0.3435874,0.43338865,0.5231899,0.8706817,1.2142692,1.5617609,1.9053483,2.2489357,3.0532427,3.853645,4.657952,5.4583545,6.262661,5.610626,4.958591,4.3065557,3.6506162,2.998581,2.8111696,2.6237583,2.436347,2.2489357,2.0615244,1.7843118,1.5070993,1.2298868,0.95267415,0.6754616,0.5388075,0.40605783,0.26940376,0.13665408,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.48414588,0.94486535,1.4055848,1.8663043,2.3231194,2.4519646,2.5808098,2.7057507,2.8345962,2.9634414,3.0805733,3.2016098,3.3226464,3.4436827,3.5608149,4.493967,5.423215,6.3524623,7.28171,8.210958,7.2192397,6.223617,5.2279944,4.2323723,3.2367494,2.912684,2.5886188,2.260649,1.9365835,1.6125181,1.5227169,1.4329157,1.3431144,1.2533131,1.1635119,1.1986516,1.2337911,1.2689307,1.3040704,1.33921,1.1986516,1.0580931,0.91753453,0.77697605,0.63641757,0.5192855,0.39824903,0.27721256,0.15617609,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.113227665,0.113227665,0.113227665,0.113227665,0.113227665,0.21083772,0.30844778,0.40605783,0.5036679,0.60127795,0.4958591,0.39044023,0.28502136,0.1796025,0.07418364,0.359205,0.64032197,0.92143893,1.2064602,1.4875772,1.1908426,0.8941081,0.59346914,0.29673457,0.0,0.05466163,0.10932326,0.1639849,0.21864653,0.27330816,0.23426414,0.19522011,0.15617609,0.113227665,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21864653,0.43338865,0.6520352,0.8706817,1.0893283,1.2181735,1.3470187,1.475864,1.6086137,1.737459,1.6008049,1.4680552,1.3314011,1.1986516,1.0619974,1.2337911,1.4055848,1.5812829,1.7530766,1.9248703,1.7686942,1.6164225,1.4602464,1.3040704,1.1517987,1.077615,1.0034313,0.93315214,0.8589685,0.78868926,0.659844,0.5309987,0.40605783,0.27721256,0.14836729,2.2567444,4.365122,6.473499,8.581876,10.686349,10.085071,9.483793,8.878611,8.277332,7.676055,6.688241,5.704332,4.7204223,3.736513,2.7486992,2.3738766,1.999054,1.6242313,1.2494087,0.8745861,0.7301232,0.58566034,0.44119745,0.29673457,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,0.39044023,0.37872702,0.3709182,0.359205,0.3513962,0.3318742,0.31625658,0.29673457,0.28111696,0.26159495,0.22645533,0.18741131,0.14836729,0.113227665,0.07418364,0.08980125,0.10541886,0.12103647,0.13665408,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.12103647,0.15227169,0.1835069,0.21864653,0.24988174,0.28502136,0.32016098,0.3553006,0.39044023,0.42557985,0.42557985,0.42948425,0.43338865,0.43338865,0.43729305,0.47633708,0.5192855,0.5583295,0.59737355,0.63641757,0.659844,0.6832704,0.7066968,0.7262188,0.74964523,0.80430686,0.8550641,0.9058213,0.96048295,1.0112402,0.9878138,0.96438736,0.93705654,0.9136301,0.8862993,0.8199245,0.75354964,0.6832704,0.61689556,0.5505207,0.57785153,0.60518235,0.63251317,0.659844,0.6871748,0.679366,0.6676528,0.6559396,0.6481308,0.63641757,0.71841,0.79649806,0.8784905,0.95657855,1.038571,1.1088502,1.183034,1.2533131,1.3274968,1.4016805,2.0107672,2.6237583,3.2367494,3.8497405,4.462732,3.9083066,3.357786,2.803361,2.25284,1.698415,1.6710842,1.639849,1.6086137,1.5812829,1.5500476,1.3509232,1.1517987,0.94876975,0.74964523,0.5505207,0.5466163,0.5466163,0.5427119,0.5388075,0.5388075,1.0346665,1.53443,2.0302892,2.5261483,3.0259118,2.5261483,2.0263848,1.5266213,1.0268579,0.5231899,0.42557985,0.3240654,0.22645533,0.12494087,0.023426414,0.12494087,0.22645533,0.3240654,0.42557985,0.5231899,0.46462387,0.40605783,0.3435874,0.28502136,0.22645533,0.20302892,0.1796025,0.15617609,0.13665408,0.113227665,0.113227665,0.113227665,0.113227665,0.113227665,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.031235218,0.03513962,0.039044023,0.046852827,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.039044023,0.042948425,0.046852827,0.046852827,0.05075723,0.10932326,0.1717937,0.23035973,0.28892577,0.3513962,0.58175594,0.80821127,1.038571,1.2689307,1.4992905,2.0341935,2.5690966,3.1039999,3.638903,4.173806,3.7404175,3.3031244,2.8697357,2.436347,1.999054,1.8741131,1.7491722,1.6242313,1.4992905,1.3743496,1.1908426,1.0034313,0.8199245,0.63641757,0.44900626,0.359205,0.26940376,0.1796025,0.08980125,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.339683,0.6442264,0.94486535,1.2494087,1.5500476,1.6359446,1.7218413,1.8038338,1.8897307,1.9756275,2.0537157,2.135708,2.2137961,2.2957885,2.3738766,2.9946766,3.6154766,4.2362766,4.853172,5.473972,4.83365,4.1894236,3.5491016,2.9048753,2.260649,2.2879796,2.3114061,2.338737,2.3621633,2.3855898,2.241127,2.0927596,1.9443923,1.796025,1.6515622,1.678893,1.7062237,1.7335546,1.7608855,1.7882162,1.5656652,1.3431144,1.1205635,0.8980125,0.6754616,0.5466163,0.41386664,0.28502136,0.15617609,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.14055848,0.20693332,0.26940376,0.3357786,0.39824903,0.3435874,0.28502136,0.22645533,0.1717937,0.113227665,0.5309987,0.94876975,1.3665408,1.7843118,2.1981785,1.7608855,1.319688,0.8784905,0.44119745,0.0,0.07027924,0.14055848,0.21083772,0.28111696,0.3513962,0.28892577,0.23035973,0.1717937,0.10932326,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15617609,0.31625658,0.47243267,0.62860876,0.78868926,1.0190489,1.2533131,1.4836729,1.717937,1.9482968,1.8741131,1.796025,1.717937,1.639849,1.5617609,1.6515622,1.7413634,1.8311646,1.9209659,2.0107672,1.8311646,1.6476578,1.4641509,1.2806439,1.1010414,0.98390937,0.8706817,0.75354964,0.64032197,0.5231899,0.46462387,0.40605783,0.3435874,0.28502136,0.22645533,1.7062237,3.1859922,4.6657605,6.1455293,7.6252975,7.9532676,8.281238,8.609207,8.933272,9.261242,8.148487,7.0318284,5.919074,4.802415,3.6857557,3.0883822,2.4871042,1.8858263,1.2884527,0.6871748,0.5700427,0.45291066,0.3357786,0.21864653,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.12103647,0.23816854,0.359205,0.48024148,0.60127795,0.5349031,0.46852827,0.40605783,0.339683,0.27330816,0.25378615,0.23426414,0.21474212,0.19522011,0.1756981,0.14836729,0.12494087,0.10151446,0.07418364,0.05075723,0.058566034,0.07027924,0.078088045,0.08980125,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.12884527,0.16008049,0.19131571,0.21864653,0.24988174,0.27721256,0.30454338,0.3318742,0.359205,0.38653582,0.39824903,0.40605783,0.41777104,0.42557985,0.43729305,0.48414588,0.5309987,0.58175594,0.62860876,0.6754616,0.6910792,0.7066968,0.71841,0.7340276,0.74964523,0.8238289,0.8941081,0.96829176,1.038571,1.1127546,1.1361811,1.1635119,1.1869383,1.2142692,1.2376955,1.1557031,1.0737107,0.9917182,0.9058213,0.8238289,0.8589685,0.8941081,0.92924774,0.96438736,0.999527,0.97219616,0.94486535,0.91753453,0.8902037,0.8628729,0.9956226,1.1283722,1.261122,1.3938715,1.5266213,1.6164225,1.7062237,1.796025,1.8858263,1.9756275,2.8385005,3.7013733,4.564246,5.423215,6.2860875,5.364649,4.4432096,3.521771,2.5964274,1.6749885,1.6164225,1.5617609,1.5031948,1.4446288,1.3860629,1.2494087,1.1127546,0.97610056,0.8394465,0.698888,0.6637484,0.62860876,0.59346914,0.5583295,0.5231899,0.8277333,1.1283722,1.4329157,1.7335546,2.0380979,1.7491722,1.4641509,1.175225,0.8862993,0.60127795,0.48805028,0.37482262,0.26159495,0.14836729,0.039044023,0.10151446,0.1639849,0.22645533,0.28892577,0.3513962,0.30844778,0.26940376,0.23035973,0.19131571,0.14836729,0.13665408,0.12103647,0.10541886,0.08980125,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.13665408,0.10932326,0.08199245,0.05466163,0.027330816,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.046852827,0.05075723,0.058566034,0.06637484,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.046852827,0.039044023,0.03513962,0.031235218,0.023426414,0.05466163,0.08589685,0.113227665,0.14446288,0.1756981,0.28892577,0.40605783,0.5192855,0.63641757,0.74964523,1.0190489,1.2845483,1.5539521,1.8194515,2.0888553,1.8702087,1.6515622,1.43682,1.2181735,0.999527,0.93705654,0.8745861,0.81211567,0.74964523,0.6871748,0.59346914,0.5036679,0.40996224,0.31625658,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.19522011,0.339683,0.48414588,0.62860876,0.77307165,0.8160201,0.8589685,0.9019169,0.94486535,0.9878138,1.0268579,1.0659018,1.1088502,1.1478943,1.1869383,1.4992905,1.8077383,2.1161861,2.4285383,2.736986,2.4480603,2.1591344,1.8663043,1.5773785,1.2884527,1.6632754,2.0380979,2.4129205,2.787743,3.1625657,2.9556324,2.7526035,2.5456703,2.3426414,2.135708,2.1591344,2.1786566,2.1981785,2.2177005,2.2372224,1.9326792,1.6281357,1.3235924,1.0190489,0.7106012,0.57394713,0.43338865,0.29283017,0.15227169,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.07027924,0.10151446,0.13665408,0.1678893,0.19912452,0.19131571,0.1796025,0.1717937,0.16008049,0.14836729,0.7027924,1.2533131,1.8077383,2.358259,2.912684,2.330928,1.7491722,1.1635119,0.58175594,0.0,0.08589685,0.1717937,0.25378615,0.339683,0.42557985,0.3435874,0.26549935,0.1835069,0.10541886,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09761006,0.19522011,0.29283017,0.39044023,0.48805028,0.8238289,1.1557031,1.4914817,1.8272603,2.1630387,2.1435168,2.1239948,2.1005683,2.0810463,2.0615244,2.069333,2.077142,2.084951,2.0927596,2.1005683,1.8897307,1.678893,1.4680552,1.261122,1.0502841,0.8941081,0.7340276,0.57785153,0.42167544,0.26159495,0.26940376,0.27721256,0.28502136,0.29283017,0.30063897,1.1517987,2.0068626,2.8580225,3.7091823,4.564246,5.8214636,7.0786815,8.335898,9.593117,10.850334,9.60483,8.359325,7.113821,5.8683167,4.6267166,3.7989833,2.9751544,2.1513257,1.3235924,0.4997635,0.40996224,0.32016098,0.23035973,0.14055848,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.16008049,0.32016098,0.48024148,0.64032197,0.80040246,0.679366,0.5583295,0.44119745,0.32016098,0.19912452,0.1756981,0.15617609,0.13274968,0.10932326,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.031235218,0.03513962,0.039044023,0.046852827,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.14055848,0.1678893,0.19522011,0.22255093,0.24988174,0.26940376,0.28892577,0.30844778,0.3318742,0.3513962,0.3670138,0.38653582,0.40215343,0.42167544,0.43729305,0.49195468,0.5466163,0.60127795,0.6559396,0.7106012,0.71841,0.7262188,0.7340276,0.7418364,0.74964523,0.8433509,0.93315214,1.0268579,1.1205635,1.2142692,1.2884527,1.3626363,1.43682,1.5110037,1.5890918,1.4914817,1.3938715,1.2962615,1.1986516,1.1010414,1.1439898,1.1869383,1.2259823,1.2689307,1.3118792,1.2689307,1.2220778,1.1791295,1.1322767,1.0893283,1.2728351,1.456342,1.6437533,1.8272603,2.0107672,2.1200905,2.2294137,2.3348327,2.4441557,2.5495746,3.6623292,4.775084,5.8878384,7.000593,8.113348,6.8209906,5.5286336,4.2362766,2.9439192,1.6515622,1.5656652,1.4797685,1.3938715,1.3118792,1.2259823,1.1517987,1.0737107,0.999527,0.92534333,0.8511597,0.78088045,0.7145056,0.6481308,0.58175594,0.5114767,0.62079996,0.7262188,0.8355421,0.94096094,1.0502841,0.97610056,0.9019169,0.8238289,0.74964523,0.6754616,0.5505207,0.42557985,0.30063897,0.1756981,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.1756981,0.15617609,0.13665408,0.113227665,0.093705654,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.12884527,0.09761006,0.06637484,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.058566034,0.07027924,0.078088045,0.08980125,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,1.038571,1.7608855,2.4871042,3.213323,3.9356375,3.6740425,3.4124475,3.1508527,2.8892577,2.6237583,2.639376,2.6510892,2.6628022,2.6745155,2.6862288,2.2996929,1.9131571,1.5266213,1.1361811,0.74964523,0.60127795,0.44900626,0.30063897,0.14836729,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.8745861,1.5617609,2.2489357,2.9361105,3.6232853,2.900971,2.174752,1.4485333,0.7262188,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.62470436,1.0619974,1.4992905,1.9365835,2.3738766,2.4129205,2.4480603,2.4871042,2.5261483,2.5612879,2.4871042,2.4129205,2.338737,2.260649,2.1864653,1.9482968,1.7140326,1.475864,1.2376955,0.999527,0.80040246,0.60127795,0.39824903,0.19912452,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.60127795,0.8238289,1.0502841,1.2767396,1.4992905,3.6857557,5.8761253,8.062591,10.249056,12.439425,11.061172,9.686822,8.312472,6.9381227,5.563773,4.513489,3.4632049,2.4129205,1.3626363,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.0,0.0,0.0,0.0,0.0,0.19912452,0.39824903,0.60127795,0.80040246,0.999527,0.8238289,0.6481308,0.47633708,0.30063897,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.1756981,0.19912452,0.22645533,0.24988174,0.26159495,0.27330816,0.28892577,0.30063897,0.31235218,0.3357786,0.3631094,0.38653582,0.41386664,0.43729305,0.4997635,0.5622339,0.62470436,0.6871748,0.74964523,0.74964523,0.74964523,0.74964523,0.74964523,0.74964523,0.8628729,0.97610056,1.0893283,1.1986516,1.3118792,1.43682,1.5617609,1.6867018,1.8116426,1.9365835,1.8233559,1.7140326,1.6008049,1.4875772,1.3743496,1.4251068,1.475864,1.5266213,1.5734742,1.6242313,1.5617609,1.4992905,1.43682,1.3743496,1.3118792,1.5500476,1.7882162,2.0263848,2.260649,2.4988174,2.6237583,2.7486992,2.87364,2.998581,3.1235218,4.4861584,5.8487945,7.211431,8.574067,9.936704,8.273428,6.6140575,4.950782,3.2875066,1.6242313,1.5110037,1.4016805,1.2884527,1.175225,1.0619974,1.0502841,1.038571,1.0268579,1.0112402,0.999527,0.9019169,0.80040246,0.698888,0.60127795,0.4997635,0.41386664,0.3240654,0.23816854,0.14836729,0.062470436,0.19912452,0.3357786,0.47633708,0.61299115,0.74964523,0.61299115,0.47633708,0.3357786,0.19912452,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22255093,0.44510186,0.6676528,0.8902037,1.1127546,0.93315214,0.75745404,0.58175594,0.40215343,0.22645533,0.27330816,0.32016098,0.3670138,0.41386664,0.46071947,0.3709182,0.28111696,0.19131571,0.10151446,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.8316377,1.4094892,1.9912452,2.5690966,3.1508527,2.9751544,2.7994564,2.6237583,2.4480603,2.2762666,2.280171,2.2840753,2.2918842,2.2957885,2.2996929,1.9639144,1.6281357,1.2962615,0.96048295,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.78088045,1.4133936,2.0459068,2.67842,3.310933,2.7018464,2.0888553,1.475864,0.8628729,0.24988174,0.359205,0.46462387,0.57394713,0.679366,0.78868926,0.6442264,0.4958591,0.3513962,0.20693332,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.37482262,0.43338865,0.4958591,0.5544251,0.61689556,0.6754616,0.5661383,0.45681506,0.3435874,0.23426414,0.12494087,0.14836729,0.1756981,0.19912452,0.22645533,0.24988174,0.59346914,0.94096094,1.2845483,1.6281357,1.9756275,1.9912452,2.0068626,2.018576,2.0341935,2.0498111,2.0810463,2.1083772,2.1396124,2.1708477,2.1981785,2.1786566,2.15523,2.1318035,2.1083772,2.0888553,1.8038338,1.5188124,1.2337911,0.94876975,0.6637484,0.6754616,0.6871748,0.698888,0.7106012,0.7262188,0.8784905,1.0307622,1.183034,1.3353056,1.4875772,3.377308,5.267039,7.1567693,9.0465,10.936231,9.706344,8.476458,7.2465706,6.016684,4.786797,3.900498,3.018103,2.1318035,1.2494087,0.3631094,0.31625658,0.27330816,0.22645533,0.1835069,0.13665408,0.10932326,0.08199245,0.05466163,0.027330816,0.0,0.16008049,0.32016098,0.48024148,0.64032197,0.80040246,0.659844,0.5192855,0.37872702,0.23816854,0.10151446,0.093705654,0.08980125,0.08589685,0.078088045,0.07418364,0.08980125,0.10541886,0.12103647,0.13665408,0.14836729,0.13274968,0.113227665,0.09761006,0.078088045,0.062470436,0.07418364,0.08199245,0.093705654,0.10151446,0.113227665,0.10151446,0.093705654,0.08199245,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.12103647,0.14446288,0.1678893,0.19131571,0.21083772,0.22645533,0.23816854,0.24988174,0.26159495,0.27330816,0.30454338,0.3357786,0.3631094,0.39434463,0.42557985,0.48414588,0.5466163,0.60518235,0.6637484,0.7262188,0.71841,0.7106012,0.7027924,0.6949836,0.6871748,0.78868926,0.8941081,0.9956226,1.097137,1.1986516,1.3938715,1.5890918,1.7843118,1.979532,2.174752,1.9834363,1.7882162,1.5969005,1.4055848,1.2142692,1.3899672,1.5656652,1.7452679,1.9209659,2.1005683,2.084951,2.069333,2.0537157,2.0380979,2.0263848,2.0654287,2.1044729,2.1435168,2.1864653,2.2255092,2.5612879,2.893162,3.2289407,3.5647192,3.900498,4.806319,5.716045,6.621866,7.531592,8.437413,7.0903945,5.743376,4.396357,3.049338,1.698415,1.5812829,1.4641509,1.3470187,1.2298868,1.1127546,1.1361811,1.1557031,1.1791295,1.2025559,1.2259823,1.1088502,0.9956226,0.8784905,0.76526284,0.6481308,0.58566034,0.5192855,0.45681506,0.39044023,0.3240654,0.42557985,0.5231899,0.62470436,0.7262188,0.8238289,0.7301232,0.63641757,0.5388075,0.44510186,0.3513962,0.3631094,0.37482262,0.38653582,0.39824903,0.41386664,0.3318742,0.24597734,0.1639849,0.08199245,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.039044023,0.06637484,0.093705654,0.12103647,0.14836729,0.12884527,0.10541886,0.08199245,0.058566034,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.093705654,0.10932326,0.12884527,0.14446288,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.44510186,0.8902037,1.3353056,1.7804074,2.2255092,1.8702087,1.5149081,1.1596074,0.80430686,0.44900626,0.5466163,0.64032197,0.7340276,0.8316377,0.92534333,0.74574083,0.5661383,0.38653582,0.20693332,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.62079996,1.0580931,1.4914817,1.9287747,2.3621633,2.2762666,2.1864653,2.1005683,2.0107672,1.9248703,1.9209659,1.9209659,1.9170616,1.9131571,1.9131571,1.6281357,1.3470187,1.0659018,0.78088045,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.6910792,1.2689307,1.8467822,2.4207294,2.998581,2.4988174,1.999054,1.4992905,0.999527,0.4997635,0.61689556,0.7301232,0.8433509,0.96048295,1.0737107,0.8862993,0.6949836,0.5036679,0.31625658,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,0.74964523,0.8706817,0.9917182,1.1088502,1.2298868,1.3509232,1.1283722,0.9097257,0.6910792,0.46852827,0.24988174,0.26159495,0.27330816,0.28892577,0.30063897,0.31235218,0.5661383,0.8160201,1.0698062,1.3235924,1.5734742,1.5656652,1.5617609,1.5539521,1.5461433,1.5383345,1.6710842,1.8077383,1.9443923,2.077142,2.2137961,2.4051118,2.5964274,2.7916477,2.9829633,3.174279,2.803361,2.436347,2.0654287,1.6945106,1.3235924,1.2767396,1.2259823,1.175225,1.1244678,1.0737107,1.1557031,1.2337911,1.3157835,1.3938715,1.475864,3.06886,4.661856,6.250948,7.843944,9.43694,8.351517,7.266093,6.180669,5.099149,4.0137253,3.2914112,2.5730011,1.8506867,1.1322767,0.41386664,0.38653582,0.359205,0.3318742,0.30063897,0.27330816,0.21864653,0.1639849,0.10932326,0.05466163,0.0,0.12103647,0.23816854,0.359205,0.48024148,0.60127795,0.4958591,0.39044023,0.28502136,0.1796025,0.07418364,0.08980125,0.10541886,0.12103647,0.13665408,0.14836729,0.1796025,0.21083772,0.23816854,0.26940376,0.30063897,0.26549935,0.23035973,0.19522011,0.16008049,0.12494087,0.14446288,0.1639849,0.1835069,0.20693332,0.22645533,0.20693332,0.1835069,0.1639849,0.14446288,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.093705654,0.113227665,0.13665408,0.15617609,0.1756981,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.27330816,0.30844778,0.3435874,0.37872702,0.41386664,0.46852827,0.5270943,0.58566034,0.6442264,0.698888,0.6832704,0.6715572,0.6559396,0.64032197,0.62470436,0.71841,0.80821127,0.9019169,0.9956226,1.0893283,1.3509232,1.6164225,1.8819219,2.1474214,2.4129205,2.1396124,1.8663043,1.5969005,1.3235924,1.0502841,1.3548276,1.6593709,1.9639144,2.2684577,2.5769055,2.6081407,2.639376,2.6706111,2.7057507,2.736986,2.5808098,2.4207294,2.2645533,2.1083772,1.9482968,2.494913,3.0415294,3.5842414,4.1308575,4.6735697,5.12648,5.579391,6.0323014,6.4852123,6.9381227,5.903456,4.872694,3.8380275,2.8072653,1.7765031,1.6515622,1.5305257,1.4055848,1.2845483,1.1635119,1.2181735,1.2767396,1.3353056,1.3938715,1.4485333,1.319688,1.1908426,1.0580931,0.92924774,0.80040246,0.75745404,0.7145056,0.6715572,0.62860876,0.58566034,0.6481308,0.7106012,0.77307165,0.8394465,0.9019169,0.8472553,0.79649806,0.7418364,0.6910792,0.63641757,0.6754616,0.7106012,0.74964523,0.78868926,0.8238289,0.659844,0.4958591,0.3318742,0.1639849,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.042948425,0.058566034,0.078088045,0.093705654,0.113227665,0.10541886,0.09761006,0.08980125,0.08199245,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.10932326,0.13274968,0.15617609,0.1756981,0.19912452,0.1756981,0.14836729,0.12494087,0.10151446,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6676528,1.3353056,2.0029583,2.6706111,3.338264,2.803361,2.2723622,1.7413634,1.2064602,0.6754616,0.8160201,0.96048295,1.1010414,1.2455044,1.3860629,1.116659,0.8472553,0.57785153,0.30844778,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.41386664,0.7066968,0.9956226,1.2845483,1.5734742,1.5734742,1.5734742,1.5734742,1.5734742,1.5734742,1.5656652,1.5539521,1.5461433,1.53443,1.5266213,1.2962615,1.0659018,0.8355421,0.60518235,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.59737355,1.1205635,1.6437533,2.1669433,2.6862288,2.2996929,1.9131571,1.5266213,1.1361811,0.74964523,0.8706817,0.9956226,1.116659,1.2415999,1.3626363,1.1283722,0.8941081,0.6559396,0.42167544,0.18741131,0.37482262,0.5622339,0.74964523,0.93705654,1.1244678,1.3040704,1.4836729,1.6632754,1.8467822,2.0263848,1.6945106,1.3665408,1.0346665,0.7066968,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.5349031,0.6949836,0.8550641,1.0151446,1.175225,1.1439898,1.116659,1.0854238,1.0541886,1.0268579,1.2650263,1.5031948,1.7452679,1.9834363,2.2255092,2.631567,3.0415294,3.4475873,3.853645,4.263607,3.8067923,3.3538816,2.8970666,2.4441557,1.9873407,1.8741131,1.7608855,1.6515622,1.5383345,1.4251068,1.4329157,1.4407244,1.4485333,1.456342,1.4641509,2.7565079,4.0527697,5.349031,6.6413884,7.9376497,6.996689,6.055728,5.1186714,4.1777105,3.2367494,2.6823244,2.1278992,1.5734742,1.0190489,0.46071947,0.45291066,0.44119745,0.43338865,0.42167544,0.41386664,0.3318742,0.24597734,0.1639849,0.08199245,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,0.3318742,0.26159495,0.19131571,0.12103647,0.05075723,0.08589685,0.12103647,0.15617609,0.19131571,0.22645533,0.26940376,0.31625658,0.359205,0.40605783,0.44900626,0.39824903,0.3435874,0.29283017,0.23816854,0.18741131,0.21864653,0.24597734,0.27721256,0.30844778,0.3357786,0.30844778,0.27721256,0.24597734,0.21864653,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.06637484,0.08589685,0.10151446,0.12103647,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.19912452,0.23816854,0.28111696,0.32016098,0.359205,0.39824903,0.45681506,0.5114767,0.5661383,0.62079996,0.6754616,0.6520352,0.62860876,0.60908675,0.58566034,0.5622339,0.6442264,0.7262188,0.80821127,0.8941081,0.97610056,1.3118792,1.6437533,1.979532,2.3153105,2.6510892,2.2957885,1.9443923,1.5929961,1.2415999,0.8862993,1.319688,1.7530766,2.1864653,2.6159496,3.049338,3.1313305,3.2094188,3.2914112,3.3694992,3.4514916,3.096191,2.7408905,2.3855898,2.0302892,1.6749885,2.4285383,3.1859922,3.9395418,4.6930914,5.4505453,5.446641,5.446641,5.4427366,5.4388323,5.4388323,4.7204223,4.0020123,3.2836022,2.5690966,1.8506867,1.7218413,1.5969005,1.4680552,1.33921,1.2142692,1.3040704,1.397776,1.4914817,1.5812829,1.6749885,1.5305257,1.3860629,1.2415999,1.0932326,0.94876975,0.92924774,0.9097257,0.8902037,0.8706817,0.8511597,0.8745861,0.9019169,0.92534333,0.94876975,0.97610056,0.96438736,0.95657855,0.94486535,0.93315214,0.92534333,0.9878138,1.0502841,1.1127546,1.175225,1.2376955,0.9917182,0.7418364,0.4958591,0.24597734,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.046852827,0.05075723,0.058566034,0.06637484,0.07418364,0.08199245,0.08980125,0.09761006,0.10541886,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.12884527,0.15617609,0.1835069,0.21083772,0.23816854,0.21083772,0.18741131,0.1639849,0.13665408,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.8902037,1.7804074,2.6706111,3.5608149,4.4510183,3.7404175,3.0298162,2.3192148,1.6086137,0.9019169,1.0893283,1.2806439,1.4719596,1.6593709,1.8506867,1.4914817,1.1283722,0.76916724,0.40996224,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.20693332,0.3513962,0.4958591,0.6442264,0.78868926,0.8745861,0.96438736,1.0502841,1.1361811,1.2259823,1.2064602,1.1908426,1.1713207,1.1557031,1.1361811,0.96048295,0.78088045,0.60518235,0.42557985,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.5036679,0.97219616,1.4407244,1.9092526,2.3738766,2.1005683,1.8233559,1.5500476,1.2767396,0.999527,1.1283722,1.261122,1.3899672,1.5188124,1.6515622,1.3704453,1.0893283,0.80821127,0.5309987,0.24988174,0.4997635,0.74964523,0.999527,1.2494087,1.4992905,1.7413634,1.979532,2.2216048,2.4597735,2.7018464,2.260649,1.8194515,1.3782539,0.94096094,0.4997635,0.48805028,0.47633708,0.46071947,0.44900626,0.43729305,0.5036679,0.57394713,0.64032197,0.7066968,0.77307165,0.7223144,0.6715572,0.61689556,0.5661383,0.5114767,0.8589685,1.2025559,1.5461433,1.893635,2.2372224,2.8619268,3.4827268,4.1035266,4.728231,5.349031,4.8102236,4.271416,3.7287042,3.1898966,2.6510892,2.475391,2.2996929,2.1239948,1.9482968,1.7765031,1.7101282,1.6437533,1.5812829,1.5149081,1.4485333,2.4480603,3.4436827,4.4432096,5.4388323,6.4383593,5.6418614,4.8492675,4.0527697,3.2562714,2.463678,2.0732377,1.6827974,1.2923572,0.9019169,0.5114767,0.5192855,0.5270943,0.5349031,0.5427119,0.5505207,0.44119745,0.3318742,0.21864653,0.10932326,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.1639849,0.12884527,0.093705654,0.058566034,0.023426414,0.078088045,0.13665408,0.19131571,0.24597734,0.30063897,0.359205,0.42167544,0.48024148,0.5388075,0.60127795,0.5309987,0.46071947,0.39044023,0.32016098,0.24988174,0.28892577,0.3318742,0.3709182,0.40996224,0.44900626,0.40996224,0.3709182,0.3318742,0.28892577,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.039044023,0.05466163,0.07027924,0.08589685,0.10151446,0.113227665,0.12494087,0.13665408,0.14836729,0.1639849,0.20693332,0.25378615,0.29673457,0.3435874,0.38653582,0.44119745,0.49195468,0.5466163,0.59737355,0.6481308,0.62079996,0.58956474,0.5583295,0.5309987,0.4997635,0.57394713,0.6442264,0.71841,0.78868926,0.8628729,1.2689307,1.6710842,2.077142,2.4831998,2.8892577,2.455869,2.0224805,1.5890918,1.1557031,0.7262188,1.2845483,1.8467822,2.4051118,2.9634414,3.5256753,3.6506162,3.7794614,3.9083066,4.0332475,4.1620927,3.611572,3.057147,2.5066261,1.9522011,1.4016805,2.366068,3.330455,4.2948427,5.2592297,6.223617,5.7668023,5.309987,4.853172,4.396357,3.9356375,3.533484,3.1313305,2.7291772,2.3270237,1.9248703,1.7921207,1.6593709,1.5266213,1.3938715,1.261122,1.3899672,1.5188124,1.6437533,1.7725986,1.901444,1.7413634,1.5812829,1.4212024,1.261122,1.1010414,1.1010414,1.1049459,1.1088502,1.1088502,1.1127546,1.1010414,1.0893283,1.0737107,1.0619974,1.0502841,1.0815194,1.116659,1.1478943,1.1791295,1.2142692,1.3001659,1.3860629,1.475864,1.5617609,1.6515622,1.319688,0.9917182,0.659844,0.3318742,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.046852827,0.046852827,0.042948425,0.039044023,0.039044023,0.058566034,0.08199245,0.10541886,0.12884527,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.14446288,0.1756981,0.21083772,0.24207294,0.27330816,0.24988174,0.22645533,0.19912452,0.1756981,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1127546,2.2255092,3.338264,4.4510183,5.563773,4.6735697,3.78727,2.900971,2.0107672,1.1244678,1.3626363,1.6008049,1.8389735,2.0732377,2.3114061,1.8623998,1.4133936,0.96438736,0.5114767,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1756981,0.3513962,0.5231899,0.698888,0.8745861,0.8511597,0.8238289,0.80040246,0.77307165,0.74964523,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.41386664,0.8238289,1.2376955,1.6515622,2.0615244,1.901444,1.737459,1.5734742,1.4133936,1.2494087,1.3860629,1.5266213,1.6632754,1.7999294,1.9365835,1.6125181,1.2884527,0.96438736,0.63641757,0.31235218,0.62470436,0.93705654,1.2494087,1.5617609,1.8741131,2.174752,2.475391,2.77603,3.076669,3.3734035,2.8267872,2.2762666,1.7257458,1.175225,0.62470436,0.60127795,0.57394713,0.5505207,0.5231899,0.4997635,0.47633708,0.44900626,0.42557985,0.39824903,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.44900626,0.9019169,1.3509232,1.7999294,2.2489357,3.0883822,3.9239242,4.7633705,5.5989127,6.4383593,5.813655,5.1889505,4.564246,3.9356375,3.310933,3.076669,2.8385005,2.6003318,2.3621633,2.1239948,1.9873407,1.8506867,1.7140326,1.5734742,1.43682,2.135708,2.8385005,3.5373883,4.2362766,4.939069,4.2870336,3.638903,2.9868677,2.338737,1.6867018,1.4641509,1.2376955,1.0112402,0.78868926,0.5622339,0.58566034,0.61299115,0.63641757,0.6637484,0.6871748,0.5505207,0.41386664,0.27330816,0.13665408,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.44900626,0.5231899,0.60127795,0.6754616,0.74964523,0.6637484,0.57394713,0.48805028,0.39824903,0.31235218,0.3631094,0.41386664,0.46071947,0.5114767,0.5622339,0.5114767,0.46071947,0.41386664,0.3631094,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.1756981,0.22645533,0.27330816,0.3240654,0.37482262,0.42557985,0.47633708,0.5231899,0.57394713,0.62470436,0.58566034,0.5505207,0.5114767,0.47633708,0.43729305,0.4997635,0.5622339,0.62470436,0.6871748,0.74964523,1.2259823,1.698415,2.174752,2.6510892,3.1235218,2.612045,2.1005683,1.5890918,1.0737107,0.5622339,1.2494087,1.9365835,2.6237583,3.310933,3.998108,4.173806,4.349504,4.5252023,4.7009,4.8765984,4.123049,3.3734035,2.6237583,1.8741131,1.1244678,2.2996929,3.474918,4.650143,5.825368,7.000593,6.086963,5.173333,4.263607,3.349977,2.436347,2.35045,2.260649,2.174752,2.0888553,1.999054,1.8623998,1.7257458,1.5890918,1.4485333,1.3118792,1.475864,1.6359446,1.7999294,1.9639144,2.1239948,1.9482968,1.7765031,1.6008049,1.4251068,1.2494087,1.2767396,1.3001659,1.3235924,1.3509232,1.3743496,1.3235924,1.2767396,1.2259823,1.175225,1.1244678,1.1986516,1.2767396,1.3509232,1.4251068,1.4992905,1.6125181,1.7257458,1.8389735,1.9482968,2.0615244,1.6515622,1.2376955,0.8238289,0.41386664,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.1639849,0.19912452,0.23816854,0.27330816,0.31235218,0.28892577,0.26159495,0.23816854,0.21083772,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.92924774,1.8584955,2.7916477,3.7208953,4.650143,4.2557983,3.8653584,3.4710135,3.0805733,2.6862288,2.5769055,2.463678,2.35045,2.2372224,2.1239948,1.7101282,1.2962615,0.8784905,0.46462387,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14055848,0.28111696,0.42167544,0.5583295,0.698888,0.679366,0.659844,0.64032197,0.62079996,0.60127795,0.5036679,0.40605783,0.30844778,0.21083772,0.113227665,0.09761006,0.08199245,0.06637484,0.05075723,0.039044023,0.031235218,0.027330816,0.023426414,0.015617609,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.08589685,0.1639849,0.23816854,0.31235218,0.38653582,0.31625658,0.24207294,0.1717937,0.09761006,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.3318742,0.659844,0.9917182,1.319688,1.6515622,1.5227169,1.3938715,1.2689307,1.1400855,1.0112402,1.1283722,1.2494087,1.3665408,1.4836729,1.6008049,1.3860629,1.1713207,0.95657855,0.7418364,0.5231899,0.7301232,0.93315214,1.1400855,1.3431144,1.5500476,1.8038338,2.0615244,2.3153105,2.5690966,2.8267872,2.5066261,2.1903696,1.8741131,1.5539521,1.2376955,1.5070993,1.7765031,2.0459068,2.3192148,2.5886188,2.1435168,1.698415,1.2533131,0.80821127,0.3631094,0.48024148,0.59737355,0.7145056,0.8316377,0.94876975,1.1205635,1.2884527,1.4602464,1.6281357,1.7999294,2.4910088,3.1859922,3.8770714,4.5681505,5.263134,4.802415,4.3416953,3.8809757,3.4241607,2.9634414,2.8619268,2.7643168,2.6628022,2.5612879,2.463678,2.2684577,2.0732377,1.8780174,1.6827974,1.4875772,2.1239948,2.7565079,3.3929255,4.029343,4.661856,4.2362766,3.8067923,3.3812122,2.951728,2.5261483,2.1630387,1.7999294,1.43682,1.0737107,0.7106012,0.6832704,0.6559396,0.62860876,0.60127795,0.57394713,0.46071947,0.3435874,0.23035973,0.113227665,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.39434463,0.47243267,0.5544251,0.63251317,0.7106012,0.62079996,0.5309987,0.44119745,0.3513962,0.26159495,0.30063897,0.3357786,0.37482262,0.41386664,0.44900626,0.40996224,0.3709182,0.3318742,0.28892577,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.06637484,0.078088045,0.093705654,0.10932326,0.12494087,0.1678893,0.21083772,0.25378615,0.29673457,0.3357786,0.38263142,0.42557985,0.47243267,0.5192855,0.5622339,0.5427119,0.5231899,0.5036679,0.48414588,0.46071947,0.5231899,0.58566034,0.6481308,0.7106012,0.77307165,1.1557031,1.53443,1.9131571,2.2957885,2.6745155,2.2567444,1.8350691,1.4133936,0.9956226,0.57394713,1.1205635,1.6632754,2.2098918,2.7565079,3.2992198,3.455396,3.611572,3.7638438,3.9200199,4.0761957,3.6506162,3.2289407,2.8072653,2.3855898,1.9639144,2.8385005,3.716991,4.5954814,5.473972,6.348558,5.5989127,4.845363,4.0918136,3.338264,2.5886188,2.4480603,2.3075018,2.1669433,2.0263848,1.8858263,1.7413634,1.5969005,1.4524376,1.3079748,1.1635119,1.2806439,1.397776,1.5149081,1.6320401,1.7491722,1.6008049,1.4485333,1.3001659,1.1517987,0.999527,1.0229534,1.0463798,1.0659018,1.0893283,1.1127546,1.1127546,1.1127546,1.1127546,1.1127546,1.1127546,1.175225,1.2376955,1.3001659,1.3626363,1.4251068,1.5539521,1.678893,1.8077383,1.9365835,2.0615244,1.678893,1.2923572,0.9058213,0.5231899,0.13665408,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.08589685,0.093705654,0.10541886,0.113227665,0.12494087,0.13274968,0.14055848,0.14836729,0.15617609,0.1639849,0.14446288,0.12884527,0.10932326,0.093705654,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.19522011,0.22645533,0.26159495,0.29283017,0.3240654,0.30844778,0.28892577,0.27330816,0.25378615,0.23816854,0.19912452,0.15617609,0.11713207,0.078088045,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.74574083,1.4953861,2.241127,2.9907722,3.736513,3.8419318,3.9434462,4.044961,4.1464753,4.251894,3.78727,3.3265507,2.8619268,2.4012074,1.9365835,1.5578566,1.1791295,0.79649806,0.41777104,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10541886,0.21083772,0.31625658,0.42167544,0.5231899,0.5114767,0.4958591,0.48024148,0.46462387,0.44900626,0.37872702,0.30844778,0.23816854,0.1717937,0.10151446,0.093705654,0.08980125,0.08589685,0.078088045,0.07418364,0.06637484,0.05466163,0.046852827,0.03513962,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.1756981,0.3240654,0.47633708,0.62470436,0.77307165,0.62860876,0.48414588,0.339683,0.19522011,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.24597734,0.4958591,0.7418364,0.9917182,1.2376955,1.1439898,1.0541886,0.96048295,0.8667773,0.77307165,0.8706817,0.96829176,1.0659018,1.1635119,1.261122,1.1557031,1.0541886,0.94876975,0.8433509,0.737932,0.8355421,0.93315214,1.0307622,1.1283722,1.2259823,1.43682,1.6437533,1.8545911,2.0654287,2.2762666,2.1903696,2.1044729,2.018576,1.9365835,1.8506867,2.416825,2.979059,3.5451972,4.1113358,4.6735697,3.8106966,2.9439192,2.0810463,1.2142692,0.3513962,0.659844,0.96829176,1.2806439,1.5890918,1.901444,1.7882162,1.678893,1.5695697,1.4602464,1.3509232,1.8975395,2.4441557,2.9907722,3.541293,4.087909,3.7911747,3.4983444,3.2016098,2.9087796,2.612045,2.6510892,2.6862288,2.7252727,2.7643168,2.7994564,2.5456703,2.2957885,2.0420024,1.7882162,1.5383345,2.1083772,2.67842,3.2484627,3.8185053,4.388548,4.181615,3.978586,3.7716527,3.5686235,3.3616903,2.8619268,2.3621633,1.8623998,1.3626363,0.8628729,0.78088045,0.7027924,0.62079996,0.5427119,0.46071947,0.3709182,0.27721256,0.1835069,0.093705654,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.3357786,0.42167544,0.5036679,0.58956474,0.6754616,0.58175594,0.49195468,0.39824903,0.30454338,0.21083772,0.23816854,0.26159495,0.28892577,0.31235218,0.3357786,0.30844778,0.27721256,0.24597734,0.21864653,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.05466163,0.07418364,0.08980125,0.10932326,0.12494087,0.16008049,0.19522011,0.23035973,0.26549935,0.30063897,0.339683,0.37872702,0.42167544,0.46071947,0.4997635,0.4958591,0.4958591,0.49195468,0.48805028,0.48805028,0.5505207,0.61299115,0.6754616,0.737932,0.80040246,1.0854238,1.3704453,1.6554666,1.9404879,2.2255092,1.8975395,1.5695697,1.2415999,0.9136301,0.58566034,0.9917182,1.3938715,1.796025,2.1981785,2.6003318,2.7330816,2.8697357,3.0063896,3.1391394,3.2757936,3.1781836,3.084478,2.9907722,2.893162,2.7994564,3.3812122,3.959064,4.5408196,5.1186714,5.700427,5.1069584,4.513489,3.9239242,3.330455,2.736986,2.5456703,2.3543546,2.1591344,1.9678187,1.7765031,1.6242313,1.4680552,1.3157835,1.1635119,1.0112402,1.0854238,1.1557031,1.2298868,1.3040704,1.3743496,1.2494087,1.1244678,0.999527,0.8745861,0.74964523,0.76916724,0.78868926,0.80821127,0.8316377,0.8511597,0.9019169,0.94876975,0.999527,1.0502841,1.1010414,1.1517987,1.1986516,1.2494087,1.3001659,1.3509232,1.4914817,1.6359446,1.7765031,1.9209659,2.0615244,1.7062237,1.3470187,0.9917182,0.63251317,0.27330816,0.23816854,0.19912452,0.1639849,0.12494087,0.08589685,0.12103647,0.15227169,0.1835069,0.21864653,0.24988174,0.22645533,0.20693332,0.1835069,0.16008049,0.13665408,0.14055848,0.14055848,0.14446288,0.14836729,0.14836729,0.13665408,0.12103647,0.10541886,0.08980125,0.07418364,0.10151446,0.12494087,0.14836729,0.1756981,0.19912452,0.22645533,0.25378615,0.28111696,0.30844778,0.3357786,0.3279698,0.31625658,0.30844778,0.29673457,0.28892577,0.24597734,0.20302892,0.16008049,0.11713207,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5661383,1.1283722,1.6945106,2.260649,2.8267872,3.4241607,4.0215344,4.618908,5.2162814,5.813655,5.001539,4.1894236,3.3734035,2.5612879,1.7491722,1.4055848,1.0580931,0.7145056,0.3709182,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07027924,0.14055848,0.21083772,0.28111696,0.3513962,0.339683,0.3318742,0.32016098,0.30844778,0.30063897,0.25769055,0.21474212,0.1717937,0.12884527,0.08589685,0.093705654,0.09761006,0.10151446,0.10932326,0.113227665,0.09761006,0.08199245,0.06637484,0.05075723,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.26159495,0.48805028,0.7106012,0.93705654,1.1635119,0.94486535,0.7262188,0.5114767,0.29283017,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.1639849,0.3318742,0.4958591,0.659844,0.8238289,0.76916724,0.7106012,0.6520352,0.59346914,0.5388075,0.61689556,0.6910792,0.76916724,0.8472553,0.92534333,0.92924774,0.93315214,0.94096094,0.94486535,0.94876975,0.94096094,0.92924774,0.92143893,0.9097257,0.9019169,1.0659018,1.2298868,1.3938715,1.5617609,1.7257458,1.8741131,2.018576,2.1669433,2.3153105,2.463678,3.3226464,4.181615,5.040583,5.903456,6.7624245,5.477876,4.193328,2.9087796,1.6242313,0.3357786,0.8394465,1.3431144,1.8467822,2.3465457,2.8502135,2.4597735,2.069333,1.678893,1.2884527,0.9019169,1.3040704,1.7062237,2.1083772,2.5105307,2.912684,2.7838387,2.6510892,2.522244,2.3933985,2.260649,2.436347,2.612045,2.787743,2.9634414,3.1391394,2.8267872,2.5183394,2.2059872,1.8975395,1.5890918,2.0927596,2.5964274,3.1039999,3.6076677,4.1113358,4.1308575,4.1464753,4.165997,4.181615,4.2011366,3.5608149,2.9243972,2.2879796,1.6515622,1.0112402,0.8784905,0.74574083,0.61689556,0.48414588,0.3513962,0.28111696,0.21083772,0.14055848,0.07027924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.27721256,0.3670138,0.45681506,0.5466163,0.63641757,0.5427119,0.44900626,0.3513962,0.25769055,0.1639849,0.1756981,0.18741131,0.19912452,0.21083772,0.22645533,0.20693332,0.1835069,0.1639849,0.14446288,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.046852827,0.06637484,0.08589685,0.10541886,0.12494087,0.15227169,0.1796025,0.20693332,0.23426414,0.26159495,0.29673457,0.3318742,0.3670138,0.40215343,0.43729305,0.45291066,0.46852827,0.48414588,0.4958591,0.5114767,0.57394713,0.63641757,0.698888,0.76135844,0.8238289,1.0151446,1.2064602,1.3938715,1.5851873,1.7765031,1.5383345,1.3040704,1.0698062,0.8355421,0.60127795,0.8589685,1.1205635,1.3782539,1.639849,1.901444,2.0146716,2.1318035,2.2450314,2.358259,2.475391,2.7057507,2.9400148,3.174279,3.4046388,3.638903,3.9200199,4.2011366,4.4861584,4.7672753,5.0483923,4.618908,4.185519,3.7521305,3.3187418,2.8892577,2.6432803,2.397303,2.1513257,1.9092526,1.6632754,1.5031948,1.3431144,1.183034,1.0229534,0.8628729,0.8902037,0.91753453,0.94486535,0.97219616,0.999527,0.9019169,0.80040246,0.698888,0.60127795,0.4997635,0.5192855,0.5349031,0.5544251,0.5700427,0.58566034,0.6871748,0.78868926,0.8862993,0.9878138,1.0893283,1.1244678,1.1635119,1.1986516,1.2376955,1.2767396,1.4329157,1.5890918,1.7491722,1.9053483,2.0615244,1.7335546,1.4016805,1.0737107,0.7418364,0.41386664,0.3513962,0.28892577,0.22645533,0.1639849,0.10151446,0.15617609,0.21083772,0.26549935,0.32016098,0.37482262,0.3240654,0.26940376,0.21864653,0.1639849,0.113227665,0.13665408,0.15617609,0.1796025,0.20302892,0.22645533,0.20302892,0.1796025,0.15617609,0.13665408,0.113227665,0.13665408,0.1639849,0.18741131,0.21083772,0.23816854,0.26159495,0.28111696,0.30454338,0.3279698,0.3513962,0.3474918,0.3435874,0.3435874,0.339683,0.3357786,0.29283017,0.24597734,0.20302892,0.15617609,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.38263142,0.76526284,1.1478943,1.5305257,1.9131571,3.0063896,4.095718,5.1889505,6.282183,7.375416,6.211904,5.0483923,3.8887846,2.7252727,1.5617609,1.2533131,0.94096094,0.63251317,0.3240654,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.1717937,0.1639849,0.16008049,0.15617609,0.14836729,0.13665408,0.12103647,0.10541886,0.08980125,0.07418364,0.08980125,0.10541886,0.12103647,0.13665408,0.14836729,0.12884527,0.10932326,0.08980125,0.07027924,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.3513962,0.6481308,0.94876975,1.2494087,1.5500476,1.261122,0.96829176,0.679366,0.39044023,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.08199245,0.1639849,0.24597734,0.3318742,0.41386664,0.39044023,0.3670138,0.3435874,0.3240654,0.30063897,0.359205,0.41386664,0.47243267,0.5309987,0.58566034,0.7027924,0.8160201,0.93315214,1.0463798,1.1635119,1.0463798,0.92924774,0.80821127,0.6910792,0.57394713,0.6949836,0.8160201,0.93315214,1.0541886,1.175225,1.5539521,1.9365835,2.3153105,2.6940374,3.076669,4.2284675,5.3841705,6.5398736,7.6955767,8.85128,7.1450562,5.4388323,3.736513,2.0302892,0.3240654,1.0190489,1.7140326,2.4090161,3.1039999,3.7989833,3.1313305,2.4597735,1.7882162,1.1205635,0.44900626,0.7066968,0.96438736,1.2220778,1.4797685,1.737459,1.7725986,1.8077383,1.8428779,1.8780174,1.9131571,2.2255092,2.5378613,2.8502135,3.1625657,3.474918,3.1079042,2.7408905,2.3738766,2.0068626,1.6359446,2.077142,2.5183394,2.9556324,3.39683,3.8380275,4.0761957,4.318269,4.5564375,4.7985106,5.036679,4.263607,3.4866312,2.7135596,1.9365835,1.1635119,0.97610056,0.79259366,0.60908675,0.42167544,0.23816854,0.19131571,0.14055848,0.093705654,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.21864653,0.31625658,0.40996224,0.5036679,0.60127795,0.5036679,0.40605783,0.30844778,0.21083772,0.113227665,0.113227665,0.113227665,0.113227665,0.113227665,0.113227665,0.10151446,0.093705654,0.08199245,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.03513962,0.058566034,0.078088045,0.10151446,0.12494087,0.14446288,0.1639849,0.1835069,0.20693332,0.22645533,0.25378615,0.28502136,0.31625658,0.3435874,0.37482262,0.40605783,0.44119745,0.47243267,0.5036679,0.5388075,0.60127795,0.6637484,0.7262188,0.78868926,0.8511597,0.94486535,1.038571,1.1361811,1.2298868,1.3235924,1.183034,1.038571,0.8980125,0.75354964,0.61299115,0.7301232,0.8472553,0.96438736,1.0815194,1.1986516,1.2962615,1.3899672,1.4836729,1.5812829,1.6749885,2.233318,2.795552,3.3538816,3.9161155,4.474445,4.4588275,4.4432096,4.4314966,4.415879,4.4002614,4.126953,3.853645,3.5842414,3.310933,3.0376248,2.7408905,2.4441557,2.1435168,1.8467822,1.5500476,1.3821584,1.2142692,1.0463798,0.8784905,0.7106012,0.6949836,0.679366,0.659844,0.6442264,0.62470436,0.5505207,0.47633708,0.39824903,0.3240654,0.24988174,0.26549935,0.28111696,0.29673457,0.30844778,0.3240654,0.47633708,0.62470436,0.77307165,0.92534333,1.0737107,1.1010414,1.1244678,1.1517987,1.175225,1.1986516,1.3743496,1.5461433,1.717937,1.8897307,2.0615244,1.7608855,1.456342,1.1557031,0.8511597,0.5505207,0.46071947,0.37482262,0.28892577,0.19912452,0.113227665,0.19131571,0.26940376,0.3435874,0.42167544,0.4997635,0.41777104,0.3357786,0.25378615,0.1717937,0.08589685,0.12884527,0.1717937,0.21474212,0.25769055,0.30063897,0.26940376,0.23816854,0.21083772,0.1796025,0.14836729,0.1756981,0.19912452,0.22645533,0.24988174,0.27330816,0.29283017,0.30844778,0.3279698,0.3435874,0.3631094,0.3670138,0.3709182,0.37872702,0.38263142,0.38653582,0.339683,0.29283017,0.24597734,0.19912452,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19912452,0.39824903,0.60127795,0.80040246,0.999527,2.5886188,4.173806,5.7628975,7.348085,8.937177,7.426173,5.911265,4.4002614,2.8892577,1.3743496,1.1010414,0.8238289,0.5505207,0.27330816,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.43729305,0.81211567,1.1869383,1.5617609,1.9365835,1.5734742,1.2142692,0.8511597,0.48805028,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.10151446,0.13665408,0.1756981,0.21083772,0.24988174,0.47633708,0.698888,0.92534333,1.1517987,1.3743496,1.1517987,0.92534333,0.698888,0.47633708,0.24988174,0.3240654,0.39824903,0.47633708,0.5505207,0.62470436,1.2376955,1.8506867,2.463678,3.076669,3.6857557,5.138193,6.5867267,8.039165,9.487698,10.936231,8.812236,6.688241,4.564246,2.436347,0.31235218,1.1986516,2.0888553,2.9751544,3.8614538,4.7516575,3.7989833,2.8502135,1.901444,0.94876975,0.0,0.113227665,0.22645533,0.3357786,0.44900626,0.5622339,0.76135844,0.96438736,1.1635119,1.3626363,1.5617609,2.0107672,2.463678,2.912684,3.3616903,3.8106966,3.3890212,2.9634414,2.5378613,2.1122816,1.6867018,2.0615244,2.436347,2.8111696,3.1859922,3.5608149,4.025439,4.4861584,4.950782,5.4115014,5.8761253,4.9624953,4.0488653,3.1391394,2.2255092,1.3118792,1.0737107,0.8394465,0.60127795,0.3631094,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.1639849,0.26159495,0.3631094,0.46071947,0.5622339,0.46071947,0.3631094,0.26159495,0.1639849,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.21083772,0.23816854,0.26159495,0.28892577,0.31235218,0.3631094,0.41386664,0.46071947,0.5114767,0.5622339,0.62470436,0.6871748,0.74964523,0.81211567,0.8745861,0.8745861,0.8745861,0.8745861,0.8745861,0.8745861,0.8238289,0.77307165,0.7262188,0.6754616,0.62470436,0.60127795,0.57394713,0.5505207,0.5231899,0.4997635,0.57394713,0.6481308,0.7262188,0.80040246,0.8745861,1.7608855,2.6510892,3.5373883,4.423688,5.3138914,5.001539,4.689187,4.376835,4.0605783,3.7482262,3.638903,3.5256753,3.4124475,3.2992198,3.1859922,2.8385005,2.4871042,2.135708,1.7882162,1.43682,1.261122,1.0893283,0.9136301,0.737932,0.5622339,0.4997635,0.43729305,0.37482262,0.31235218,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.26159495,0.46071947,0.6637484,0.8628729,1.0619974,1.0737107,1.0893283,1.1010414,1.1127546,1.1244678,1.3118792,1.4992905,1.6867018,1.8741131,2.0615244,1.7882162,1.5110037,1.2376955,0.96438736,0.6871748,0.57394713,0.46071947,0.3513962,0.23816854,0.12494087,0.22645533,0.3240654,0.42557985,0.5231899,0.62470436,0.5114767,0.39824903,0.28892577,0.1756981,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.37482262,0.3357786,0.30063897,0.26159495,0.22645533,0.18741131,0.21083772,0.23816854,0.26159495,0.28892577,0.31235218,0.3240654,0.3357786,0.3513962,0.3631094,0.37482262,0.38653582,0.39824903,0.41386664,0.42557985,0.43729305,0.38653582,0.3357786,0.28892577,0.23816854,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16008049,0.32016098,0.48024148,0.64032197,0.80040246,2.069333,3.338264,4.6110992,5.8800297,7.1489606,5.938596,4.728231,3.521771,2.3114061,1.1010414,0.8784905,0.659844,0.44119745,0.21864653,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.07027924,0.08980125,0.10932326,0.12884527,0.14836729,0.13274968,0.113227665,0.09761006,0.078088045,0.062470436,0.058566034,0.058566034,0.05466163,0.05075723,0.05075723,0.3513962,0.6481308,0.94876975,1.2494087,1.5500476,1.261122,0.96829176,0.679366,0.39044023,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.13665408,0.1717937,0.20693332,0.23816854,0.27330816,0.24988174,0.22645533,0.19912452,0.1756981,0.14836729,0.1835069,0.21864653,0.25378615,0.28892577,0.3240654,0.5114767,0.6949836,0.8784905,1.0659018,1.2494087,1.0424755,0.8355421,0.62860876,0.42167544,0.21083772,0.30454338,0.39824903,0.49195468,0.58175594,0.6754616,1.1400855,1.6047094,2.069333,2.533957,2.998581,4.181615,5.364649,6.547683,7.7307167,8.913751,7.211431,5.5130157,3.8106966,2.1122816,0.41386664,1.2415999,2.069333,2.893162,3.7208953,4.548629,3.6506162,2.7486992,1.8506867,0.94876975,0.05075723,0.12884527,0.21083772,0.28892577,0.3709182,0.44900626,0.60908675,0.76916724,0.92924774,1.0893283,1.2494087,1.737459,2.2255092,2.7135596,3.2016098,3.6857557,3.338264,2.9907722,2.6432803,2.2957885,1.9482968,2.436347,2.920493,3.4046388,3.8887846,4.376835,4.521298,4.6696653,4.8180323,4.9663997,5.1108627,4.3416953,3.5725281,2.803361,2.0341935,1.261122,1.077615,0.8941081,0.7066968,0.5231899,0.3357786,0.26940376,0.20302892,0.13665408,0.06637484,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.13274968,0.21474212,0.29673457,0.37872702,0.46071947,0.37872702,0.29673457,0.21474212,0.13274968,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.10151446,0.1756981,0.24988174,0.3240654,0.39824903,0.5192855,0.64032197,0.76135844,0.8784905,0.999527,1.116659,1.2337911,1.3509232,1.4719596,1.5890918,1.6008049,1.6164225,1.6320401,1.6476578,1.6632754,1.5969005,1.53443,1.4680552,1.4016805,1.33921,1.3235924,1.3079748,1.2923572,1.2767396,1.261122,1.2415999,1.2181735,1.1947471,1.1713207,1.1517987,1.1986516,1.2494087,1.3001659,1.3509232,1.4016805,1.2923572,1.1869383,1.077615,0.96829176,0.8628729,1.5929961,2.3231194,3.0532427,3.7833657,4.513489,4.3612175,4.21285,4.0605783,3.912211,3.7638438,3.6818514,3.6037633,3.521771,3.4436827,3.3616903,2.9751544,2.5886188,2.1981785,1.8116426,1.4251068,1.2415999,1.0580931,0.8784905,0.6949836,0.5114767,0.45681506,0.39824903,0.339683,0.28111696,0.22645533,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.3435874,0.5231899,0.7027924,0.8823949,1.0619974,1.1010414,1.1361811,1.175225,1.2142692,1.2494087,1.3860629,1.5188124,1.6554666,1.7882162,1.9248703,1.7491722,1.5695697,1.3938715,1.2142692,1.038571,0.91753453,0.79649806,0.679366,0.5583295,0.43729305,0.46852827,0.4958591,0.5270943,0.5583295,0.58566034,0.5700427,0.5544251,0.5349031,0.5192855,0.4997635,0.46071947,0.42557985,0.38653582,0.3513962,0.31235218,0.28892577,0.26159495,0.23816854,0.21083772,0.18741131,0.21864653,0.25378615,0.28502136,0.31625658,0.3513962,0.3631094,0.37872702,0.39434463,0.40996224,0.42557985,0.43729305,0.44900626,0.46071947,0.47633708,0.48805028,0.44900626,0.40605783,0.3670138,0.3279698,0.28892577,0.24597734,0.20693332,0.1678893,0.12884527,0.08589685,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12103647,0.23816854,0.359205,0.48024148,0.60127795,1.5539521,2.5066261,3.4593005,4.40807,5.3607445,4.454923,3.5491016,2.639376,1.7335546,0.8238289,0.659844,0.4958591,0.3318742,0.1639849,0.0,0.12103647,0.23816854,0.359205,0.48024148,0.60127795,0.48024148,0.359205,0.23816854,0.12103647,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.05075723,0.06637484,0.08199245,0.09761006,0.113227665,0.10151446,0.093705654,0.08199245,0.07418364,0.062470436,0.058566034,0.05075723,0.046852827,0.042948425,0.039044023,0.26159495,0.48805028,0.7106012,0.93705654,1.1635119,0.94486535,0.7262188,0.5114767,0.29283017,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.26940376,0.339683,0.40996224,0.48024148,0.5505207,0.48805028,0.42557985,0.3631094,0.30063897,0.23816854,0.26940376,0.30063897,0.3357786,0.3670138,0.39824903,0.5466163,0.6910792,0.8355421,0.98000497,1.1244678,0.93315214,0.74574083,0.5544251,0.3631094,0.1756981,0.28502136,0.39434463,0.5036679,0.61689556,0.7262188,1.0424755,1.358732,1.678893,1.9951496,2.3114061,3.2289407,4.142571,5.056201,5.9737353,6.8873653,5.610626,4.337791,3.0610514,1.7882162,0.5114767,1.2806439,2.0459068,2.815074,3.5842414,4.349504,3.4983444,2.6510892,1.7999294,0.94876975,0.10151446,0.14836729,0.19522011,0.24207294,0.28892577,0.3357786,0.45681506,0.57785153,0.698888,0.8160201,0.93705654,1.4641509,1.9873407,2.514435,3.0376248,3.5608149,3.2914112,3.0220075,2.7526035,2.4831998,2.2137961,2.8072653,3.4007344,3.998108,4.591577,5.1889505,5.0210614,4.853172,4.6852827,4.5173936,4.349504,3.7208953,3.096191,2.4675822,1.8389735,1.2142692,1.0815194,0.94876975,0.8160201,0.6832704,0.5505207,0.44119745,0.3318742,0.21864653,0.10932326,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.10151446,0.1678893,0.23426414,0.29673457,0.3631094,0.29673457,0.23426414,0.1678893,0.10151446,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.1756981,0.30063897,0.42557985,0.5505207,0.6754616,0.9019169,1.1283722,1.358732,1.5851873,1.8116426,2.0224805,2.233318,2.4441557,2.6510892,2.8619268,2.8424048,2.822883,2.803361,2.7838387,2.7643168,2.5690966,2.377781,2.1864653,1.9912452,1.7999294,1.7686942,1.7413634,1.7101282,1.678893,1.6515622,1.6554666,1.6593709,1.6632754,1.6710842,1.6749885,1.7999294,1.9248703,2.0498111,2.174752,2.2996929,2.0107672,1.7218413,1.4290112,1.1400855,0.8511597,1.4212024,1.9951496,2.5690966,3.1391394,3.7130866,3.7247996,3.736513,3.7482262,3.7638438,3.775557,3.7287042,3.6818514,3.631094,3.5842414,3.5373883,3.1118085,2.6862288,2.260649,1.8389735,1.4133936,1.2220778,1.0307622,0.8433509,0.6520352,0.46071947,0.40996224,0.359205,0.30454338,0.25378615,0.19912452,0.1756981,0.14836729,0.12494087,0.10151446,0.07418364,0.113227665,0.14836729,0.18741131,0.22645533,0.26159495,0.42167544,0.58175594,0.7418364,0.9019169,1.0619974,1.1244678,1.1869383,1.2494087,1.3118792,1.3743496,1.456342,1.5383345,1.6242313,1.7062237,1.7882162,1.7062237,1.6281357,1.5461433,1.4680552,1.3860629,1.261122,1.1322767,1.0034313,0.8784905,0.74964523,0.7106012,0.6715572,0.62860876,0.58956474,0.5505207,0.62860876,0.7066968,0.78088045,0.8589685,0.93705654,0.80040246,0.6637484,0.5231899,0.38653582,0.24988174,0.23816854,0.22645533,0.21083772,0.19912452,0.18741131,0.22645533,0.26940376,0.30844778,0.3474918,0.38653582,0.40605783,0.42167544,0.44119745,0.45681506,0.47633708,0.48805028,0.4997635,0.5114767,0.5231899,0.5388075,0.5075723,0.47633708,0.44900626,0.41777104,0.38653582,0.3435874,0.30063897,0.26159495,0.21864653,0.1756981,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,1.0346665,1.6710842,2.3035975,2.9400148,3.5764325,2.97125,2.366068,1.7608855,1.1557031,0.5505207,0.44119745,0.3318742,0.21864653,0.10932326,0.0,0.1796025,0.359205,0.5388075,0.71841,0.9019169,0.71841,0.5388075,0.359205,0.1796025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.03513962,0.046852827,0.05466163,0.06637484,0.07418364,0.07418364,0.07027924,0.06637484,0.06637484,0.062470436,0.05466163,0.046852827,0.039044023,0.031235218,0.023426414,0.1756981,0.3240654,0.47633708,0.62470436,0.77307165,0.62860876,0.48414588,0.339683,0.19522011,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.40605783,0.5114767,0.61689556,0.71841,0.8238289,0.7262188,0.62470436,0.5231899,0.42557985,0.3240654,0.3553006,0.38653582,0.41386664,0.44510186,0.47633708,0.58175594,0.6832704,0.78868926,0.8941081,0.999527,0.8277333,0.6559396,0.48414588,0.30844778,0.13665408,0.26549935,0.39434463,0.5192855,0.6481308,0.77307165,0.94486535,1.116659,1.2845483,1.456342,1.6242313,2.2723622,2.920493,3.5686235,4.2167544,4.860981,4.0137253,3.1625657,2.3114061,1.4641509,0.61299115,1.319688,2.0263848,2.7330816,3.4436827,4.1503797,3.349977,2.5495746,1.7491722,0.94876975,0.14836729,0.1639849,0.1796025,0.19522011,0.21083772,0.22645533,0.30454338,0.38653582,0.46462387,0.5466163,0.62470436,1.1869383,1.7491722,2.3114061,2.87364,3.435874,3.2445583,3.0532427,2.8619268,2.6667068,2.475391,3.1781836,3.8848803,4.591577,5.2943697,6.001066,5.5169206,5.036679,4.552533,4.068387,3.5881457,3.1039999,2.6159496,2.1318035,1.6476578,1.1635119,1.0815194,1.0034313,0.92143893,0.8433509,0.76135844,0.60908675,0.45681506,0.30454338,0.15227169,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.07418364,0.12103647,0.1678893,0.21474212,0.26159495,0.21474212,0.1678893,0.12103647,0.07418364,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.24988174,0.42557985,0.60127795,0.77307165,0.94876975,1.2845483,1.620327,1.9561055,2.2918842,2.6237583,2.9283018,3.2289407,3.533484,3.8341231,4.138666,4.084005,4.029343,3.970777,3.9161155,3.8614538,3.541293,3.2211318,2.900971,2.5808098,2.260649,2.2177005,2.1708477,2.1278992,2.0810463,2.0380979,2.069333,2.1005683,2.135708,2.1669433,2.1981785,2.4012074,2.6003318,2.7994564,2.998581,3.2016098,2.7291772,2.2567444,1.7843118,1.3118792,0.8394465,1.2533131,1.6671798,2.0810463,2.4988174,2.912684,3.0883822,3.2640803,3.435874,3.611572,3.78727,3.7716527,3.7560349,3.7443218,3.7287042,3.7130866,3.2484627,2.787743,2.3231194,1.8623998,1.4016805,1.2025559,1.0034313,0.80821127,0.60908675,0.41386664,0.3631094,0.31625658,0.26940376,0.22255093,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.113227665,0.1639849,0.21083772,0.26159495,0.31235218,0.3631094,0.5036679,0.6442264,0.78088045,0.92143893,1.0619974,1.1517987,1.2376955,1.3235924,1.4133936,1.4992905,1.5305257,1.5617609,1.5890918,1.620327,1.6515622,1.6671798,1.6867018,1.7023194,1.7218413,1.737459,1.6008049,1.4680552,1.3314011,1.1986516,1.0619974,0.95267415,0.8433509,0.7340276,0.62079996,0.5114767,0.6832704,0.8589685,1.0307622,1.2025559,1.3743496,1.1361811,0.9019169,0.6637484,0.42557985,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.23426414,0.28111696,0.3318742,0.37872702,0.42557985,0.44510186,0.46462387,0.48414588,0.5036679,0.5231899,0.5388075,0.5505207,0.5622339,0.57394713,0.58566034,0.5661383,0.5466163,0.5270943,0.5075723,0.48805028,0.44119745,0.39824903,0.3513962,0.30844778,0.26159495,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.5192855,0.8355421,1.1517987,1.4680552,1.7882162,1.4836729,1.183034,0.8784905,0.57785153,0.27330816,0.21864653,0.1639849,0.10932326,0.05466163,0.0,0.23816854,0.48024148,0.71841,0.96048295,1.1986516,0.96048295,0.71841,0.48024148,0.23816854,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.015617609,0.023426414,0.027330816,0.031235218,0.039044023,0.042948425,0.046852827,0.05075723,0.058566034,0.062470436,0.05075723,0.042948425,0.031235218,0.023426414,0.011713207,0.08589685,0.1639849,0.23816854,0.31235218,0.38653582,0.31625658,0.24207294,0.1717937,0.09761006,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,0.5388075,0.679366,0.8199245,0.96048295,1.1010414,0.96438736,0.8238289,0.6871748,0.5505207,0.41386664,0.44119745,0.46852827,0.4958591,0.5231899,0.5505207,0.61689556,0.679366,0.74574083,0.80821127,0.8745861,0.71841,0.5661383,0.40996224,0.25378615,0.10151446,0.24597734,0.39044023,0.5349031,0.679366,0.8238289,0.8472553,0.8706817,0.8941081,0.9136301,0.93705654,1.3157835,1.698415,2.077142,2.455869,2.8385005,2.4129205,1.9873407,1.5617609,1.1361811,0.7106012,1.358732,2.0068626,2.6549935,3.3031244,3.951255,3.2016098,2.4519646,1.698415,0.94876975,0.19912452,0.1835069,0.1639849,0.14836729,0.12884527,0.113227665,0.15227169,0.19131571,0.23426414,0.27330816,0.31235218,0.9136301,1.5110037,2.1122816,2.7135596,3.310933,3.1977055,3.0805733,2.9673457,2.854118,2.736986,3.5530062,4.369026,5.181142,5.997162,6.813182,6.016684,5.2162814,4.4197836,3.6232853,2.8267872,2.4831998,2.1396124,1.796025,1.456342,1.1127546,1.0854238,1.0580931,1.0307622,1.0034313,0.97610056,0.78088045,0.58566034,0.39044023,0.19522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.042948425,0.07418364,0.10151446,0.13274968,0.1639849,0.13274968,0.10151446,0.07418364,0.042948425,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.3240654,0.5505207,0.77307165,0.999527,1.2259823,1.6671798,2.1083772,2.5534792,2.9946766,3.435874,3.8341231,4.2284675,4.6228123,5.017157,5.4115014,5.3217,5.2318993,5.142098,5.0522966,4.9624953,4.513489,4.068387,3.619381,3.174279,2.7252727,2.6667068,2.6042364,2.5456703,2.4831998,2.4246337,2.4831998,2.5456703,2.6042364,2.6667068,2.7252727,2.998581,3.2757936,3.5491016,3.8263142,4.0996222,3.4436827,2.7916477,2.135708,1.4797685,0.8238289,1.0815194,1.33921,1.5969005,1.8545911,2.1122816,2.4480603,2.787743,3.1235218,3.4632049,3.7989833,3.8185053,3.8341231,3.853645,3.8692627,3.8887846,3.3890212,2.8892577,2.3855898,1.8858263,1.3860629,1.183034,0.97610056,0.77307165,0.5661383,0.3631094,0.32016098,0.27721256,0.23426414,0.19131571,0.14836729,0.14836729,0.14836729,0.14836729,0.14836729,0.14836729,0.21083772,0.27330816,0.3357786,0.39824903,0.46071947,0.58175594,0.7027924,0.8238289,0.94096094,1.0619974,1.175225,1.2884527,1.4016805,1.5110037,1.6242313,1.6008049,1.5812829,1.5578566,1.53443,1.5110037,1.6281357,1.7413634,1.8584955,1.9717231,2.0888553,1.9443923,1.8038338,1.6593709,1.5188124,1.3743496,1.1947471,1.0151446,0.8355421,0.6559396,0.47633708,0.7418364,1.0112402,1.2767396,1.5461433,1.8116426,1.475864,1.1361811,0.80040246,0.46071947,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.24207294,0.29673457,0.3513962,0.40605783,0.46071947,0.48414588,0.5075723,0.5309987,0.5544251,0.57394713,0.58566034,0.60127795,0.61299115,0.62470436,0.63641757,0.62860876,0.61689556,0.60908675,0.59737355,0.58566034,0.5388075,0.49195468,0.44510186,0.39824903,0.3513962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.30063897,0.60127795,0.9019169,1.1986516,1.4992905,1.1986516,0.9019169,0.60127795,0.30063897,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.6754616,0.8511597,1.0268579,1.1986516,1.3743496,1.1986516,1.0268579,0.8511597,0.6754616,0.4997635,0.5231899,0.5505207,0.57394713,0.60127795,0.62470436,0.6481308,0.6754616,0.698888,0.7262188,0.74964523,0.61299115,0.47633708,0.3357786,0.19912452,0.062470436,0.22645533,0.38653582,0.5505207,0.7106012,0.8745861,0.74964523,0.62470436,0.4997635,0.37482262,0.24988174,0.3631094,0.47633708,0.58566034,0.698888,0.81211567,0.81211567,0.81211567,0.81211567,0.81211567,0.81211567,1.4016805,1.9873407,2.5769055,3.1625657,3.7482262,3.049338,2.35045,1.6515622,0.94876975,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.63641757,1.2767396,1.9131571,2.5495746,3.1859922,3.1508527,3.1118085,3.076669,3.0376248,2.998581,3.9239242,4.8492675,5.774611,6.699954,7.6252975,6.5125427,5.3997884,4.2870336,3.174279,2.0615244,1.8623998,1.6632754,1.4641509,1.261122,1.0619974,1.0893283,1.1127546,1.1361811,1.1635119,1.1869383,0.94876975,0.7106012,0.47633708,0.23816854,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.39824903,0.6754616,0.94876975,1.2259823,1.4992905,2.0498111,2.6003318,3.1508527,3.7013733,4.251894,4.73604,5.22409,5.7121406,6.2001905,6.688241,6.5633,6.4383593,6.3134184,6.1884775,6.0635366,5.4856853,4.911738,4.337791,3.7638438,3.1859922,3.1118085,3.0376248,2.9634414,2.8892577,2.8111696,2.900971,2.9868677,3.076669,3.1625657,3.2484627,3.5998588,3.951255,4.298747,4.650143,5.001539,4.1620927,3.3265507,2.4871042,1.6515622,0.81211567,0.9136301,1.0112402,1.1127546,1.2142692,1.3118792,1.8116426,2.3114061,2.8111696,3.310933,3.8106966,3.8614538,3.912211,3.9629683,4.0137253,4.0605783,3.5256753,2.9868677,2.4480603,1.9131571,1.3743496,1.1635119,0.94876975,0.737932,0.5231899,0.31235218,0.27330816,0.23816854,0.19912452,0.1639849,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.26159495,0.3357786,0.41386664,0.48805028,0.5622339,0.6637484,0.76135844,0.8628729,0.96438736,1.0619974,1.1986516,1.33921,1.475864,1.6125181,1.7491722,1.6749885,1.6008049,1.5266213,1.4485333,1.3743496,1.5890918,1.7999294,2.0107672,2.2255092,2.436347,2.2879796,2.135708,1.9873407,1.8389735,1.6867018,1.43682,1.1869383,0.93705654,0.6871748,0.43729305,0.80040246,1.1635119,1.5266213,1.8858263,2.2489357,1.8116426,1.3743496,0.93705654,0.4997635,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.24988174,0.31235218,0.37482262,0.43729305,0.4997635,0.5231899,0.5505207,0.57394713,0.60127795,0.62470436,0.63641757,0.6481308,0.6637484,0.6754616,0.6871748,0.6871748,0.6871748,0.6871748,0.6871748,0.6871748,0.63641757,0.58566034,0.5388075,0.48805028,0.43729305,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23816854,0.48024148,0.71841,0.96048295,1.1986516,0.96048295,0.71841,0.48024148,0.23816854,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08199245,0.1639849,0.24597734,0.3318742,0.41386664,0.5505207,0.6871748,0.8238289,0.96438736,1.1010414,0.96438736,0.8238289,0.6871748,0.5505207,0.41386664,0.42948425,0.44900626,0.46462387,0.48414588,0.4997635,0.5231899,0.5466163,0.5661383,0.58956474,0.61299115,0.5270943,0.44119745,0.359205,0.27330816,0.18741131,0.30844778,0.43338865,0.5544251,0.679366,0.80040246,0.7027924,0.60518235,0.5075723,0.40996224,0.31235218,0.5466163,0.77697605,1.0112402,1.2415999,1.475864,1.3782539,1.2845483,1.1908426,1.0932326,0.999527,1.456342,1.9092526,2.366068,2.8189783,3.2757936,2.7565079,2.233318,1.7140326,1.1947471,0.6754616,0.5466163,0.41386664,0.28502136,0.15617609,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.5661383,1.1283722,1.6945106,2.260649,2.8267872,2.8619268,2.893162,2.9283018,2.9634414,2.998581,3.7013733,4.4002614,5.099149,5.801942,6.5008297,5.591104,4.6813784,3.7716527,2.8619268,1.9482968,1.7608855,1.5695697,1.3782539,1.1908426,0.999527,0.9917182,0.98390937,0.97610056,0.96829176,0.96438736,0.77307165,0.58566034,0.39824903,0.21083772,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.3240654,0.5466163,0.76916724,0.9917182,1.2142692,1.6632754,2.1161861,2.5690966,3.0220075,3.474918,3.8809757,4.290938,4.6969957,5.1030536,5.5130157,5.423215,5.337318,5.251421,5.1616197,5.0757227,4.6696653,4.263607,3.8614538,3.455396,3.049338,3.06886,3.084478,3.1039999,3.1196175,3.1391394,3.1118085,3.0883822,3.0610514,3.0376248,3.0141985,3.2953155,3.5764325,3.8614538,4.142571,4.423688,3.8341231,3.240654,2.6471848,2.0537157,1.4641509,1.5383345,1.6125181,1.6867018,1.7608855,1.8389735,2.3465457,2.854118,3.3616903,3.8692627,4.376835,4.154284,3.9317331,3.7091823,3.4866312,3.2640803,2.8306916,2.4012074,1.9717231,1.542239,1.1127546,0.94096094,0.76916724,0.59346914,0.42167544,0.24988174,0.21864653,0.19131571,0.16008049,0.12884527,0.10151446,0.113227665,0.12494087,0.13665408,0.14836729,0.1639849,0.22255093,0.28111696,0.3435874,0.40215343,0.46071947,0.5466163,0.63251317,0.71841,0.80430686,0.8862993,1.0151446,1.1439898,1.2689307,1.397776,1.5266213,1.5110037,1.4953861,1.4797685,1.4641509,1.4485333,1.6827974,1.9131571,2.1474214,2.3816853,2.612045,2.5573835,2.5027218,2.4480603,2.3933985,2.338737,2.018576,1.7023194,1.3860629,1.0659018,0.74964523,1.0737107,1.4016805,1.7257458,2.0498111,2.3738766,2.084951,1.796025,1.5031948,1.2142692,0.92534333,0.77697605,0.62860876,0.48414588,0.3357786,0.18741131,0.25378615,0.31625658,0.38263142,0.44900626,0.5114767,0.5270943,0.5427119,0.5583295,0.57394713,0.58566034,0.61689556,0.6442264,0.6715572,0.698888,0.7262188,0.7301232,0.7340276,0.7418364,0.74574083,0.74964523,0.698888,0.6481308,0.60127795,0.5505207,0.4997635,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1796025,0.359205,0.5388075,0.71841,0.9019169,0.71841,0.5388075,0.359205,0.1796025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06637484,0.12884527,0.19522011,0.26159495,0.3240654,0.42557985,0.5231899,0.62470436,0.7262188,0.8238289,0.7262188,0.62470436,0.5231899,0.42557985,0.3240654,0.3357786,0.3435874,0.3553006,0.3631094,0.37482262,0.39434463,0.41386664,0.43338865,0.45681506,0.47633708,0.44119745,0.40996224,0.37872702,0.3435874,0.31235218,0.39434463,0.47633708,0.5583295,0.6442264,0.7262188,0.6559396,0.58566034,0.5153811,0.44510186,0.37482262,0.7262188,1.0815194,1.4329157,1.7843118,2.135708,1.9482968,1.756981,1.5656652,1.3782539,1.1869383,1.5110037,1.8311646,2.15523,2.4792955,2.7994564,2.4597735,2.1200905,1.7804074,1.4407244,1.1010414,0.8902037,0.679366,0.46852827,0.26159495,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.49195468,0.98390937,1.475864,1.9717231,2.463678,2.5690966,2.67842,2.7838387,2.893162,2.998581,3.474918,3.951255,4.423688,4.900025,5.376362,4.6657605,3.959064,3.252367,2.5456703,1.8389735,1.6593709,1.475864,1.2962615,1.116659,0.93705654,0.8980125,0.8589685,0.8160201,0.77697605,0.737932,0.60127795,0.46071947,0.3240654,0.18741131,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.24597734,0.41386664,0.58566034,0.75354964,0.92534333,1.2806439,1.6359446,1.9912452,2.3465457,2.7018464,3.0259118,3.3538816,3.6818514,4.009821,4.337791,4.2870336,4.2362766,4.1894236,4.138666,4.087909,3.853645,3.619381,3.3812122,3.1469483,2.912684,3.0220075,3.1313305,3.240654,3.3538816,3.4632049,3.3265507,3.1859922,3.049338,2.912684,2.77603,2.9907722,3.2055142,3.4202564,3.6349986,3.8497405,3.5022488,3.154757,2.8072653,2.4597735,2.1122816,2.1630387,2.2137961,2.260649,2.3114061,2.3621633,2.8775444,3.3929255,3.9083066,4.423688,4.939069,4.4432096,3.9473507,3.4514916,2.9556324,2.463678,2.1396124,1.8194515,1.4953861,1.1713207,0.8511597,0.71841,0.58566034,0.45291066,0.32016098,0.18741131,0.1639849,0.14055848,0.12103647,0.09761006,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.13665408,0.1835069,0.22645533,0.27330816,0.31625658,0.3631094,0.43338865,0.5036679,0.57394713,0.6442264,0.7106012,0.8316377,0.94876975,1.0659018,1.183034,1.3001659,1.3431144,1.3899672,1.43682,1.4797685,1.5266213,1.7765031,2.0302892,2.2840753,2.533957,2.787743,2.8267872,2.8658314,2.9087796,2.9478238,2.9868677,2.6042364,2.2177005,1.8311646,1.4485333,1.0619974,1.3509232,1.6359446,1.9248703,2.2137961,2.4988174,2.358259,2.2137961,2.0732377,1.9287747,1.7882162,1.4680552,1.1478943,0.8277333,0.5075723,0.18741131,0.25378615,0.3240654,0.39044023,0.45681506,0.5231899,0.5309987,0.5349031,0.5388075,0.5466163,0.5505207,0.59346914,0.63641757,0.679366,0.71841,0.76135844,0.77307165,0.78088045,0.79259366,0.80430686,0.81211567,0.76135844,0.7106012,0.6637484,0.61299115,0.5622339,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12103647,0.23816854,0.359205,0.48024148,0.60127795,0.48024148,0.359205,0.23816854,0.12103647,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.093705654,0.14055848,0.19131571,0.23816854,0.30063897,0.3631094,0.42557985,0.48805028,0.5505207,0.48805028,0.42557985,0.3631094,0.30063897,0.23816854,0.23816854,0.24207294,0.24597734,0.24597734,0.24988174,0.26940376,0.28502136,0.30063897,0.32016098,0.3357786,0.359205,0.37872702,0.39824903,0.41777104,0.43729305,0.48024148,0.5231899,0.5661383,0.60908675,0.6481308,0.60908675,0.5661383,0.5231899,0.48024148,0.43729305,0.9097257,1.3821584,1.8545911,2.3270237,2.7994564,2.514435,2.2294137,1.9443923,1.6593709,1.3743496,1.5656652,1.7530766,1.9443923,2.135708,2.3231194,2.1669433,2.0068626,1.8467822,1.6867018,1.5266213,1.2337911,0.94486535,0.6559396,0.3631094,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.42167544,0.8394465,1.261122,1.678893,2.1005683,2.280171,2.4597735,2.639376,2.8189783,2.998581,3.2484627,3.4983444,3.7482262,3.998108,4.251894,3.7443218,3.240654,2.7330816,2.2294137,1.7257458,1.5539521,1.3860629,1.2142692,1.0463798,0.8745861,0.80430686,0.7301232,0.6559396,0.58566034,0.5114767,0.42557985,0.3357786,0.24988174,0.1639849,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.1678893,0.28502136,0.40215343,0.5192855,0.63641757,0.8941081,1.1517987,1.4094892,1.6671798,1.9248703,2.1708477,2.4207294,2.6667068,2.9165885,3.1625657,3.1508527,3.1391394,3.1235218,3.1118085,3.1000953,3.0337205,2.97125,2.9048753,2.8385005,2.77603,2.979059,3.1781836,3.3812122,3.5842414,3.78727,3.5373883,3.2875066,3.0376248,2.787743,2.5378613,2.6862288,2.8306916,2.979059,3.1274261,3.2757936,3.174279,3.06886,2.9673457,2.8658314,2.7643168,2.787743,2.8111696,2.8385005,2.8619268,2.8892577,3.408543,3.9317331,4.454923,4.9781127,5.5013027,4.732136,3.9668727,3.1977055,2.4285383,1.6632754,1.4485333,1.2337911,1.0190489,0.80430686,0.58566034,0.4958591,0.40215343,0.30844778,0.21864653,0.12494087,0.10932326,0.093705654,0.078088045,0.06637484,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.14055848,0.1717937,0.20302892,0.23426414,0.26159495,0.31625658,0.3709182,0.42557985,0.48414588,0.5388075,0.6442264,0.75354964,0.8589685,0.96829176,1.0737107,1.1791295,1.2845483,1.3899672,1.4953861,1.6008049,1.8741131,2.1435168,2.416825,2.690133,2.9634414,3.096191,3.232845,3.3655949,3.5022488,3.638903,3.1859922,2.7330816,2.280171,1.8272603,1.3743496,1.6242313,1.8741131,2.1239948,2.3738766,2.6237583,2.631567,2.6354716,2.639376,2.6432803,2.6510892,2.1591344,1.6632754,1.1713207,0.679366,0.18741131,0.25769055,0.3279698,0.39824903,0.46852827,0.5388075,0.5309987,0.5270943,0.5231899,0.5192855,0.5114767,0.5700427,0.62860876,0.6832704,0.7418364,0.80040246,0.8160201,0.8316377,0.8433509,0.8589685,0.8745861,0.8238289,0.77307165,0.7262188,0.6754616,0.62470436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.1756981,0.19912452,0.22645533,0.24988174,0.27330816,0.24988174,0.22645533,0.19912452,0.1756981,0.14836729,0.14446288,0.14055848,0.13665408,0.12884527,0.12494087,0.14055848,0.15617609,0.1717937,0.1835069,0.19912452,0.27330816,0.3435874,0.41777104,0.48805028,0.5622339,0.5661383,0.5661383,0.5700427,0.57394713,0.57394713,0.5583295,0.5466163,0.5309987,0.5153811,0.4997635,1.0932326,1.6867018,2.2762666,2.8697357,3.4632049,3.0805733,2.7018464,2.3231194,1.9443923,1.5617609,1.620327,1.678893,1.7335546,1.7921207,1.8506867,1.8702087,1.8897307,1.9092526,1.9287747,1.9482968,1.5812829,1.2103647,0.8394465,0.46852827,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.3474918,0.6949836,1.0424755,1.3899672,1.737459,1.9912452,2.241127,2.494913,2.7486992,2.998581,3.0259118,3.049338,3.076669,3.1000953,3.1235218,2.822883,2.5183394,2.2177005,1.9131571,1.6125181,1.4524376,1.2923572,1.1322767,0.97219616,0.81211567,0.7066968,0.60127795,0.4958591,0.39434463,0.28892577,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.08980125,0.15617609,0.21864653,0.28502136,0.3513962,0.5114767,0.6715572,0.8316377,0.9917182,1.1517987,1.3157835,1.4836729,1.6515622,1.8194515,1.9873407,2.0107672,2.0380979,2.0615244,2.0888553,2.1122816,2.2177005,2.3231194,2.4285383,2.533957,2.639376,2.9322062,3.2289407,3.521771,3.8185053,4.1113358,3.7482262,3.3890212,3.0259118,2.6628022,2.2996929,2.3816853,2.4597735,2.541766,2.619854,2.7018464,2.8424048,2.9868677,3.1274261,3.2718892,3.4124475,3.4124475,3.4124475,3.4124475,3.4124475,3.4124475,3.9434462,4.4705405,5.001539,5.532538,6.0635366,5.0210614,3.9824903,2.9439192,1.901444,0.8628729,0.75354964,0.6481308,0.5388075,0.43338865,0.3240654,0.27330816,0.21864653,0.1678893,0.113227665,0.062470436,0.05466163,0.046852827,0.039044023,0.031235218,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.11713207,0.13274968,0.14836729,0.1639849,0.20302892,0.24207294,0.28111696,0.3240654,0.3631094,0.46071947,0.5583295,0.6559396,0.75354964,0.8511597,1.0151446,1.1791295,1.3431144,1.5110037,1.6749885,1.9678187,2.260649,2.5534792,2.8463092,3.1391394,3.3655949,3.5959544,3.8263142,4.056674,4.2870336,3.767748,3.2484627,2.7291772,2.2059872,1.6867018,1.901444,2.1122816,2.3231194,2.5378613,2.7486992,2.900971,3.0532427,3.2094188,3.3616903,3.513962,2.8463092,2.182561,1.5188124,0.8511597,0.18741131,0.26159495,0.3318742,0.40605783,0.47633708,0.5505207,0.5349031,0.5192855,0.5036679,0.48805028,0.47633708,0.5466163,0.62079996,0.6910792,0.76526284,0.8394465,0.8589685,0.8784905,0.8980125,0.91753453,0.93705654,0.8862993,0.8394465,0.78868926,0.737932,0.6871748,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.18741131,0.31235218,0.43729305,0.5622339,0.6871748,0.6481308,0.61299115,0.57394713,0.5388075,0.4997635,0.5114767,0.5231899,0.5388075,0.5505207,0.5622339,1.2767396,1.9873407,2.7018464,3.4124475,4.123049,3.6506162,3.174279,2.7018464,2.2255092,1.7491722,1.6749885,1.6008049,1.5266213,1.4485333,1.3743496,1.5734742,1.7765031,1.9756275,2.174752,2.3738766,1.9248703,1.475864,1.0268579,0.57394713,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.27330816,0.5505207,0.8238289,1.1010414,1.3743496,1.698415,2.0263848,2.35045,2.6745155,2.998581,2.7994564,2.6003318,2.4012074,2.1981785,1.999054,1.901444,1.7999294,1.698415,1.6008049,1.4992905,1.3509232,1.1986516,1.0502841,0.9019169,0.74964523,0.61299115,0.47633708,0.3357786,0.19912452,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.37482262,0.46071947,0.5505207,0.63641757,0.7262188,0.81211567,0.8745861,0.93705654,0.999527,1.0619974,1.1244678,1.4016805,1.6749885,1.9482968,2.2255092,2.4988174,2.8892577,3.2757936,3.6623292,4.0488653,4.4393053,3.9629683,3.4866312,3.0141985,2.5378613,2.0615244,2.0732377,2.0888553,2.1005683,2.1122816,2.1239948,2.514435,2.900971,3.2875066,3.6740425,4.0605783,4.037152,4.0137253,3.9863946,3.9629683,3.9356375,4.474445,5.0132523,5.548156,6.086963,6.6257706,5.3138914,3.998108,2.6862288,1.3743496,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.27330816,0.3631094,0.44900626,0.5388075,0.62470436,0.8511597,1.0737107,1.3001659,1.5266213,1.7491722,2.0615244,2.3738766,2.6862288,2.998581,3.310933,3.638903,3.9629683,4.2870336,4.6110992,4.939069,4.349504,3.7638438,3.174279,2.5886188,1.999054,2.174752,2.35045,2.5261483,2.7018464,2.87364,3.174279,3.474918,3.775557,4.0761957,4.376835,3.5373883,2.7018464,1.8623998,1.0268579,0.18741131,0.26159495,0.3357786,0.41386664,0.48805028,0.5622339,0.5388075,0.5114767,0.48805028,0.46071947,0.43729305,0.5231899,0.61299115,0.698888,0.78868926,0.8745861,0.9019169,0.92534333,0.94876975,0.97610056,0.999527,0.94876975,0.9019169,0.8511597,0.80040246,0.74964523,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.1639849,0.27330816,0.38653582,0.4997635,0.61299115,0.60127795,0.58566034,0.57394713,0.5622339,0.5505207,0.6559396,0.76135844,0.8667773,0.96829176,1.0737107,1.6710842,2.2645533,2.8619268,3.455396,4.0488653,3.611572,3.174279,2.736986,2.2996929,1.8623998,1.8038338,1.7413634,1.6827974,1.6242313,1.5617609,1.8311646,2.096664,2.366068,2.631567,2.900971,2.436347,1.9756275,1.5110037,1.0502841,0.58566034,0.5505207,0.5114767,0.47633708,0.43729305,0.39824903,0.5427119,0.6832704,0.8277333,0.96829176,1.1127546,1.3743496,1.6320401,1.893635,2.1513257,2.4129205,2.2879796,2.1630387,2.0380979,1.9131571,1.7882162,1.8194515,1.8467822,1.8780174,1.9092526,1.9365835,1.7413634,1.542239,1.3431144,1.1478943,0.94876975,0.8238289,0.6949836,0.5661383,0.44119745,0.31235218,0.28111696,0.25378615,0.22255093,0.19131571,0.1639849,0.13665408,0.10932326,0.078088045,0.05075723,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.30063897,0.38263142,0.46462387,0.5466163,0.62860876,0.7106012,0.78868926,0.8667773,0.94486535,1.0229534,1.1010414,1.4172981,1.7335546,2.0537157,2.3699722,2.6862288,3.076669,3.4671092,3.8575494,4.2479897,4.6384296,4.415879,4.1972322,3.978586,3.7560349,3.5373883,3.3812122,3.2211318,3.0649557,2.9087796,2.7486992,3.1079042,3.4632049,3.8224099,4.181615,4.5369153,4.4119744,4.2870336,4.1620927,4.037152,3.912211,4.220659,4.533011,4.841459,5.153811,5.462259,4.388548,3.3187418,2.2450314,1.1713207,0.10151446,0.093705654,0.08980125,0.08589685,0.078088045,0.07418364,0.06637484,0.05466163,0.046852827,0.03513962,0.023426414,0.031235218,0.039044023,0.046852827,0.05466163,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.25769055,0.3279698,0.39824903,0.46852827,0.5388075,0.737932,0.93705654,1.1361811,1.33921,1.5383345,1.8350691,2.1318035,2.4285383,2.7291772,3.0259118,3.3460727,3.6701381,3.9942036,4.3143644,4.6384296,4.271416,3.9044023,3.533484,3.1664703,2.7994564,2.8385005,2.87364,2.912684,2.951728,2.9868677,3.2992198,3.611572,3.9239242,4.2362766,4.548629,3.8692627,3.1859922,2.5027218,1.8194515,1.1361811,1.0463798,0.95267415,0.8589685,0.76916724,0.6754616,0.63251317,0.58956474,0.5466163,0.5036679,0.46071947,0.5231899,0.58175594,0.6442264,0.7027924,0.76135844,0.79259366,0.8238289,0.8511597,0.8823949,0.9136301,0.9019169,0.8941081,0.8823949,0.8706817,0.8628729,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.13665408,0.23816854,0.3357786,0.43729305,0.5388075,0.5505207,0.5622339,0.57394713,0.58566034,0.60127795,0.79649806,0.9956226,1.1908426,1.3899672,1.5890918,2.0654287,2.541766,3.018103,3.4983444,3.9746814,3.5764325,3.174279,2.77603,2.3738766,1.9756275,1.9287747,1.8858263,1.8389735,1.796025,1.7491722,2.084951,2.4207294,2.7565079,3.0883822,3.4241607,2.951728,2.475391,1.999054,1.5266213,1.0502841,0.999527,0.94876975,0.9019169,0.8511597,0.80040246,0.80821127,0.8199245,0.8316377,0.8394465,0.8511597,1.0463798,1.2415999,1.43682,1.6281357,1.8233559,1.7765031,1.7257458,1.6749885,1.6242313,1.5734742,1.7335546,1.893635,2.0537157,2.2137961,2.3738766,2.1318035,1.8858263,1.639849,1.3938715,1.1517987,1.0307622,0.9136301,0.79649806,0.679366,0.5622339,0.48805028,0.41777104,0.3435874,0.27330816,0.19912452,0.1717937,0.14055848,0.10932326,0.078088045,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.22645533,0.30063897,0.37872702,0.45681506,0.5349031,0.61299115,0.7066968,0.79649806,0.8902037,0.98390937,1.0737107,1.43682,1.796025,2.15523,2.514435,2.87364,3.2679846,3.6584249,4.0527697,4.4432096,4.8375545,4.872694,4.9078336,4.942973,4.9781127,5.0132523,4.6852827,4.357313,4.029343,3.7013733,3.3734035,3.7013733,4.029343,4.357313,4.6852827,5.0132523,4.786797,4.564246,4.337791,4.1113358,3.8887846,3.970777,4.0527697,4.134762,4.2167544,4.298747,3.4671092,2.6354716,1.8038338,0.96829176,0.13665408,0.12884527,0.11713207,0.10932326,0.09761006,0.08589685,0.078088045,0.07418364,0.06637484,0.058566034,0.05075723,0.06637484,0.078088045,0.093705654,0.10932326,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.23816854,0.29283017,0.3435874,0.39824903,0.44900626,0.62470436,0.80040246,0.97610056,1.1517987,1.3235924,1.6086137,1.8897307,2.1708477,2.455869,2.736986,3.057147,3.377308,3.697469,4.01763,4.337791,4.1894236,4.041056,3.8965936,3.7482262,3.5998588,3.4983444,3.4007344,3.2992198,3.2016098,3.1000953,3.4241607,3.7482262,4.0761957,4.4002614,4.7243266,4.1972322,3.6701381,3.1430438,2.6159496,2.0888553,1.8272603,1.5656652,1.3079748,1.0463798,0.78868926,0.7262188,0.6676528,0.60908675,0.5466163,0.48805028,0.5192855,0.5544251,0.58566034,0.61689556,0.6481308,0.6832704,0.71841,0.75354964,0.78868926,0.8238289,0.8550641,0.8862993,0.9136301,0.94486535,0.97610056,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.113227665,0.19912452,0.28892577,0.37482262,0.46071947,0.4997635,0.5388075,0.57394713,0.61299115,0.6481308,0.94096094,1.2298868,1.5188124,1.8116426,2.1005683,2.4597735,2.8189783,3.1781836,3.541293,3.900498,3.5373883,3.174279,2.8111696,2.4480603,2.0888553,2.05762,2.0263848,1.999054,1.9678187,1.9365835,2.338737,2.7408905,3.1469483,3.5491016,3.951255,3.4632049,2.9751544,2.4871042,1.999054,1.5110037,1.4485333,1.3860629,1.3235924,1.261122,1.1986516,1.077615,0.95657855,0.8316377,0.7106012,0.58566034,0.71841,0.8472553,0.97610056,1.1088502,1.2376955,1.261122,1.2884527,1.3118792,1.33921,1.3626363,1.6515622,1.9443923,2.233318,2.522244,2.8111696,2.5183394,2.2294137,1.9365835,1.6437533,1.3509232,1.2415999,1.1361811,1.0268579,0.92143893,0.81211567,0.698888,0.58175594,0.46852827,0.3513962,0.23816854,0.20693332,0.1717937,0.14055848,0.10932326,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.22255093,0.29673457,0.3670138,0.44119745,0.5114767,0.62079996,0.7262188,0.8355421,0.94096094,1.0502841,1.4524376,1.8545911,2.2567444,2.6588979,3.0610514,3.4593005,3.853645,4.2479897,4.6423345,5.036679,5.3256044,5.618435,5.9073606,6.196286,6.4891167,5.989353,5.493494,4.9937305,4.4978714,3.998108,4.298747,4.5954814,4.892216,5.1889505,5.4856853,5.1616197,4.8375545,4.513489,4.1894236,3.8614538,3.716991,3.5725281,3.4280653,3.2836022,3.1391394,2.5456703,1.9522011,1.358732,0.76916724,0.1756981,0.16008049,0.14446288,0.12884527,0.113227665,0.10151446,0.093705654,0.08980125,0.08589685,0.078088045,0.07418364,0.09761006,0.12103647,0.14055848,0.1639849,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.23816854,0.22645533,0.21083772,0.19912452,0.18741131,0.22255093,0.25769055,0.29283017,0.3279698,0.3631094,0.5114767,0.6637484,0.81211567,0.96438736,1.1127546,1.3782539,1.6476578,1.9131571,2.182561,2.4480603,2.7682211,3.084478,3.4007344,3.7208953,4.037152,4.1113358,4.181615,4.2557983,4.3260775,4.4002614,4.1620927,3.9239242,3.6857557,3.4514916,3.213323,3.5491016,3.8887846,4.224563,4.564246,4.900025,4.5291066,4.154284,3.7833657,3.408543,3.0376248,2.6081407,2.182561,1.7530766,1.3274968,0.9019169,0.8238289,0.74574083,0.6676528,0.58956474,0.5114767,0.5192855,0.5231899,0.5270943,0.5309987,0.5388075,0.57785153,0.61689556,0.6559396,0.698888,0.737932,0.80821127,0.8784905,0.94876975,1.0190489,1.0893283,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.08589685,0.1639849,0.23816854,0.31235218,0.38653582,0.44900626,0.5114767,0.57394713,0.63641757,0.698888,1.0815194,1.4641509,1.8467822,2.2294137,2.612045,2.854118,3.096191,3.338264,3.5842414,3.8263142,3.4983444,3.174279,2.8502135,2.5261483,2.1981785,2.1864653,2.1708477,2.15523,2.1396124,2.1239948,2.5964274,3.0649557,3.533484,4.0059166,4.474445,3.9746814,3.474918,2.9751544,2.475391,1.9756275,1.901444,1.8233559,1.7491722,1.6749885,1.6008049,1.3431144,1.0893283,0.8355421,0.58175594,0.3240654,0.39044023,0.45681506,0.5192855,0.58566034,0.6481308,0.74964523,0.8511597,0.94876975,1.0502841,1.1517987,1.5695697,1.9912452,2.4090161,2.8306916,3.2484627,2.9087796,2.5690966,2.2294137,1.8897307,1.5500476,1.4524376,1.3548276,1.2572175,1.1596074,1.0619974,0.9058213,0.74574083,0.58956474,0.43338865,0.27330816,0.23816854,0.20693332,0.1717937,0.13665408,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.14055848,0.21083772,0.27721256,0.3435874,0.41386664,0.5349031,0.6559396,0.78088045,0.9019169,1.0268579,1.4719596,1.9131571,2.358259,2.803361,3.2484627,3.6467118,4.044961,4.4432096,4.841459,5.2358036,5.7824197,6.329036,6.871748,7.4183645,7.9610763,7.2934237,6.6257706,5.958118,5.2943697,4.6267166,4.892216,5.1616197,5.4271193,5.6965227,5.9620223,5.5364423,5.1108627,4.689187,4.263607,3.8380275,3.4632049,3.0922866,2.7213683,2.3465457,1.9756275,1.6242313,1.2689307,0.91753453,0.5661383,0.21083772,0.19131571,0.1717937,0.15227169,0.13274968,0.113227665,0.10932326,0.10932326,0.10541886,0.10151446,0.10151446,0.12884527,0.16008049,0.19131571,0.21864653,0.24988174,0.26159495,0.27330816,0.28892577,0.30063897,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.28892577,0.26159495,0.23816854,0.21083772,0.18741131,0.20693332,0.22255093,0.23816854,0.25769055,0.27330816,0.39824903,0.5231899,0.6481308,0.77307165,0.9019169,1.1517987,1.4055848,1.6593709,1.9092526,2.1630387,2.4792955,2.7916477,3.1079042,3.4241607,3.736513,4.029343,4.322173,4.6150036,4.9078336,5.2006636,4.825841,4.4510183,4.0761957,3.7013733,3.3265507,3.6740425,4.025439,4.376835,4.7243266,5.0757227,4.8570766,4.6384296,4.423688,4.2050414,3.9863946,3.3929255,2.795552,2.2020829,1.6086137,1.0112402,0.91753453,0.8238289,0.7262188,0.63251317,0.5388075,0.5153811,0.49195468,0.46852827,0.44900626,0.42557985,0.46852827,0.5153811,0.5583295,0.60518235,0.6481308,0.76135844,0.8706817,0.98000497,1.0893283,1.1986516,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.39824903,0.48805028,0.57394713,0.6637484,0.74964523,1.2259823,1.698415,2.174752,2.6510892,3.1235218,3.2484627,3.3734035,3.4983444,3.6232853,3.7482262,3.4632049,3.174279,2.8892577,2.6003318,2.3114061,2.3114061,2.3114061,2.3114061,2.3114061,2.3114061,2.8502135,3.3890212,3.9239242,4.462732,5.001539,4.4861584,3.9746814,3.4632049,2.951728,2.436347,2.35045,2.260649,2.174752,2.0888553,1.999054,1.6125181,1.2259823,0.8355421,0.44900626,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.23816854,0.41386664,0.58566034,0.76135844,0.93705654,1.4875772,2.0380979,2.5886188,3.1391394,3.6857557,3.2992198,2.912684,2.5261483,2.135708,1.7491722,1.6632754,1.5734742,1.4875772,1.4016805,1.3118792,1.1127546,0.9136301,0.7106012,0.5114767,0.31235218,0.27330816,0.23816854,0.19912452,0.1639849,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.44900626,0.58566034,0.7262188,0.8628729,0.999527,1.4875772,1.9756275,2.463678,2.951728,3.435874,3.8380275,4.2362766,4.6384296,5.036679,5.4388323,6.239235,7.0357327,7.8361354,8.636538,9.43694,8.601398,7.7619514,6.9264097,6.086963,5.251421,5.4856853,5.7238536,5.9620223,6.2001905,6.4383593,5.911265,5.388075,4.860981,4.337791,3.8106966,3.213323,2.612045,2.0107672,1.4133936,0.81211567,0.698888,0.58566034,0.47633708,0.3631094,0.24988174,0.22645533,0.19912452,0.1756981,0.14836729,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.1639849,0.19912452,0.23816854,0.27330816,0.31235218,0.3240654,0.3357786,0.3513962,0.3631094,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.3357786,0.30063897,0.26159495,0.22645533,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.28892577,0.38653582,0.48805028,0.58566034,0.6871748,0.92534333,1.1635119,1.4016805,1.6359446,1.8741131,2.1864653,2.4988174,2.8111696,3.1235218,3.435874,3.951255,4.462732,4.9742084,5.4856853,6.001066,5.4856853,4.9742084,4.462732,3.951255,3.435874,3.7989833,4.1620927,4.5252023,4.8883114,5.251421,5.1889505,5.12648,5.0640097,5.001539,4.939069,4.173806,3.4124475,2.6510892,1.8858263,1.1244678,1.0112402,0.9019169,0.78868926,0.6754616,0.5622339,0.5114767,0.46071947,0.41386664,0.3631094,0.31235218,0.3631094,0.41386664,0.46071947,0.5114767,0.5622339,0.7106012,0.8628729,1.0112402,1.1635119,1.3118792,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.015617609,0.015617609,0.019522011,0.023426414,0.023426414,0.07027924,0.113227665,0.16008049,0.20693332,0.24988174,0.3240654,0.39824903,0.47633708,0.5505207,0.62470436,1.0541886,1.4797685,1.9092526,2.3348327,2.7643168,2.8580225,2.951728,3.049338,3.1430438,3.2367494,3.0259118,2.8189783,2.6081407,2.397303,2.1864653,2.330928,2.4714866,2.6159496,2.7565079,2.900971,3.3812122,3.8614538,4.3416953,4.8219366,5.298274,4.9468775,4.591577,4.2362766,3.8809757,3.5256753,3.4007344,3.279698,3.1586614,3.0337205,2.912684,2.631567,2.3465457,2.0654287,1.7843118,1.4992905,1.2181735,0.94096094,0.659844,0.37872702,0.10151446,0.31625658,0.5349031,0.75354964,0.96829176,1.1869383,1.5656652,1.9482968,2.3270237,2.7057507,3.0883822,2.8189783,2.5456703,2.2762666,2.0068626,1.737459,1.6359446,1.5383345,1.43682,1.33921,1.2376955,1.1010414,0.96438736,0.8238289,0.6871748,0.5505207,0.46852827,0.39044023,0.30844778,0.23035973,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05466163,0.10932326,0.1639849,0.21864653,0.27330816,0.39044023,0.5036679,0.62079996,0.7340276,0.8511597,1.3938715,1.9404879,2.4831998,3.0298162,3.5764325,3.978586,4.380739,4.7828927,5.185046,5.5871997,6.3134184,7.043542,7.7697606,8.495979,9.226103,8.699008,8.171914,7.6409154,7.113821,6.5867267,6.6413884,6.6921453,6.746807,6.7975645,6.8483214,6.1572423,5.466163,4.7711797,4.0801005,3.3890212,2.8814487,2.3738766,1.8663043,1.358732,0.8511597,0.7262188,0.60127795,0.47633708,0.3513962,0.22645533,0.20693332,0.1835069,0.1639849,0.14446288,0.12494087,0.12884527,0.12884527,0.13274968,0.13665408,0.13665408,0.1678893,0.19912452,0.22645533,0.25769055,0.28892577,0.30063897,0.31235218,0.3240654,0.3357786,0.3513962,0.3513962,0.3513962,0.3513962,0.3513962,0.3513962,0.3318742,0.31625658,0.29673457,0.28111696,0.26159495,0.26159495,0.25769055,0.25378615,0.25378615,0.24988174,0.3513962,0.44900626,0.5505207,0.6481308,0.74964523,0.93705654,1.1244678,1.3118792,1.4992905,1.6867018,2.0341935,2.3816853,2.7291772,3.076669,3.4241607,3.8692627,4.31046,4.7516575,5.196759,5.6379566,5.2943697,4.950782,4.6110992,4.267512,3.9239242,4.2362766,4.548629,4.860981,5.173333,5.4856853,5.5442514,5.5989127,5.6535745,5.708236,5.7628975,4.845363,3.9278288,3.0102942,2.0927596,1.175225,1.0932326,1.0151446,0.93315214,0.8550641,0.77307165,0.7223144,0.6715572,0.61689556,0.5661383,0.5114767,0.5427119,0.57394713,0.60127795,0.63251317,0.6637484,0.8316377,0.9956226,1.1635119,1.3314011,1.4992905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.031235218,0.03513962,0.039044023,0.046852827,0.05075723,0.078088045,0.10541886,0.13274968,0.16008049,0.18741131,0.24988174,0.31235218,0.37482262,0.43729305,0.4997635,0.8784905,1.261122,1.639849,2.018576,2.4012074,2.463678,2.5300527,2.5964274,2.6588979,2.7252727,2.592523,2.4597735,2.3270237,2.194274,2.0615244,2.3465457,2.631567,2.9165885,3.2016098,3.4866312,3.9083066,4.3338866,4.755562,5.1772375,5.5989127,5.4036927,5.2045684,5.009348,4.8102236,4.6110992,4.454923,4.298747,4.138666,3.9824903,3.8263142,3.6467118,3.4710135,3.2914112,3.1157131,2.9361105,2.377781,1.8194515,1.2572175,0.698888,0.13665408,0.39824903,0.6559396,0.91753453,1.1791295,1.43682,1.6476578,1.8584955,2.069333,2.2762666,2.4871042,2.3348327,2.182561,2.0302892,1.8780174,1.7257458,1.6125181,1.4992905,1.3860629,1.2767396,1.1635119,1.0893283,1.0112402,0.93705654,0.8628729,0.78868926,0.6637484,0.5427119,0.42167544,0.29673457,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.093705654,0.14055848,0.19131571,0.23816854,0.3318742,0.42167544,0.5153811,0.60908675,0.698888,1.3040704,1.9053483,2.5066261,3.1118085,3.7130866,4.1191444,4.521298,4.927356,5.3334136,5.735567,6.3915067,7.0474463,7.703386,8.359325,9.01136,8.796618,8.577971,8.359325,8.140678,7.9259367,7.793187,7.660437,7.5276875,7.394938,7.262188,6.4032197,5.5442514,4.6813784,3.8224099,2.9634414,2.5456703,2.1318035,1.717937,1.3040704,0.8862993,0.74964523,0.61299115,0.47633708,0.3357786,0.19912452,0.1835069,0.1717937,0.15617609,0.14055848,0.12494087,0.12884527,0.13665408,0.14055848,0.14446288,0.14836729,0.1717937,0.19522011,0.21864653,0.23816854,0.26159495,0.27330816,0.28892577,0.30063897,0.31235218,0.3240654,0.3240654,0.3240654,0.3240654,0.3240654,0.3240654,0.3279698,0.3318742,0.3318742,0.3357786,0.3357786,0.3318742,0.3279698,0.3240654,0.31625658,0.31235218,0.41386664,0.5114767,0.61299115,0.7106012,0.81211567,0.94876975,1.0893283,1.2259823,1.3626363,1.4992905,1.8819219,2.2645533,2.6471848,3.0298162,3.4124475,3.7833657,4.1581883,4.5291066,4.903929,5.2748475,5.1030536,4.93126,4.755562,4.5837684,4.4119744,4.6735697,4.939069,5.2006636,5.462259,5.7238536,5.8956475,6.0713453,6.2431393,6.4149327,6.5867267,5.5130157,4.4432096,3.3694992,2.2957885,1.2259823,1.1791295,1.1283722,1.0815194,1.0346665,0.9878138,0.93315214,0.8784905,0.8238289,0.76916724,0.7106012,0.7223144,0.7340276,0.7418364,0.75354964,0.76135844,0.94876975,1.1322767,1.3157835,1.5031948,1.6867018,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.046852827,0.05075723,0.058566034,0.06637484,0.07418364,0.08589685,0.093705654,0.10541886,0.113227665,0.12494087,0.1756981,0.22645533,0.27330816,0.3240654,0.37482262,0.7066968,1.038571,1.3743496,1.7062237,2.0380979,2.0732377,2.1083772,2.1435168,2.1786566,2.2137961,2.1591344,2.1005683,2.0459068,1.9912452,1.9365835,2.366068,2.7916477,3.2211318,3.6467118,4.0761957,4.4393053,4.806319,5.169429,5.5364423,5.899552,5.860508,5.8214636,5.7785153,5.7394714,5.700427,5.5091114,5.3138914,5.1225758,4.93126,4.73604,4.6657605,4.591577,4.521298,4.447114,4.376835,3.533484,2.6940374,1.8545911,1.0151446,0.1756981,0.47633708,0.78088045,1.0815194,1.3860629,1.6867018,1.7257458,1.7686942,1.8077383,1.8467822,1.8858263,1.8506867,1.8194515,1.7843118,1.7491722,1.7140326,1.5890918,1.4641509,1.33921,1.2142692,1.0893283,1.0737107,1.0619974,1.0502841,1.038571,1.0268579,0.8589685,0.6949836,0.5309987,0.3631094,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.26940376,0.339683,0.40996224,0.48024148,0.5505207,1.2103647,1.8702087,2.5300527,3.1898966,3.8497405,4.2557983,4.6657605,5.0718184,5.481781,5.8878384,6.4695945,7.0513506,7.633106,8.218767,8.800523,8.894228,8.98403,9.077735,9.171441,9.261242,8.944985,8.628729,8.308568,7.9923115,7.676055,6.649197,5.618435,4.591577,3.5647192,2.5378613,2.2137961,1.893635,1.5695697,1.2494087,0.92534333,0.77307165,0.62470436,0.47633708,0.3240654,0.1756981,0.1639849,0.15617609,0.14446288,0.13665408,0.12494087,0.13274968,0.14055848,0.14836729,0.15617609,0.1639849,0.1756981,0.19131571,0.20693332,0.22255093,0.23816854,0.24988174,0.26159495,0.27330816,0.28892577,0.30063897,0.30063897,0.30063897,0.30063897,0.30063897,0.30063897,0.3240654,0.3435874,0.3670138,0.39044023,0.41386664,0.40605783,0.39824903,0.39044023,0.38263142,0.37482262,0.47633708,0.57394713,0.6754616,0.77307165,0.8745861,0.96438736,1.0502841,1.1361811,1.2259823,1.3118792,1.7296503,2.1474214,2.5651922,2.9829633,3.4007344,3.7013733,4.0059166,4.3065557,4.6110992,4.911738,4.911738,4.9078336,4.903929,4.903929,4.900025,5.1108627,5.3256044,5.5364423,5.7511845,5.9620223,6.250948,6.5437784,6.832704,7.1216297,7.4105554,6.184573,4.958591,3.7287042,2.5027218,1.2767396,1.261122,1.2455044,1.2298868,1.2142692,1.1986516,1.1439898,1.0854238,1.0268579,0.96829176,0.9136301,0.9019169,0.8941081,0.8823949,0.8706817,0.8628729,1.0659018,1.2689307,1.4680552,1.6710842,1.8741131,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.058566034,0.07027924,0.078088045,0.08980125,0.10151446,0.093705654,0.08589685,0.078088045,0.07027924,0.062470436,0.10151446,0.13665408,0.1756981,0.21083772,0.24988174,0.5349031,0.8199245,1.1049459,1.3899672,1.6749885,1.678893,1.6867018,1.6906061,1.6945106,1.698415,1.7218413,1.7452679,1.7686942,1.7882162,1.8116426,2.3816853,2.951728,3.521771,4.0918136,4.661856,4.970304,5.278752,5.5832953,5.891743,6.2001905,6.3173227,6.434455,6.551587,6.6687193,6.785851,6.559396,6.3329406,6.1064854,5.8761253,5.64967,5.6809053,5.716045,5.74728,5.7785153,5.813655,4.6930914,3.5725281,2.4519646,1.3314011,0.21083772,0.5583295,0.9019169,1.2494087,1.5929961,1.9365835,1.8077383,1.678893,1.5461433,1.4172981,1.2884527,1.3704453,1.4524376,1.53443,1.6164225,1.698415,1.5617609,1.4251068,1.2884527,1.1517987,1.0112402,1.0619974,1.1127546,1.1635119,1.2142692,1.261122,1.0541886,0.8472553,0.64032197,0.43338865,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.06637484,0.09761006,0.12884527,0.1639849,0.21083772,0.25769055,0.30454338,0.3513962,0.39824903,1.116659,1.8350691,2.5534792,3.2718892,3.9863946,4.396357,4.806319,5.2162814,5.6262436,6.036206,6.547683,7.0591593,7.5667315,8.078208,8.58578,8.991838,9.393991,9.796145,10.198298,10.600452,10.096785,9.593117,9.093353,8.589685,8.086017,6.89127,5.6965227,4.5017757,3.3070288,2.1122816,1.8819219,1.6515622,1.4212024,1.1908426,0.96438736,0.80040246,0.63641757,0.47633708,0.31235218,0.14836729,0.14446288,0.14055848,0.13665408,0.12884527,0.12494087,0.13665408,0.14446288,0.15617609,0.1639849,0.1756981,0.1835069,0.19131571,0.19912452,0.20693332,0.21083772,0.22645533,0.23816854,0.24988174,0.26159495,0.27330816,0.27330816,0.27330816,0.27330816,0.27330816,0.27330816,0.31625658,0.359205,0.40215343,0.44510186,0.48805028,0.47633708,0.46852827,0.45681506,0.44900626,0.43729305,0.5388075,0.63641757,0.737932,0.8394465,0.93705654,0.97610056,1.0112402,1.0502841,1.0893283,1.1244678,1.5773785,2.0302892,2.4831998,2.9361105,3.3890212,3.619381,3.853645,4.084005,4.318269,4.548629,4.716518,4.884407,5.0522966,5.2201858,5.388075,5.548156,5.7121406,5.8761253,6.036206,6.2001905,6.606249,7.016211,7.422269,7.8283267,8.238289,6.8561306,5.473972,4.0918136,2.7057507,1.3235924,1.3431144,1.358732,1.3782539,1.3938715,1.4133936,1.3509232,1.2923572,1.2337911,1.1713207,1.1127546,1.0815194,1.0541886,1.0229534,0.9917182,0.96438736,1.183034,1.4016805,1.6242313,1.8428779,2.0615244,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.3631094,0.60127795,0.8394465,1.0737107,1.3118792,1.2884527,1.261122,1.2376955,1.2142692,1.1869383,1.2884527,1.3860629,1.4875772,1.5890918,1.6867018,2.4012074,3.1118085,3.8263142,4.5369153,5.251421,5.5013027,5.7511845,6.001066,6.250948,6.5008297,6.774138,7.0513506,7.3246584,7.601871,7.8751793,7.6135845,7.348085,7.08649,6.824895,6.5633,6.699954,6.8366084,6.9732623,7.113821,7.250475,5.8487945,4.4510183,3.049338,1.6515622,0.24988174,0.63641757,1.0268579,1.4133936,1.7999294,2.1864653,1.8858263,1.5890918,1.2884527,0.9878138,0.6871748,0.8862993,1.0893283,1.2884527,1.4875772,1.6867018,1.5383345,1.3860629,1.2376955,1.0893283,0.93705654,1.0502841,1.1635119,1.2767396,1.3860629,1.4992905,1.2494087,0.999527,0.74964523,0.4997635,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.1756981,0.19912452,0.22645533,0.24988174,1.0268579,1.7999294,2.5769055,3.349977,4.123049,4.5369153,4.950782,5.3607445,5.774611,6.1884775,6.6257706,7.0630636,7.5003567,7.9376497,8.374943,9.089449,9.80005,10.510651,11.225157,11.935758,11.248583,10.561408,9.874233,9.187058,8.499884,7.137247,5.774611,4.4119744,3.049338,1.6867018,1.5500476,1.4133936,1.2767396,1.1361811,0.999527,0.8238289,0.6481308,0.47633708,0.30063897,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.31235218,0.37482262,0.43729305,0.4997635,0.5622339,0.5505207,0.5388075,0.5231899,0.5114767,0.4997635,0.60127795,0.698888,0.80040246,0.9019169,0.999527,0.9878138,0.97610056,0.96438736,0.94876975,0.93705654,1.4251068,1.9131571,2.4012074,2.8892577,3.3734035,3.5373883,3.7013733,3.8614538,4.025439,4.1894236,4.5252023,4.860981,5.2006636,5.5364423,5.8761253,5.989353,6.098676,6.211904,6.3251314,6.4383593,6.9615493,7.4886436,8.011833,8.538928,9.062118,7.523783,5.985449,4.4510183,2.912684,1.3743496,1.4251068,1.475864,1.5266213,1.5734742,1.6242313,1.5617609,1.4992905,1.43682,1.3743496,1.3118792,1.261122,1.2142692,1.1635119,1.1127546,1.0619974,1.3001659,1.5383345,1.7765031,2.0107672,2.2489357,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.058566034,0.07027924,0.078088045,0.08980125,0.10151446,0.08199245,0.06637484,0.046852827,0.031235218,0.011713207,0.039044023,0.062470436,0.08589685,0.113227665,0.13665408,0.3318742,0.5270943,0.7223144,0.91753453,1.1127546,1.1088502,1.1010414,1.097137,1.0932326,1.0893283,1.1557031,1.2259823,1.2962615,1.3665408,1.43682,2.0732377,2.7057507,3.3421683,3.978586,4.6110992,5.2318993,5.8487945,6.46569,7.082586,7.699481,7.621393,7.5394006,7.461313,7.37932,7.3012323,7.1177254,6.9342184,6.7507114,6.571109,6.387602,6.5359693,6.6843367,6.8287997,6.9771667,7.125534,5.9542136,4.786797,3.6154766,2.4441557,1.2767396,1.4446288,1.6164225,1.7843118,1.9561055,2.1239948,1.8663043,1.6047094,1.3431144,1.0854238,0.8238289,1.1088502,1.3899672,1.6710842,1.9561055,2.2372224,1.9522011,1.6671798,1.3821584,1.097137,0.81211567,0.9097257,1.0073358,1.1049459,1.2025559,1.3001659,1.1049459,0.9097257,0.7145056,0.5192855,0.3240654,0.26940376,0.21474212,0.16008049,0.10541886,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.12494087,0.14836729,0.1756981,0.19912452,0.22645533,0.8628729,1.4992905,2.135708,2.77603,3.4124475,3.8380275,4.263607,4.689187,5.1108627,5.5364423,6.329036,7.1216297,7.914223,8.706817,9.499411,9.897659,10.295909,10.694158,11.088503,11.486752,11.174399,10.858143,10.541886,10.22563,9.913278,8.402273,6.89127,5.3841705,3.873167,2.3621633,2.1239948,1.8819219,1.6437533,1.4016805,1.1635119,0.94876975,0.737932,0.5231899,0.31235218,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10932326,0.12103647,0.12884527,0.14055848,0.14836729,0.15227169,0.15617609,0.15617609,0.16008049,0.1639849,0.1756981,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.25378615,0.26940376,0.28502136,0.30063897,0.3474918,0.39434463,0.44119745,0.48805028,0.5388075,0.5349031,0.5309987,0.5309987,0.5270943,0.5231899,0.60127795,0.679366,0.75745404,0.8355421,0.9136301,0.96438736,1.0112402,1.0619974,1.1127546,1.1635119,1.5773785,1.9912452,2.4090161,2.822883,3.2367494,3.474918,3.7130866,3.951255,4.1894236,4.423688,4.814128,5.2006636,5.5871997,5.9737353,6.364176,6.364176,6.364176,6.364176,6.364176,6.364176,6.852226,7.3441806,7.832231,8.324185,8.812236,7.601871,6.387602,5.173333,3.9629683,2.7486992,2.5456703,2.3465457,2.1435168,1.9404879,1.737459,1.7062237,1.678893,1.6476578,1.6164225,1.5890918,1.4836729,1.3821584,1.2806439,1.1791295,1.0737107,1.261122,1.4485333,1.6359446,1.8233559,2.0107672,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.046852827,0.05075723,0.058566034,0.06637484,0.07418364,0.06637484,0.05466163,0.046852827,0.03513962,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.30063897,0.45681506,0.60908675,0.76135844,0.9136301,0.92924774,0.94096094,0.95657855,0.97219616,0.9878138,1.0268579,1.0659018,1.1088502,1.1478943,1.1869383,1.7452679,2.3035975,2.8619268,3.416352,3.9746814,4.958591,5.9464045,6.930314,7.914223,8.898132,8.464745,8.031356,7.5940623,7.1606736,6.7233806,6.621866,6.520352,6.4188375,6.3134184,6.211904,6.36808,6.5281606,6.6843367,6.844417,7.000593,6.0596323,5.1186714,4.181615,3.240654,2.2996929,2.25284,2.2059872,2.1591344,2.1083772,2.0615244,1.8428779,1.6242313,1.4016805,1.183034,0.96438736,1.3274968,1.6906061,2.05762,2.4207294,2.787743,2.366068,1.9482968,1.5266213,1.1088502,0.6871748,0.76916724,0.8511597,0.93315214,1.0190489,1.1010414,0.96048295,0.8199245,0.679366,0.5388075,0.39824903,0.339683,0.28111696,0.21864653,0.16008049,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.10151446,0.12494087,0.14836729,0.1756981,0.19912452,0.698888,1.1986516,1.698415,2.1981785,2.7018464,3.1391394,3.5764325,4.0137253,4.4510183,4.8883114,6.036206,7.1841,8.32809,9.475985,10.6238785,10.705871,10.791768,10.87376,10.955752,11.037745,11.096312,11.150972,11.209538,11.268105,11.326671,9.6673,8.011833,6.3524623,4.6969957,3.0376248,2.6940374,2.3543546,2.0107672,1.6671798,1.3235924,1.0737107,0.8238289,0.57394713,0.3240654,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.08199245,0.08980125,0.09761006,0.10541886,0.113227665,0.11713207,0.12103647,0.12884527,0.13274968,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.19912452,0.23035973,0.26159495,0.28892577,0.32016098,0.3513962,0.38263142,0.41386664,0.44900626,0.48024148,0.5114767,0.5192855,0.5270943,0.5349031,0.5427119,0.5505207,0.60518235,0.659844,0.7145056,0.76916724,0.8238289,0.93705654,1.0502841,1.1635119,1.2767396,1.3860629,1.7296503,2.0732377,2.416825,2.7565079,3.1000953,3.4124475,3.7247996,4.037152,4.349504,4.661856,5.099149,5.5364423,5.9737353,6.4110284,6.8483214,6.7389984,6.6257706,6.5125427,6.3993154,6.2860875,6.7429028,7.195813,7.6526284,8.105539,8.562354,7.676055,6.785851,5.899552,5.0132523,4.126953,3.6701381,3.213323,2.7604125,2.3035975,1.8506867,1.8506867,1.8545911,1.8584955,1.8584955,1.8623998,1.7062237,1.5539521,1.397776,1.2415999,1.0893283,1.2259823,1.3626363,1.4992905,1.6359446,1.7765031,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.031235218,0.03513962,0.039044023,0.046852827,0.05075723,0.046852827,0.046852827,0.042948425,0.039044023,0.039044023,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.27330816,0.38263142,0.49195468,0.60127795,0.7106012,0.74574083,0.78088045,0.8160201,0.8511597,0.8862993,0.8980125,0.9058213,0.91753453,0.92924774,0.93705654,1.4172981,1.8975395,2.377781,2.8580225,3.338264,4.689187,6.044015,7.394938,8.745861,10.100689,9.308095,8.519405,7.7307167,6.9381227,6.1494336,6.126007,6.1064854,6.083059,6.0596323,6.036206,6.2040954,6.3719845,6.5398736,6.707763,6.8756523,6.165051,5.45445,4.743849,4.0332475,3.3265507,3.0610514,2.795552,2.5300527,2.2645533,1.999054,1.8194515,1.639849,1.4602464,1.2806439,1.1010414,1.5461433,1.9951496,2.4441557,2.8892577,3.338264,2.7838387,2.2294137,1.6710842,1.116659,0.5622339,0.62860876,0.698888,0.76526284,0.8316377,0.9019169,0.8160201,0.7301232,0.6442264,0.5583295,0.47633708,0.40996224,0.3435874,0.28111696,0.21474212,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.1756981,0.5388075,0.9019169,1.261122,1.6242313,1.9873407,2.436347,2.8892577,3.338264,3.78727,4.2362766,5.7394714,7.2426662,8.745861,10.249056,11.748346,11.517986,11.283723,11.053363,10.819098,10.588739,11.018223,11.447707,11.877192,12.306676,12.73616,10.932326,9.128492,7.320754,5.5169206,3.7130866,3.2679846,2.822883,2.377781,1.9326792,1.4875772,1.1986516,0.9136301,0.62470436,0.3357786,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05466163,0.058566034,0.06637484,0.07027924,0.07418364,0.08199245,0.08980125,0.09761006,0.10541886,0.113227665,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.21864653,0.26549935,0.30844778,0.3553006,0.39824903,0.41777104,0.43338865,0.45291066,0.46852827,0.48805028,0.5036679,0.5231899,0.5388075,0.5583295,0.57394713,0.60908675,0.64032197,0.6715572,0.7066968,0.737932,0.9136301,1.0893283,1.261122,1.43682,1.6125181,1.8819219,2.1513257,2.4207294,2.6940374,2.9634414,3.349977,3.736513,4.126953,4.513489,4.900025,5.388075,5.8761253,6.364176,6.8483214,7.336372,7.113821,6.8873653,6.66091,6.4383593,6.211904,6.6335793,7.0513506,7.473026,7.890797,8.312472,7.7502384,7.1880045,6.6257706,6.0635366,5.5013027,4.7907014,4.084005,3.377308,2.6706111,1.9639144,1.999054,2.0341935,2.069333,2.1005683,2.135708,1.9287747,1.7218413,1.5149081,1.3079748,1.1010414,1.1869383,1.2767396,1.3626363,1.4485333,1.5383345,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.015617609,0.015617609,0.019522011,0.023426414,0.023426414,0.031235218,0.03513962,0.039044023,0.046852827,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.1756981,0.24207294,0.30844778,0.37872702,0.44510186,0.5114767,0.5661383,0.62079996,0.679366,0.7340276,0.78868926,0.76916724,0.74574083,0.7262188,0.7066968,0.6871748,1.0893283,1.4914817,1.893635,2.2957885,2.7018464,4.4197836,6.141625,7.859562,9.581403,11.29934,10.155351,9.01136,7.8634663,6.719476,5.575486,5.6340523,5.688714,5.74728,5.805846,5.8644123,6.04011,6.2158084,6.395411,6.571109,6.7507114,6.27047,5.7902284,5.309987,4.829746,4.349504,3.8692627,3.3851168,2.900971,2.4207294,1.9365835,1.796025,1.6593709,1.5188124,1.3782539,1.2376955,1.7686942,2.2957885,2.8267872,3.357786,3.8887846,3.1977055,2.5066261,1.815547,1.1283722,0.43729305,0.48805028,0.5427119,0.59346914,0.6481308,0.698888,0.6715572,0.64032197,0.60908675,0.58175594,0.5505207,0.48024148,0.40996224,0.339683,0.26940376,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.37482262,0.60127795,0.8238289,1.0502841,1.2767396,1.737459,2.1981785,2.6628022,3.1235218,3.5881457,5.446641,7.3012323,9.159728,11.018223,12.8767185,12.326198,11.779582,11.232965,10.686349,10.135828,10.940135,11.740538,12.544845,13.349152,14.149553,12.197352,10.2451515,8.292951,6.3407493,4.388548,3.8380275,3.2914112,2.7447948,2.1981785,1.6515622,1.3235924,0.999527,0.6754616,0.3513962,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.027330816,0.031235218,0.031235218,0.03513962,0.039044023,0.046852827,0.058566034,0.06637484,0.078088045,0.08589685,0.10151446,0.113227665,0.12494087,0.13665408,0.14836729,0.21083772,0.26940376,0.3318742,0.39044023,0.44900626,0.45291066,0.45681506,0.45681506,0.46071947,0.46071947,0.48805028,0.5192855,0.5466163,0.57394713,0.60127795,0.60908675,0.62079996,0.62860876,0.64032197,0.6481308,0.8862993,1.1244678,1.3626363,1.6008049,1.8389735,2.0341935,2.233318,2.4285383,2.6276627,2.8267872,3.2875066,3.7482262,4.21285,4.6735697,5.138193,5.6730967,6.211904,6.7507114,7.2856145,7.824422,7.4886436,7.1489606,6.813182,6.473499,6.13772,6.524256,6.9068875,7.2934237,7.676055,8.062591,7.824422,7.5862536,7.348085,7.113821,6.8756523,5.9151692,4.9546866,3.9942036,3.0337205,2.0732377,2.1435168,2.2098918,2.2762666,2.3465457,2.4129205,2.1513257,1.893635,1.6320401,1.3743496,1.1127546,1.1517987,1.1869383,1.2259823,1.261122,1.3001659,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.21083772,0.23816854,0.26159495,0.28892577,0.31235218,0.38653582,0.46071947,0.5388075,0.61299115,0.6871748,0.63641757,0.58566034,0.5388075,0.48805028,0.43729305,0.76135844,1.0893283,1.4133936,1.737459,2.0615244,4.1503797,6.239235,8.324185,10.413041,12.501896,10.998701,9.499411,8.00012,6.5008297,5.001539,5.138193,5.2748475,5.4115014,5.548156,5.688714,5.8761253,6.0635366,6.250948,6.4383593,6.6257706,6.375889,6.126007,5.8761253,5.6262436,5.376362,4.6735697,3.9746814,3.2757936,2.5769055,1.8741131,1.7765031,1.6749885,1.5734742,1.475864,1.3743496,1.9873407,2.6003318,3.213323,3.8263142,4.4393053,3.611572,2.787743,1.9639144,1.1361811,0.31235218,0.3513962,0.38653582,0.42557985,0.46071947,0.4997635,0.5231899,0.5505207,0.57394713,0.60127795,0.62470436,0.5505207,0.47633708,0.39824903,0.3240654,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.21083772,0.30063897,0.38653582,0.47633708,0.5622339,1.038571,1.5110037,1.9873407,2.463678,2.9361105,5.1499066,7.363703,9.573594,11.787391,14.001186,13.138313,12.27544,11.412568,10.549695,9.686822,10.862047,12.037272,13.212498,14.387722,15.562947,13.462379,11.361811,9.261242,7.164578,5.0640097,4.4119744,3.7638438,3.1118085,2.463678,1.8116426,1.4485333,1.0893283,0.7262188,0.3631094,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.19912452,0.27330816,0.3513962,0.42557985,0.4997635,0.48805028,0.47633708,0.46071947,0.44900626,0.43729305,0.47633708,0.5114767,0.5505207,0.58566034,0.62470436,0.61299115,0.60127795,0.58566034,0.57394713,0.5622339,0.8628729,1.1635119,1.4641509,1.7608855,2.0615244,2.1864653,2.3114061,2.436347,2.5612879,2.6862288,3.2250361,3.7638438,4.298747,4.8375545,5.376362,5.9620223,6.551587,7.137247,7.726812,8.312472,7.8634663,7.4105554,6.9615493,6.5125427,6.0635366,6.4110284,6.7624245,7.113821,7.461313,7.812709,7.898606,7.988407,8.074304,8.164105,8.250002,7.0357327,5.825368,4.6110992,3.4007344,2.1864653,2.2879796,2.3855898,2.4871042,2.5886188,2.6862288,2.3738766,2.0615244,1.7491722,1.43682,1.1244678,1.1127546,1.1010414,1.0893283,1.0737107,1.0619974,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19912452,0.39434463,0.59346914,0.78868926,0.9878138,0.78868926,0.59346914,0.39434463,0.19912452,0.0,0.0,0.0,0.0,0.0,0.0,0.042948425,0.08589685,0.12884527,0.1717937,0.21083772,0.1717937,0.12884527,0.08589685,0.042948425,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.093705654,0.10932326,0.12884527,0.14446288,0.1639849,0.19912452,0.23426414,0.26940376,0.30063897,0.3357786,0.37872702,0.42167544,0.46462387,0.5075723,0.5505207,0.5349031,0.5192855,0.5036679,0.48805028,0.47633708,0.96829176,1.4641509,1.9600099,2.455869,2.951728,4.6852827,6.4188375,8.156297,9.889851,11.623405,10.2451515,8.866898,7.4847393,6.1064854,4.7243266,4.939069,5.1499066,5.3607445,5.575486,5.786324,5.9425,6.098676,6.250948,6.407124,6.5633,6.3173227,6.0713453,5.8292727,5.5832953,5.337318,4.6930914,4.0527697,3.408543,2.7682211,2.1239948,2.0107672,1.901444,1.7882162,1.6749885,1.5617609,2.018576,2.4792955,2.9361105,3.3929255,3.8497405,3.174279,2.4988174,1.8233559,1.1517987,0.47633708,0.5192855,0.5661383,0.60908675,0.6559396,0.698888,0.6715572,0.64032197,0.60908675,0.58175594,0.5505207,0.48414588,0.41386664,0.3474918,0.28111696,0.21083772,0.1796025,0.14836729,0.113227665,0.08199245,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.1717937,0.24597734,0.31625658,0.39044023,0.46071947,0.8511597,1.2415999,1.6320401,2.0224805,2.4129205,4.2362766,6.0635366,7.8868923,9.714153,11.537509,10.928422,10.323239,9.714153,9.108971,8.499884,9.6243515,10.748819,11.873287,13.001659,14.126127,12.263727,10.401327,8.538928,6.676528,4.814128,4.154284,3.49444,2.8306916,2.1708477,1.5110037,1.2142692,0.9136301,0.61299115,0.31235218,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.058566034,0.07027924,0.078088045,0.08980125,0.10151446,0.1639849,0.22645533,0.28892577,0.3513962,0.41386664,0.40215343,0.39434463,0.38263142,0.3709182,0.3631094,0.40215343,0.44119745,0.48414588,0.5231899,0.5622339,0.5583295,0.5544251,0.5466163,0.5427119,0.5388075,0.78868926,1.038571,1.2884527,1.5383345,1.7882162,1.9326792,2.077142,2.2216048,2.366068,2.514435,3.0415294,3.5725281,4.1035266,4.630621,5.1616197,6.0518236,6.9381227,7.824422,8.710721,9.600925,8.859089,8.113348,7.3715115,6.629675,5.8878384,6.914696,7.941554,8.968412,9.999174,11.0260315,10.416945,9.803954,9.194867,8.58578,7.9766936,7.141152,6.3056097,5.4700675,4.6345253,3.7989833,3.677947,3.5569105,3.4319696,3.310933,3.1859922,2.8658314,2.5456703,2.2294137,1.9092526,1.5890918,1.5578566,1.5266213,1.4992905,1.4680552,1.43682,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.39434463,0.78868926,1.1869383,1.5812829,1.9756275,1.5812829,1.1869383,0.78868926,0.39434463,0.0,0.0,0.0,0.0,0.0,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.09761006,0.10932326,0.11713207,0.12884527,0.13665408,0.1835069,0.22645533,0.27330816,0.31625658,0.3631094,0.3709182,0.38263142,0.39434463,0.40215343,0.41386664,0.43338865,0.45291066,0.47243267,0.49195468,0.5114767,1.1791295,1.8428779,2.5066261,3.174279,3.8380275,5.2201858,6.602344,7.984503,9.366661,10.748819,9.491602,8.23048,6.969358,5.708236,4.4510183,4.73604,5.024966,5.3138914,5.5989127,5.8878384,6.008875,6.133816,6.2548523,6.375889,6.5008297,6.2587566,6.0205884,5.7785153,5.5403466,5.298274,4.716518,4.1308575,3.5451972,2.959537,2.3738766,2.2489357,2.1239948,1.999054,1.8741131,1.7491722,2.0537157,2.3543546,2.6588979,2.959537,3.2640803,2.736986,2.2137961,1.6867018,1.1635119,0.63641757,0.6910792,0.7418364,0.79649806,0.8472553,0.9019169,0.8160201,0.7301232,0.6442264,0.5583295,0.47633708,0.41386664,0.3553006,0.29673457,0.23426414,0.1756981,0.16008049,0.14446288,0.12884527,0.113227665,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.13274968,0.19131571,0.24597734,0.30454338,0.3631094,0.6676528,0.97219616,1.2767396,1.5812829,1.8858263,3.3265507,4.7633705,6.2001905,7.6370106,9.073831,8.722435,8.371038,8.015738,7.6643414,7.3129454,8.386656,9.464272,10.537982,11.611692,12.689307,11.061172,9.43694,7.812709,6.1884775,4.564246,3.892689,3.2211318,2.5534792,1.8819219,1.2142692,0.97610056,0.737932,0.4997635,0.26159495,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.046852827,0.05075723,0.058566034,0.06637484,0.07418364,0.12494087,0.1756981,0.22645533,0.27330816,0.3240654,0.31625658,0.30844778,0.30063897,0.29673457,0.28892577,0.3318742,0.3709182,0.41386664,0.45681506,0.4997635,0.5036679,0.5036679,0.5075723,0.5114767,0.5114767,0.7106012,0.9136301,1.1127546,1.3118792,1.5110037,1.678893,1.8428779,2.0068626,2.1708477,2.338737,2.8619268,3.3812122,3.9044023,4.4275923,4.950782,6.13772,7.3246584,8.511597,9.698535,10.889378,9.850807,8.81614,7.7814736,6.746807,5.7121406,7.4183645,9.124588,10.826907,12.533132,14.239355,12.93138,11.623405,10.315431,9.007456,7.699481,7.2426662,6.785851,6.329036,5.8683167,5.4115014,5.067914,4.7243266,4.376835,4.0332475,3.6857557,3.3616903,3.0337205,2.7057507,2.377781,2.0498111,2.0029583,1.9561055,1.9092526,1.8584955,1.8116426,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.59346914,1.183034,1.7765031,2.3699722,2.9634414,2.3699722,1.7765031,1.183034,0.59346914,0.0,0.0,0.0,0.0,0.0,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.10932326,0.08199245,0.05466163,0.027330816,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.10151446,0.10541886,0.10932326,0.10932326,0.113227665,0.1678893,0.22255093,0.27721256,0.3318742,0.38653582,0.3631094,0.3435874,0.32016098,0.29673457,0.27330816,0.3318742,0.38653582,0.44119745,0.4958591,0.5505207,1.3860629,2.2216048,3.0532427,3.8887846,4.7243266,5.755089,6.785851,7.816613,8.843472,9.874233,8.734148,7.5940623,6.453977,5.3138914,4.173806,4.5369153,4.900025,5.263134,5.6262436,5.989353,6.0791545,6.168956,6.2587566,6.348558,6.4383593,6.2040954,5.9659266,5.7316628,5.4973984,5.263134,4.73604,4.2089458,3.6818514,3.1508527,2.6237583,2.4871042,2.35045,2.2137961,2.0732377,1.9365835,2.084951,2.233318,2.3816853,2.5261483,2.6745155,2.2996929,1.9248703,1.5500476,1.175225,0.80040246,0.8589685,0.92143893,0.98000497,1.038571,1.1010414,0.96048295,0.8199245,0.679366,0.5388075,0.39824903,0.3474918,0.29673457,0.24207294,0.19131571,0.13665408,0.14055848,0.14055848,0.14446288,0.14836729,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.093705654,0.13665408,0.1756981,0.21864653,0.26159495,0.48414588,0.7027924,0.92143893,1.1439898,1.3626363,2.4129205,3.4632049,4.513489,5.563773,6.6140575,6.5164475,6.4188375,6.321227,6.223617,6.126007,7.1489606,8.175818,9.198771,10.22563,11.248583,9.86252,8.476458,7.08649,5.700427,4.3143644,3.631094,2.951728,2.2723622,1.5929961,0.9136301,0.737932,0.5622339,0.38653582,0.21083772,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.031235218,0.03513962,0.039044023,0.046852827,0.05075723,0.08589685,0.12494087,0.1639849,0.19912452,0.23816854,0.23426414,0.22645533,0.22255093,0.21864653,0.21083772,0.25769055,0.30063897,0.3474918,0.39434463,0.43729305,0.44900626,0.45681506,0.46852827,0.47633708,0.48805028,0.63641757,0.78868926,0.93705654,1.0893283,1.2376955,1.4212024,1.6086137,1.7921207,1.9756275,2.1630387,2.67842,3.193801,3.7091823,4.220659,4.73604,6.223617,7.7111945,9.198771,10.686349,12.173926,10.84643,9.518932,8.191436,6.8639393,5.5364423,7.9220324,10.303718,12.685403,15.067088,17.448774,15.445815,13.438952,11.435994,9.4291315,7.426173,7.3441806,7.266093,7.1841,7.1060123,7.0240197,6.4578815,5.891743,5.3217,4.755562,4.1894236,3.853645,3.5178664,3.182088,2.8463092,2.514435,2.4480603,2.3816853,2.3192148,2.25284,2.1864653,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.78868926,1.5812829,2.3699722,3.1586614,3.951255,3.1586614,2.3699722,1.5812829,0.78868926,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.10932326,0.10151446,0.09761006,0.093705654,0.08589685,0.15227169,0.21864653,0.28111696,0.3474918,0.41386664,0.359205,0.30063897,0.24597734,0.19131571,0.13665408,0.22645533,0.31625658,0.40605783,0.4958591,0.58566034,1.5929961,2.5964274,3.6037633,4.607195,5.610626,6.289992,6.969358,7.6448197,8.324185,8.999647,7.9805984,6.9615493,5.938596,4.919547,3.900498,4.337791,4.775084,5.212377,5.64967,6.086963,6.1455293,6.2040954,6.2587566,6.3173227,6.375889,6.1455293,5.9151692,5.6848097,5.45445,5.22409,4.755562,4.283129,3.814601,3.3460727,2.87364,2.7252727,2.5769055,2.4246337,2.2762666,2.1239948,2.1161861,2.1083772,2.1005683,2.096664,2.0888553,1.8623998,1.6359446,1.4133936,1.1869383,0.96438736,1.0307622,1.097137,1.1635119,1.2337911,1.3001659,1.1049459,0.9097257,0.7145056,0.5192855,0.3240654,0.28111696,0.23426414,0.19131571,0.14446288,0.10151446,0.12103647,0.14055848,0.16008049,0.1796025,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.05075723,0.078088045,0.10932326,0.13665408,0.1639849,0.29673457,0.43338865,0.5661383,0.7027924,0.8355421,1.4992905,2.1630387,2.8267872,3.4866312,4.1503797,4.3065557,4.466636,4.6228123,4.7789884,4.939069,5.911265,6.8873653,7.8634663,8.835662,9.811763,8.663869,7.5120697,6.364176,5.212377,4.0605783,3.3734035,2.6823244,1.9912452,1.3040704,0.61299115,0.4997635,0.38653582,0.27330816,0.1639849,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.015617609,0.015617609,0.019522011,0.023426414,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.14836729,0.14446288,0.14055848,0.14055848,0.13665408,0.1835069,0.23426414,0.28111696,0.3279698,0.37482262,0.39434463,0.40996224,0.42557985,0.44510186,0.46071947,0.5622339,0.6637484,0.76135844,0.8628729,0.96438736,1.1674163,1.3743496,1.5773785,1.7843118,1.9873407,2.494913,3.0024853,3.5100577,4.01763,4.5252023,6.3134184,8.101635,9.885946,11.674163,13.462379,11.842052,10.221725,8.601398,6.9810715,5.3607445,8.421796,11.482847,14.543899,17.601046,20.662096,17.96025,15.258404,12.556558,9.850807,7.1489606,7.445695,7.746334,8.043069,8.339804,8.636538,7.8478484,7.0591593,6.266566,5.477876,4.689187,4.3455997,4.0020123,3.6584249,3.3187418,2.9751544,2.893162,2.8111696,2.7291772,2.6432803,2.5612879,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.9878138,1.9756275,2.9634414,3.951255,4.939069,3.951255,2.9634414,1.9756275,0.9878138,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.13665408,0.21083772,0.28892577,0.3631094,0.43729305,0.3513962,0.26159495,0.1756981,0.08589685,0.0,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,1.7999294,2.9751544,4.1503797,5.3256044,6.5008297,6.824895,7.1489606,7.47693,7.800996,8.125061,7.223144,6.3251314,5.423215,4.5252023,3.6232853,4.138666,4.650143,5.1616197,5.6730967,6.1884775,6.211904,6.239235,6.262661,6.2860875,6.3134184,6.086963,5.8644123,5.6379566,5.4115014,5.1889505,4.775084,4.3612175,3.951255,3.5373883,3.1235218,2.9634414,2.7994564,2.639376,2.475391,2.3114061,2.1513257,1.9873407,1.8233559,1.6632754,1.4992905,1.4251068,1.3509232,1.2767396,1.1986516,1.1244678,1.1986516,1.2767396,1.3509232,1.4251068,1.4992905,1.2494087,0.999527,0.74964523,0.4997635,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,0.10151446,0.13665408,0.1756981,0.21083772,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.113227665,0.1639849,0.21083772,0.26159495,0.31235218,0.58566034,0.8628729,1.1361811,1.4133936,1.6867018,2.1005683,2.514435,2.9243972,3.338264,3.7482262,4.6735697,5.5989127,6.524256,7.4495993,8.374943,7.461313,6.551587,5.6379566,4.7243266,3.8106966,3.1118085,2.4129205,1.7140326,1.0112402,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.113227665,0.1639849,0.21083772,0.26159495,0.31235218,0.3357786,0.3631094,0.38653582,0.41386664,0.43729305,0.48805028,0.5388075,0.58566034,0.63641757,0.6871748,0.9136301,1.1361811,1.3626363,1.5890918,1.8116426,2.3114061,2.8111696,3.310933,3.8106966,4.3143644,6.3993154,8.488171,10.573121,12.661977,14.750832,12.837675,10.924518,9.01136,7.098203,5.1889505,8.925464,12.661977,16.398489,20.138906,23.87542,20.474686,17.073952,13.673217,10.276386,6.8756523,7.551114,8.226576,8.898132,9.573594,10.249056,9.237816,8.226576,7.211431,6.2001905,5.1889505,4.8375545,4.4861584,4.138666,3.78727,3.435874,3.338264,3.2367494,3.1391394,3.0376248,2.9361105,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.78868926,1.5812829,2.3699722,3.1586614,3.951255,3.1586614,2.3699722,1.5812829,0.78868926,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.10932326,0.1717937,0.23035973,0.28892577,0.3513962,0.28111696,0.21083772,0.14055848,0.07027924,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,1.4602464,2.4207294,3.3812122,4.3416953,5.298274,5.5989127,5.899552,6.2001905,6.5008297,6.801469,6.1884775,5.575486,4.9624953,4.349504,3.736513,4.2440853,4.7516575,5.2592297,5.7668023,6.2743745,6.2470436,6.2197127,6.192382,6.165051,6.13772,6.1025805,6.067441,6.0323014,5.997162,5.9620223,5.704332,5.4427366,5.181142,4.9234514,4.661856,4.825841,4.985922,5.1499066,5.3138914,5.473972,4.83365,4.1894236,3.5491016,2.9048753,2.260649,2.1278992,1.9912452,1.8584955,1.7218413,1.5890918,1.6242313,1.6593709,1.6906061,1.7257458,1.7608855,1.4602464,1.1557031,0.8550641,0.5544251,0.24988174,0.24597734,0.24597734,0.24207294,0.23816854,0.23816854,0.25378615,0.27330816,0.28892577,0.30844778,0.3240654,0.30844778,0.29673457,0.28111696,0.26549935,0.24988174,0.23035973,0.21083772,0.19131571,0.1717937,0.14836729,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.08980125,0.12884527,0.1717937,0.21083772,0.24988174,0.46852827,0.6910792,0.9097257,1.1283722,1.3509232,1.698415,2.0498111,2.4012074,2.7486992,3.1000953,3.9434462,4.786797,5.6262436,6.4695945,7.3129454,6.575013,5.8370814,5.099149,4.3612175,3.6232853,3.0024853,2.3816853,1.756981,1.1361811,0.5114767,0.44900626,0.38653582,0.3240654,0.26159495,0.19912452,0.22645533,0.25378615,0.28111696,0.30844778,0.3357786,0.28892577,0.24207294,0.19522011,0.14836729,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.023426414,0.031235218,0.042948425,0.05075723,0.062470436,0.058566034,0.058566034,0.05466163,0.05075723,0.05075723,0.08980125,0.12884527,0.1717937,0.21083772,0.24988174,0.26940376,0.28892577,0.30844778,0.3318742,0.3513962,0.39434463,0.43338865,0.47633708,0.5192855,0.5622339,0.75745404,0.95267415,1.1478943,1.3431144,1.5383345,1.9522011,2.366068,2.7838387,3.1977055,3.611572,5.388075,7.164578,8.937177,10.71368,12.486279,11.623405,10.760532,9.901564,9.0386915,8.175818,11.986515,15.797212,19.604004,23.4147,27.225397,24.355661,21.48983,18.623999,15.754263,12.888432,13.243732,13.599033,13.954333,14.30573,14.661031,12.861101,11.061172,9.261242,7.461313,5.661383,5.395884,5.12648,4.860981,4.591577,4.3260775,4.60329,4.884407,5.165524,5.446641,5.7238536,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.59346914,1.183034,1.7765031,2.3699722,2.9634414,2.3699722,1.7765031,1.183034,0.59346914,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.08199245,0.12884527,0.1717937,0.21864653,0.26159495,0.21083772,0.15617609,0.10541886,0.05075723,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,1.1205635,1.8663043,2.6081407,3.3538816,4.0996222,4.376835,4.650143,4.9234514,5.2006636,5.473972,5.1499066,4.825841,4.5017757,4.173806,3.8497405,4.3534083,4.853172,5.35684,5.860508,6.364176,6.282183,6.2040954,6.1221027,6.044015,5.9620223,6.1181984,6.2743745,6.426646,6.5828223,6.7389984,6.629675,6.524256,6.4149327,6.3056097,6.2001905,6.688241,7.1762915,7.6643414,8.148487,8.636538,7.5159745,6.3915067,5.270943,4.1464753,3.0259118,2.8306916,2.6354716,2.4402514,2.2450314,2.0498111,2.0459068,2.0380979,2.0341935,2.0302892,2.0263848,1.6710842,1.3157835,0.96048295,0.60518235,0.24988174,0.28111696,0.31625658,0.3474918,0.37872702,0.41386664,0.40996224,0.40605783,0.40605783,0.40215343,0.39824903,0.42167544,0.44119745,0.46071947,0.48024148,0.4997635,0.46071947,0.42167544,0.37872702,0.339683,0.30063897,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.06637484,0.09761006,0.12884527,0.15617609,0.18741131,0.3513962,0.5192855,0.6832704,0.8472553,1.0112402,1.3001659,1.5890918,1.8741131,2.1630387,2.4480603,3.2094188,3.970777,4.728231,5.4895897,6.250948,5.688714,5.12648,4.564246,3.998108,3.435874,2.893162,2.3465457,1.8038338,1.2572175,0.7106012,0.63641757,0.5622339,0.48805028,0.41386664,0.3357786,0.40605783,0.47243267,0.5388075,0.60908675,0.6754616,0.58175594,0.48414588,0.39044023,0.29673457,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.031235218,0.039044023,0.046852827,0.05466163,0.062470436,0.058566034,0.05075723,0.046852827,0.042948425,0.039044023,0.06637484,0.09761006,0.12884527,0.15617609,0.18741131,0.20302892,0.21864653,0.23426414,0.24597734,0.26159495,0.29673457,0.3318742,0.3670138,0.40215343,0.43729305,0.60127795,0.76916724,0.93315214,1.097137,1.261122,1.5929961,1.9209659,2.25284,2.5808098,2.912684,4.376835,5.8370814,7.3012323,8.761478,10.22563,10.413041,10.600452,10.787864,10.975275,11.162686,15.043662,18.928543,22.809519,26.690495,30.575375,28.240541,25.905708,23.570877,21.236044,18.90121,18.936352,18.97149,19.00663,19.041769,19.07691,16.48829,13.899672,11.311053,8.726339,6.13772,5.9542136,5.7668023,5.5832953,5.395884,5.212377,5.872221,6.532065,7.191909,7.8517528,8.511597,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.39434463,0.78868926,1.1869383,1.5812829,1.9756275,1.5812829,1.1869383,0.78868926,0.39434463,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.046852827,0.039044023,0.03513962,0.031235218,0.023426414,0.05466163,0.08589685,0.113227665,0.14446288,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.78088045,1.3118792,1.8389735,2.3699722,2.900971,3.1508527,3.4007344,3.6506162,3.900498,4.1503797,4.1113358,4.0761957,4.037152,3.998108,3.9629683,4.4588275,4.958591,5.45445,5.9542136,6.4500723,6.3173227,6.184573,6.0518236,5.919074,5.786324,6.133816,6.477403,6.8209906,7.168483,7.5120697,7.558923,7.601871,7.648724,7.6916723,7.7385254,8.550641,9.362757,10.174872,10.986988,11.799104,10.198298,8.59359,6.9927845,5.388075,3.78727,3.533484,3.2757936,3.0220075,2.7682211,2.514435,2.4675822,2.4207294,2.377781,2.330928,2.2879796,1.8819219,1.4719596,1.0659018,0.6559396,0.24988174,0.31625658,0.38653582,0.45291066,0.5192855,0.58566034,0.5661383,0.5427119,0.5192855,0.4958591,0.47633708,0.5309987,0.58566034,0.64032197,0.6949836,0.74964523,0.6910792,0.62860876,0.5700427,0.5114767,0.44900626,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.046852827,0.06637484,0.08589685,0.10541886,0.12494087,0.23426414,0.3435874,0.45681506,0.5661383,0.6754616,0.9019169,1.1244678,1.3509232,1.5734742,1.7999294,2.4792955,3.154757,3.8341231,4.5095844,5.1889505,4.7985106,4.4119744,4.025439,3.638903,3.2484627,2.7838387,2.3153105,1.8467822,1.3782539,0.9136301,0.8238289,0.737932,0.6481308,0.5622339,0.47633708,0.58175594,0.6910792,0.79649806,0.9058213,1.0112402,0.8706817,0.7262188,0.58566034,0.44119745,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.042948425,0.046852827,0.05075723,0.058566034,0.062470436,0.05466163,0.046852827,0.039044023,0.031235218,0.023426414,0.046852827,0.06637484,0.08589685,0.10541886,0.12494087,0.13665408,0.14446288,0.15617609,0.1639849,0.1756981,0.20302892,0.23035973,0.25769055,0.28502136,0.31235218,0.44900626,0.58175594,0.71841,0.8511597,0.9878138,1.2337911,1.475864,1.7218413,1.9678187,2.2137961,3.3616903,4.513489,5.661383,6.813182,7.9610763,9.198771,10.436467,11.674163,12.911859,14.149553,18.104713,22.059874,26.015032,29.970192,33.92535,32.121517,30.321589,28.517754,26.71392,24.91399,24.62897,24.343948,24.058928,23.773905,23.488884,20.111576,16.738173,13.360865,9.987461,6.6140575,6.5086384,6.407124,6.3056097,6.2040954,6.098676,7.141152,8.179723,9.218294,10.260769,11.29934,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19912452,0.39434463,0.59346914,0.78868926,0.9878138,0.78868926,0.59346914,0.39434463,0.19912452,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.019522011,0.015617609,0.015617609,0.011713207,0.027330816,0.042948425,0.058566034,0.07418364,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.44119745,0.75354964,1.0698062,1.3860629,1.698415,1.9248703,2.1513257,2.3738766,2.6003318,2.8267872,3.076669,3.3265507,3.5764325,3.8263142,4.0761957,4.5681505,5.0601053,5.55206,6.044015,6.5359693,6.3524623,6.168956,5.9815445,5.7980375,5.610626,6.1494336,6.6843367,7.2192397,7.7541428,8.289046,8.484266,8.683391,8.878611,9.077735,9.276859,10.413041,11.549222,12.689307,13.825488,14.96167,12.880623,10.795672,8.714626,6.6335793,4.548629,4.2362766,3.9200199,3.6037633,3.2914112,2.9751544,2.8892577,2.803361,2.7213683,2.6354716,2.5495746,2.0888553,1.6281357,1.1713207,0.7106012,0.24988174,0.3513962,0.45681506,0.5583295,0.659844,0.76135844,0.71841,0.679366,0.63641757,0.59346914,0.5505207,0.64032197,0.7301232,0.8199245,0.9097257,0.999527,0.92143893,0.8394465,0.76135844,0.679366,0.60127795,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.023426414,0.031235218,0.042948425,0.05075723,0.062470436,0.11713207,0.1717937,0.22645533,0.28111696,0.3357786,0.4997635,0.6637484,0.8238289,0.9878138,1.1517987,1.7452679,2.338737,2.9361105,3.5295796,4.123049,3.912211,3.7013733,3.4866312,3.2757936,3.0610514,2.6706111,2.2840753,1.893635,1.5031948,1.1127546,1.0112402,0.9136301,0.81211567,0.7106012,0.61299115,0.76135844,0.9058213,1.0541886,1.2025559,1.3509232,1.1596074,0.96829176,0.78088045,0.58956474,0.39824903,0.32016098,0.23816854,0.16008049,0.078088045,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05466163,0.058566034,0.058566034,0.062470436,0.05075723,0.042948425,0.031235218,0.023426414,0.011713207,0.023426414,0.031235218,0.042948425,0.05075723,0.062470436,0.06637484,0.07418364,0.078088045,0.08199245,0.08589685,0.10932326,0.12884527,0.14836729,0.1678893,0.18741131,0.29283017,0.39824903,0.5036679,0.60908675,0.7106012,0.8706817,1.0307622,1.1908426,1.3509232,1.5110037,2.35045,3.1859922,4.025439,4.860981,5.700427,7.988407,10.276386,12.564366,14.848442,17.136421,21.165764,25.191204,29.220547,33.245987,37.27533,36.006397,34.733562,33.46463,32.1957,30.926771,30.321589,29.716406,29.111223,28.50604,27.900858,23.738766,19.57277,15.410676,11.248583,7.08649,7.066968,7.0474463,7.027924,7.008402,6.98888,8.406178,9.82738,11.248583,12.665881,14.087084,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.698888,0.9019169,1.1010414,1.3001659,1.4992905,2.0380979,2.5769055,3.1118085,3.6506162,4.1894236,4.6735697,5.1616197,5.64967,6.13772,6.6257706,6.387602,6.1494336,5.911265,5.6730967,5.4388323,6.1611466,6.8873653,7.6135845,8.335898,9.062118,9.413514,9.761005,10.112402,10.4637985,10.81129,12.27544,13.735687,15.199838,16.663988,18.124235,15.562947,13.001659,10.436467,7.8751793,5.3138914,4.939069,4.564246,4.1894236,3.8106966,3.435874,3.310933,3.1859922,3.0610514,2.9361105,2.8111696,2.2996929,1.7882162,1.2767396,0.76135844,0.24988174,0.38653582,0.5231899,0.6637484,0.80040246,0.93705654,0.8745861,0.81211567,0.74964523,0.6871748,0.62470436,0.74964523,0.8745861,0.999527,1.1244678,1.2494087,1.1517987,1.0502841,0.94876975,0.8511597,0.74964523,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,1.0112402,1.5266213,2.0380979,2.5495746,3.0610514,3.0259118,2.9868677,2.951728,2.912684,2.87364,2.5612879,2.2489357,1.9365835,1.6242313,1.3118792,1.1986516,1.0893283,0.97610056,0.8628729,0.74964523,0.93705654,1.1244678,1.3118792,1.4992905,1.6867018,1.4485333,1.2142692,0.97610056,0.737932,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.13665408,0.21083772,0.28892577,0.3631094,0.43729305,0.5114767,0.58566034,0.6637484,0.737932,0.81211567,1.33921,1.8623998,2.3855898,2.912684,3.435874,6.774138,10.112402,13.450665,16.788929,20.12329,24.226816,28.326439,32.42606,36.525684,40.625305,39.887375,39.14944,38.41151,37.673576,36.935646,36.014206,35.088863,34.16352,33.23818,32.31283,27.362051,22.411268,17.460487,12.513609,7.562827,7.6252975,7.687768,7.7502384,7.812709,7.8751793,9.675109,11.475039,13.274967,15.074897,16.874826,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.015617609,0.015617609,0.019522011,0.023426414,0.023426414,0.023426414,0.019522011,0.015617609,0.015617609,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,0.58175594,0.76135844,0.94096094,1.1205635,1.3001659,1.7843118,2.2684577,2.7565079,3.240654,3.7247996,4.193328,4.661856,5.12648,5.5950084,6.0635366,5.9932575,5.9268827,5.860508,5.794133,5.7238536,6.3056097,6.89127,7.473026,8.054782,8.636538,8.925464,9.21439,9.499411,9.788337,10.073358,11.221252,12.365242,13.509232,14.653222,15.801116,14.215929,12.630741,11.045554,9.460366,7.8751793,7.47693,7.0786815,6.6843367,6.2860875,5.8878384,5.591104,5.2943697,4.9937305,4.6969957,4.4002614,3.8263142,3.2562714,2.6823244,2.1083772,1.5383345,1.4016805,1.2689307,1.1322767,0.9956226,0.8628729,0.79649806,0.7340276,0.6676528,0.60127795,0.5388075,0.62860876,0.7223144,0.8160201,0.9058213,0.999527,0.94486535,0.8902037,0.8355421,0.78088045,0.7262188,0.71841,0.7145056,0.7106012,0.7066968,0.698888,0.58956474,0.48024148,0.3709182,0.26159495,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,0.80821127,1.2181735,1.6281357,2.0380979,2.4480603,2.463678,2.475391,2.4871042,2.4988174,2.514435,2.2216048,1.9287747,1.6359446,1.3431144,1.0502841,0.96438736,0.8745861,0.78868926,0.698888,0.61299115,0.8316377,1.0541886,1.2728351,1.4914817,1.7140326,1.4680552,1.2259823,0.98390937,0.7418364,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.10932326,0.1717937,0.23035973,0.28892577,0.3513962,0.41386664,0.48024148,0.5466163,0.60908675,0.6754616,1.1986516,1.7257458,2.2489357,2.77603,3.2992198,6.3407493,9.382278,12.419904,15.461433,18.499058,22.36832,26.233679,30.102942,33.9683,37.837563,37.80242,37.767284,37.732143,37.697002,37.661865,37.259712,36.85756,36.455402,36.05325,35.651096,31.898966,28.15074,24.39861,20.650383,16.902157,17.10909,17.31993,17.530766,17.741604,17.948538,18.90121,19.853886,20.80656,21.759233,22.711908,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.031235218,0.03513962,0.039044023,0.046852827,0.05075723,0.046852827,0.039044023,0.03513962,0.031235218,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.46071947,0.62079996,0.78088045,0.94096094,1.1010414,1.53443,1.9639144,2.397303,2.8306916,3.2640803,3.7091823,4.1581883,4.60329,5.0522966,5.5013027,5.602817,5.704332,5.805846,5.911265,6.012779,6.453977,6.89127,7.3324676,7.773665,8.210958,8.437413,8.663869,8.886419,9.112875,9.339331,10.163159,10.990892,11.818625,12.6463585,13.4740925,12.86891,12.259823,11.650736,11.045554,10.436467,10.018696,9.597021,9.17925,8.757574,8.335898,7.8673706,7.3988423,6.9264097,6.4578815,5.989353,5.35684,4.7243266,4.0918136,3.4593005,2.8267872,2.416825,2.0107672,1.6008049,1.1947471,0.78868926,0.71841,0.6520352,0.58566034,0.5192855,0.44900626,0.5114767,0.5700427,0.62860876,0.6910792,0.74964523,0.7418364,0.7301232,0.71841,0.7106012,0.698888,0.8160201,0.92924774,1.0463798,1.1596074,1.2767396,1.0815194,0.8862993,0.6910792,0.4958591,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.60908675,0.9136301,1.2220778,1.5305257,1.8389735,1.901444,1.9639144,2.0263848,2.0888553,2.1513257,1.8780174,1.6047094,1.3314011,1.0580931,0.78868926,0.7262188,0.6637484,0.60127795,0.5388075,0.47633708,0.7262188,0.98000497,1.2337911,1.4836729,1.737459,1.4914817,1.2415999,0.9956226,0.74574083,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.08199245,0.12884527,0.1717937,0.21864653,0.26159495,0.31625658,0.3709182,0.42557985,0.48414588,0.5388075,1.0619974,1.5890918,2.1122816,2.639376,3.1625657,5.903456,8.648251,11.389141,14.133936,16.874826,20.509825,24.144823,27.779821,31.41482,35.04982,35.717472,36.385124,37.052776,37.72043,38.388084,38.50912,38.62625,38.747288,38.868324,38.98936,36.435883,33.886307,31.336733,28.787157,26.237583,26.596788,26.95209,27.311295,27.666594,28.025799,28.131218,28.236637,28.338152,28.443571,28.548988,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.046852827,0.05075723,0.058566034,0.06637484,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.339683,0.48024148,0.62079996,0.76135844,0.9019169,1.2806439,1.6593709,2.0380979,2.4207294,2.7994564,3.2289407,3.6545205,4.084005,4.5095844,4.939069,5.2084727,5.481781,5.755089,6.028397,6.3017054,6.5984397,6.8951745,7.191909,7.4886436,7.7892823,7.9493628,8.113348,8.273428,8.437413,8.601398,9.108971,9.620447,10.131924,10.639496,11.150972,11.521891,11.888905,12.259823,12.630741,13.001659,12.556558,12.11536,11.674163,11.229061,10.787864,10.143637,9.503315,8.859089,8.218767,7.57454,6.883461,6.1884775,5.4973984,4.806319,4.1113358,3.4319696,2.7526035,2.0732377,1.3938715,0.7106012,0.6442264,0.57394713,0.5036679,0.43338865,0.3631094,0.39044023,0.41777104,0.44510186,0.47243267,0.4997635,0.5349031,0.5700427,0.60518235,0.64032197,0.6754616,0.9097257,1.1439898,1.3782539,1.6164225,1.8506867,1.5695697,1.2884527,1.0112402,0.7301232,0.44900626,0.359205,0.26940376,0.1796025,0.08980125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.40605783,0.60908675,0.8160201,1.0190489,1.2259823,1.33921,1.4485333,1.5617609,1.6749885,1.7882162,1.53443,1.2806439,1.0307622,0.77697605,0.5231899,0.48805028,0.44900626,0.41386664,0.37482262,0.3357786,0.62079996,0.9058213,1.1908426,1.475864,1.7608855,1.5110037,1.2572175,1.0034313,0.75354964,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.05466163,0.08589685,0.113227665,0.14446288,0.1756981,0.21864653,0.26549935,0.30844778,0.3553006,0.39824903,0.92534333,1.4485333,1.9756275,2.4988174,3.0259118,5.4700675,7.914223,10.358379,12.806439,15.250595,18.651329,22.05597,25.456703,28.861341,32.262077,33.632523,35.002968,36.373413,37.74386,39.114304,39.754623,40.39885,41.039173,41.6834,42.32372,40.9767,39.62578,38.274857,36.92393,35.57301,36.08058,36.584248,37.09182,37.59549,38.099155,37.357323,36.615486,35.87365,35.131813,34.38607,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.058566034,0.07027924,0.078088045,0.08980125,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.21864653,0.339683,0.46071947,0.58175594,0.698888,1.0268579,1.3548276,1.6827974,2.0107672,2.338737,2.7447948,3.1508527,3.5608149,3.9668727,4.376835,4.8180323,5.2592297,5.704332,6.1455293,6.5867267,6.7429028,6.899079,7.0513506,7.2075267,7.363703,7.461313,7.562827,7.6643414,7.7619514,7.8634663,8.054782,8.246098,8.441318,8.632633,8.823949,10.170968,11.521891,12.86891,14.215929,15.562947,15.098324,14.633699,14.169076,13.704452,13.235924,12.423808,11.607788,10.791768,9.975748,9.163632,8.410083,7.656533,6.9068875,6.153338,5.3997884,4.447114,3.49444,2.541766,1.5890918,0.63641757,0.5661383,0.49195468,0.42167544,0.3474918,0.27330816,0.26940376,0.26549935,0.26159495,0.25378615,0.24988174,0.3318742,0.40996224,0.48805028,0.5700427,0.6481308,1.0034313,1.358732,1.7140326,2.069333,2.4246337,2.0615244,1.6945106,1.3314011,0.96438736,0.60127795,0.48024148,0.359205,0.23816854,0.12103647,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.20302892,0.30454338,0.40605783,0.5114767,0.61299115,0.77307165,0.93705654,1.1010414,1.261122,1.4251068,1.1908426,0.96048295,0.7262188,0.4958591,0.26159495,0.24988174,0.23816854,0.22645533,0.21083772,0.19912452,0.5192855,0.8355421,1.1517987,1.4680552,1.7882162,1.5305257,1.2728351,1.0151446,0.75745404,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.027330816,0.042948425,0.058566034,0.07418364,0.08589685,0.12103647,0.15617609,0.19131571,0.22645533,0.26159495,0.78868926,1.3118792,1.8389735,2.3621633,2.8892577,5.036679,7.1841,9.331521,11.478943,13.626364,16.796738,19.967113,23.133583,26.303959,29.474333,31.54757,33.620808,35.694046,37.76338,39.836617,41.004032,42.167545,43.331055,44.498474,45.661983,45.51362,45.361347,45.21298,45.060707,44.91234,45.564373,46.216408,46.868446,47.524384,48.17642,46.583424,44.99433,43.40524,41.816147,40.223152,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.77307165,1.0502841,1.3235924,1.6008049,1.8741131,2.260649,2.6510892,3.0376248,3.4241607,3.8106966,4.423688,5.036679,5.64967,6.262661,6.8756523,6.8873653,6.899079,6.910792,6.9264097,6.9381227,6.9732623,7.012306,7.0513506,7.08649,7.125534,7.000593,6.8756523,6.7507114,6.6257706,6.5008297,8.823949,11.150972,13.4740925,15.801116,18.124235,17.636185,17.148134,16.663988,16.175938,15.687888,14.700074,13.712261,12.724447,11.736633,10.748819,9.936704,9.124588,8.312472,7.5003567,6.688241,5.462259,4.2362766,3.0141985,1.7882162,0.5622339,0.48805028,0.41386664,0.3357786,0.26159495,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,1.1010414,1.5734742,2.0498111,2.5261483,2.998581,2.5495746,2.1005683,1.6515622,1.1986516,0.74964523,0.60127795,0.44900626,0.30063897,0.14836729,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21083772,0.42557985,0.63641757,0.8511597,1.0619974,0.8511597,0.63641757,0.42557985,0.21083772,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.41386664,0.76135844,1.1127546,1.4641509,1.8116426,1.5500476,1.2884527,1.0268579,0.76135844,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.6481308,1.175225,1.698415,2.2255092,2.7486992,4.5993857,6.4500723,8.300759,10.151445,11.998228,14.938243,17.874353,20.81437,23.750479,26.68659,29.46262,32.23865,35.010777,37.786804,40.562836,42.24954,43.936237,45.626846,47.313545,49.000248,50.050533,51.100815,52.1511,53.201385,54.25167,55.04817,55.84857,56.64897,57.449375,58.24978,55.81343,53.37318,50.936832,48.500484,46.064137,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.015617609,0.015617609,0.019522011,0.023426414,0.023426414,0.03513962,0.046852827,0.05466163,0.06637484,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.027330816,0.042948425,0.058566034,0.07418364,0.08589685,0.08199245,0.078088045,0.07418364,0.06637484,0.062470436,0.058566034,0.058566034,0.05466163,0.05075723,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.023426414,0.031235218,0.042948425,0.05075723,0.062470436,0.078088045,0.093705654,0.10932326,0.12103647,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.19912452,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.06637484,0.05466163,0.046852827,0.03513962,0.023426414,0.031235218,0.03513962,0.039044023,0.046852827,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.058566034,0.07027924,0.078088045,0.08980125,0.10151446,0.093705654,0.08589685,0.078088045,0.07027924,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,0.62860876,0.8589685,1.0893283,1.319688,1.5500476,1.9326792,2.3153105,2.697942,3.0805733,3.4632049,3.9356375,4.40807,4.8805027,5.3529353,5.825368,5.786324,5.743376,5.704332,5.6652875,5.6262436,5.8683167,6.1103897,6.3524623,6.5945354,6.8366084,7.016211,7.195813,7.37932,7.558923,7.7385254,9.546264,11.354002,13.16174,14.965574,16.773312,16.48829,16.20327,15.918248,15.633226,15.348206,14.739119,14.130032,13.520945,12.911859,12.298867,11.420377,10.541886,9.659492,8.781001,7.898606,6.7780423,5.661383,4.5408196,3.4202564,2.2996929,2.1513257,1.999054,1.8506867,1.698415,1.5500476,1.3821584,1.2142692,1.0463798,0.8784905,0.7106012,0.6715572,0.62860876,0.58566034,0.5427119,0.4997635,0.8823949,1.2650263,1.6476578,2.0302892,2.4129205,2.084951,1.756981,1.4290112,1.1010414,0.77307165,0.6559396,0.5349031,0.41386664,0.29673457,0.1756981,0.14446288,0.113227665,0.08589685,0.05466163,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12103647,0.24597734,0.3670138,0.49195468,0.61299115,0.49195468,0.3670138,0.24597734,0.12103647,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1717937,0.3435874,0.5192855,0.6910792,0.8628729,0.7027924,0.5427119,0.38263142,0.22255093,0.062470436,0.06637484,0.07418364,0.078088045,0.08199245,0.08589685,0.359205,0.63251317,0.9058213,1.1791295,1.4485333,1.2415999,1.0307622,0.8199245,0.60908675,0.39824903,0.32016098,0.23816854,0.16008049,0.078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.5192855,0.94096094,1.358732,1.7804074,2.1981785,3.6857557,5.169429,6.6531014,8.140678,9.6243515,12.201257,14.774258,17.351164,19.924164,22.50107,24.863234,27.229301,29.59537,31.961437,34.3236,36.650623,38.981552,41.308575,43.6356,45.962624,46.688843,47.418964,48.145184,48.871403,49.601524,50.355076,51.108627,51.86608,52.61963,53.37318,50.710377,48.04367,45.380867,42.71416,40.051357,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.031235218,0.03513962,0.039044023,0.046852827,0.05075723,0.058566034,0.06637484,0.07418364,0.078088045,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.042948425,0.058566034,0.078088045,0.093705654,0.113227665,0.10151446,0.093705654,0.08199245,0.07418364,0.062470436,0.058566034,0.05075723,0.046852827,0.042948425,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.046852827,0.06637484,0.08589685,0.10541886,0.12494087,0.15617609,0.1835069,0.21474212,0.24597734,0.27330816,0.30063897,0.3240654,0.3513962,0.37482262,0.39824903,0.37482262,0.3513962,0.3240654,0.30063897,0.27330816,0.23816854,0.19912452,0.1639849,0.12494087,0.08589685,0.078088045,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.046852827,0.042948425,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.046852827,0.05075723,0.058566034,0.06637484,0.07418364,0.07418364,0.07027924,0.06637484,0.06637484,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.48414588,0.6715572,0.8550641,1.038571,1.2259823,1.6008049,1.979532,2.358259,2.7330816,3.1118085,3.4436827,3.775557,4.1113358,4.4432096,4.775084,4.6813784,4.591577,4.4978714,4.4041657,4.3143644,4.759466,5.2084727,5.6535745,6.1025805,6.551587,7.0357327,7.519879,8.0040245,8.488171,8.976221,10.264673,11.553126,12.845484,14.133936,15.426293,15.344301,15.258404,15.176412,15.0944195,15.012426,14.778163,14.547803,14.313539,14.0831785,13.848915,12.90405,11.955279,11.00651,10.061645,9.112875,8.097731,7.082586,6.067441,5.0522966,4.037152,3.8106966,3.5881457,3.3616903,3.1391394,2.912684,2.6159496,2.3192148,2.018576,1.7218413,1.4251068,1.2142692,1.0034313,0.79649806,0.58566034,0.37482262,0.6637484,0.95657855,1.2455044,1.53443,1.8233559,1.620327,1.4133936,1.2103647,1.0034313,0.80040246,0.7106012,0.62079996,0.5309987,0.44119745,0.3513962,0.28892577,0.23035973,0.1717937,0.10932326,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24597734,0.48805028,0.7340276,0.98000497,1.2259823,0.98000497,0.7340276,0.48805028,0.24597734,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13274968,0.26549935,0.39824903,0.5309987,0.6637484,0.5544251,0.44900626,0.339683,0.23426414,0.12494087,0.12103647,0.12103647,0.11713207,0.113227665,0.113227665,0.30844778,0.5036679,0.698888,0.8941081,1.0893283,0.92924774,0.77307165,0.61689556,0.45681506,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.39044023,0.7066968,1.0190489,1.3353056,1.6515622,2.7682211,3.8887846,5.009348,6.1299114,7.250475,9.464272,11.674163,13.887959,16.101755,18.311647,20.267752,22.223858,24.17606,26.132164,28.08827,31.055616,34.02296,36.990307,39.957653,42.925,43.331055,43.73321,44.139267,44.545326,44.95138,45.65808,46.368683,47.07928,47.789883,48.500484,45.607323,42.71416,39.821,36.93174,34.038578,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.046852827,0.05075723,0.058566034,0.06637484,0.07418364,0.078088045,0.08589685,0.08980125,0.093705654,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.058566034,0.078088045,0.09761006,0.11713207,0.13665408,0.12103647,0.10932326,0.093705654,0.078088045,0.062470436,0.05466163,0.046852827,0.039044023,0.031235218,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.08980125,0.13665408,0.1796025,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.06637484,0.09761006,0.12884527,0.15617609,0.18741131,0.23426414,0.27721256,0.3240654,0.3670138,0.41386664,0.44900626,0.48805028,0.5231899,0.5622339,0.60127795,0.5622339,0.5231899,0.48805028,0.44900626,0.41386664,0.3513962,0.28892577,0.22645533,0.1639849,0.10151446,0.093705654,0.08980125,0.08589685,0.078088045,0.07418364,0.06637484,0.05466163,0.046852827,0.03513962,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.031235218,0.03513962,0.039044023,0.046852827,0.05075723,0.05075723,0.05466163,0.058566034,0.058566034,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.339683,0.48024148,0.62079996,0.76135844,0.9019169,1.2728351,1.6437533,2.018576,2.3894942,2.7643168,2.9556324,3.1469483,3.338264,3.533484,3.7247996,3.5803368,3.435874,3.2914112,3.1469483,2.998581,3.6506162,4.3065557,4.958591,5.610626,6.262661,7.0513506,7.843944,8.632633,9.421323,10.213917,10.986988,11.756155,12.529227,13.302299,14.07537,14.196406,14.313539,14.434575,14.555612,14.676648,14.821111,14.965574,15.110037,15.254499,15.398962,14.383818,13.368673,12.353529,11.338385,10.323239,9.413514,8.503788,7.5940623,6.6843367,5.774611,5.473972,5.173333,4.8765984,4.575959,4.2753205,3.8458362,3.4202564,2.9907722,2.5651922,2.135708,1.7608855,1.3821584,1.0034313,0.62860876,0.24988174,0.44900626,0.6442264,0.8433509,1.038571,1.2376955,1.1557031,1.0737107,0.9917182,0.9058213,0.8238289,0.76526284,0.7066968,0.6442264,0.58566034,0.5231899,0.43338865,0.3435874,0.25378615,0.1639849,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3670138,0.7340276,1.1010414,1.4680552,1.8389735,1.4680552,1.1010414,0.7340276,0.3670138,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.093705654,0.1835069,0.27721256,0.3709182,0.46071947,0.40605783,0.3513962,0.29673457,0.24207294,0.18741131,0.1756981,0.1678893,0.15617609,0.14836729,0.13665408,0.25378615,0.3709182,0.49195468,0.60908675,0.7262188,0.62079996,0.5153811,0.40996224,0.30454338,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.26159495,0.46852827,0.679366,0.8902037,1.1010414,1.8545911,2.612045,3.3655949,4.1191444,4.8765984,6.7233806,8.574067,10.424754,12.27544,14.126127,15.668366,17.21451,18.760653,20.306797,21.849035,25.456703,29.064371,32.67204,36.279705,39.887375,39.969364,40.051357,40.13335,40.219246,40.30124,40.96499,41.62874,42.29639,42.960136,43.623886,40.50427,37.38465,34.265034,31.145416,28.025799,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.058566034,0.07027924,0.078088045,0.08980125,0.10151446,0.10151446,0.10541886,0.10932326,0.10932326,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.07418364,0.093705654,0.11713207,0.14055848,0.1639849,0.14055848,0.12103647,0.10151446,0.08199245,0.062470436,0.05075723,0.042948425,0.031235218,0.023426414,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.08980125,0.12884527,0.1717937,0.21083772,0.24988174,0.30844778,0.3709182,0.42948425,0.49195468,0.5505207,0.60127795,0.6481308,0.698888,0.74964523,0.80040246,0.74964523,0.698888,0.6481308,0.60127795,0.5505207,0.46071947,0.37482262,0.28892577,0.19912452,0.113227665,0.10932326,0.10932326,0.10541886,0.10151446,0.10151446,0.08199245,0.06637484,0.046852827,0.031235218,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.015617609,0.015617609,0.019522011,0.023426414,0.023426414,0.031235218,0.039044023,0.046852827,0.05466163,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.19522011,0.28892577,0.38653582,0.48024148,0.57394713,0.94096094,1.3118792,1.678893,2.0459068,2.4129205,2.463678,2.5183394,2.5690966,2.6237583,2.6745155,2.4792955,2.280171,2.0810463,1.8858263,1.6867018,2.5456703,3.4007344,4.2597027,5.1186714,5.9737353,7.0708723,8.164105,9.261242,10.354475,11.4516115,11.705398,11.959184,12.216875,12.470661,12.724447,13.048512,13.368673,13.692739,14.016804,14.336966,14.860155,15.383345,15.906535,16.42582,16.94901,15.867491,14.785972,13.700547,12.619028,11.537509,10.733202,9.928895,9.120684,8.316377,7.5120697,7.137247,6.7624245,6.387602,6.012779,5.6379566,5.0796275,4.521298,3.9668727,3.408543,2.8502135,2.3035975,1.7608855,1.2142692,0.6715572,0.12494087,0.23035973,0.3357786,0.44119745,0.5466163,0.6481308,0.6910792,0.7301232,0.76916724,0.80821127,0.8511597,0.8199245,0.78868926,0.76135844,0.7301232,0.698888,0.58175594,0.46071947,0.339683,0.21864653,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.49195468,0.98000497,1.4719596,1.9600099,2.4480603,1.9600099,1.4719596,0.98000497,0.48805028,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10541886,0.15617609,0.21083772,0.26159495,0.26159495,0.25769055,0.25378615,0.25378615,0.24988174,0.23426414,0.21474212,0.19912452,0.1796025,0.1639849,0.20302892,0.24207294,0.28111696,0.3240654,0.3631094,0.30844778,0.25769055,0.20693332,0.15227169,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.12884527,0.23426414,0.339683,0.44510186,0.5505207,0.94096094,1.3314011,1.7218413,2.1083772,2.4988174,3.9863946,5.473972,6.9615493,8.449126,9.936704,11.072885,12.209065,13.341343,14.477524,15.613705,19.861694,24.109684,28.35377,32.601757,36.849747,36.61158,36.369507,36.13134,35.889267,35.651096,36.271896,36.888794,37.509594,38.130394,38.751194,35.401215,32.05514,28.70907,25.359093,22.01302,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.113227665,0.1639849,0.21083772,0.26159495,0.31235218,0.38653582,0.46071947,0.5388075,0.61299115,0.6871748,0.74964523,0.81211567,0.8745861,0.93705654,0.999527,0.93705654,0.8745861,0.81211567,0.74964523,0.6871748,0.57394713,0.46071947,0.3513962,0.23816854,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.61299115,0.97610056,1.33921,1.698415,2.0615244,1.9756275,1.8858263,1.7999294,1.7140326,1.6242313,1.3743496,1.1244678,0.8745861,0.62470436,0.37482262,1.43682,2.4988174,3.5608149,4.6267166,5.688714,7.08649,8.488171,9.885946,11.287627,12.689307,12.423808,12.162213,11.900618,11.639023,11.373524,11.900618,12.423808,12.950902,13.4740925,14.001186,14.899199,15.801116,16.69913,17.601046,18.499058,17.351164,16.199366,15.051471,13.899672,12.751778,12.0489855,11.350098,10.651209,9.948417,9.249529,8.800523,8.351517,7.898606,7.4495993,7.000593,6.3134184,5.6262436,4.939069,4.251894,3.5608149,2.8502135,2.135708,1.4251068,0.7106012,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.22645533,0.38653582,0.5505207,0.7106012,0.8745861,0.8745861,0.8745861,0.8745861,0.8745861,0.8745861,0.7262188,0.57394713,0.42557985,0.27330816,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.61299115,1.2259823,1.8389735,2.4480603,3.0610514,2.4480603,1.8389735,1.2259823,0.61299115,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.113227665,0.1639849,0.21083772,0.26159495,0.31235218,0.28892577,0.26159495,0.23816854,0.21083772,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,1.2494087,2.3738766,3.4983444,4.6267166,5.7511845,6.473499,7.1997175,7.9259367,8.648251,9.37447,14.262781,19.151093,24.039404,28.923813,33.812122,33.24989,32.687656,32.125423,31.563189,31.000954,31.574902,32.14885,32.7267,33.300648,33.874596,30.29816,26.725634,23.1492,19.576674,16.00024,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05466163,0.058566034,0.058566034,0.062470436,0.07418364,0.08199245,0.093705654,0.10151446,0.113227665,0.12103647,0.13274968,0.14055848,0.15227169,0.1639849,0.14836729,0.13274968,0.11713207,0.10151446,0.08589685,0.10541886,0.12103647,0.14055848,0.15617609,0.1756981,0.14836729,0.12494087,0.10151446,0.07418364,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.30063897,0.38263142,0.46462387,0.5466163,0.62860876,0.7106012,0.76135844,0.80821127,0.8550641,0.9019169,0.94876975,0.8706817,0.79649806,0.71841,0.64032197,0.5622339,0.47243267,0.38263142,0.29283017,0.20302892,0.113227665,0.10932326,0.10932326,0.10541886,0.10151446,0.10151446,0.09761006,0.093705654,0.093705654,0.08980125,0.08589685,0.10932326,0.12884527,0.14836729,0.1678893,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.13665408,0.14446288,0.15617609,0.1639849,0.1756981,0.14836729,0.12103647,0.093705654,0.06637484,0.039044023,0.03513962,0.031235218,0.031235218,0.027330816,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.49195468,0.78478485,1.077615,1.3704453,1.6632754,1.6164225,1.5656652,1.5188124,1.4719596,1.4251068,1.261122,1.0932326,0.92924774,0.76526284,0.60127795,1.5031948,2.4051118,3.3070288,4.2089458,5.1108627,6.27047,7.426173,8.58578,9.741484,10.901091,10.698062,10.495033,10.292005,10.088976,9.885946,10.577025,11.268105,11.959184,12.6463585,13.337439,14.364296,15.387249,16.414106,17.437061,18.463919,17.581524,16.69913,15.816733,14.934339,14.051944,13.314012,12.579984,11.845957,11.111929,10.373997,9.807858,9.24172,8.671678,8.105539,7.5394006,7.08649,6.6335793,6.180669,5.727758,5.2748475,4.396357,3.521771,2.6432803,1.7647898,0.8862993,0.76916724,0.6520352,0.5349031,0.41777104,0.30063897,0.39824903,0.4997635,0.60127795,0.698888,0.80040246,0.78478485,0.76916724,0.75354964,0.7418364,0.7262188,0.61689556,0.5036679,0.39434463,0.28502136,0.1756981,0.15617609,0.14055848,0.12103647,0.10541886,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.49195468,0.98000497,1.4680552,1.9600099,2.4480603,1.9600099,1.4680552,0.98000497,0.48805028,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.08980125,0.12884527,0.1717937,0.21083772,0.24988174,0.23035973,0.21083772,0.19131571,0.1717937,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.999527,1.901444,2.7994564,3.7013733,4.5993857,5.185046,5.7707067,6.356367,6.9381227,7.523783,11.435994,15.344301,19.256512,23.164818,27.073126,26.635832,26.194635,25.753437,25.316145,24.874947,25.441086,26.011127,26.577267,27.143404,27.713448,24.847616,21.981785,19.115953,16.254026,13.388195,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.042948425,0.046852827,0.05075723,0.058566034,0.062470436,0.07027924,0.078088045,0.08589685,0.093705654,0.10151446,0.12103647,0.14055848,0.16008049,0.1796025,0.19912452,0.1835069,0.1639849,0.14836729,0.12884527,0.113227665,0.12103647,0.13274968,0.14055848,0.15227169,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.08980125,0.13665408,0.1796025,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.08589685,0.13665408,0.18741131,0.23816854,0.28892577,0.37872702,0.46852827,0.5583295,0.6481308,0.737932,0.76916724,0.80430686,0.8355421,0.8667773,0.9019169,0.80821127,0.7145056,0.62079996,0.5309987,0.43729305,0.3709182,0.30063897,0.23426414,0.1678893,0.10151446,0.093705654,0.08980125,0.08589685,0.078088045,0.07418364,0.093705654,0.113227665,0.13665408,0.15617609,0.1756981,0.21474212,0.25378615,0.29673457,0.3357786,0.37482262,0.3513962,0.3240654,0.30063897,0.27330816,0.24988174,0.25769055,0.26549935,0.27330816,0.28111696,0.28892577,0.24597734,0.20302892,0.16008049,0.11713207,0.07418364,0.07027924,0.06637484,0.058566034,0.05466163,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.3709182,0.59346914,0.8160201,1.038571,1.261122,1.2533131,1.2494087,1.2415999,1.2337911,1.2259823,1.1439898,1.0659018,0.98390937,0.9058213,0.8238289,1.5656652,2.3114061,3.0532427,3.795079,4.5369153,5.45445,6.36808,7.28171,8.1992445,9.112875,8.968412,8.827853,8.683391,8.542832,8.398369,9.253433,10.108498,10.963562,11.818625,12.67369,13.825488,14.973383,16.125181,17.273075,18.424873,17.811884,17.194988,16.578093,15.965101,15.348206,14.579038,13.809871,13.040704,12.271536,11.498465,10.815194,10.131924,9.444749,8.761478,8.074304,7.8556576,7.6409154,7.422269,7.2036223,6.98888,5.9464045,4.903929,3.8614538,2.8189783,1.7765031,1.5266213,1.2806439,1.0307622,0.78478485,0.5388075,0.57394713,0.61299115,0.6481308,0.6871748,0.7262188,0.6949836,0.6637484,0.63641757,0.60518235,0.57394713,0.5036679,0.43338865,0.3631094,0.29673457,0.22645533,0.21474212,0.20693332,0.19522011,0.1835069,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3670138,0.7340276,1.1010414,1.4680552,1.8389735,1.4680552,1.1010414,0.7340276,0.3670138,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.06637484,0.09761006,0.12884527,0.15617609,0.18741131,0.1717937,0.15617609,0.14055848,0.12884527,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.74964523,1.4251068,2.1005683,2.77603,3.4514916,3.8965936,4.3416953,4.786797,5.2318993,5.6730967,8.609207,11.541413,14.473619,17.405825,20.338032,20.021774,19.701614,19.385357,19.069101,18.74894,19.311174,19.869503,20.431738,20.990067,21.548395,19.393166,17.237936,15.086611,12.93138,10.77615,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.031235218,0.039044023,0.046852827,0.05466163,0.062470436,0.06637484,0.07418364,0.078088045,0.08199245,0.08589685,0.11713207,0.14836729,0.1756981,0.20693332,0.23816854,0.21864653,0.19912452,0.1756981,0.15617609,0.13665408,0.14055848,0.14055848,0.14446288,0.14836729,0.14836729,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.07418364,0.12494087,0.1756981,0.22645533,0.27330816,0.3709182,0.46852827,0.5661383,0.6637484,0.76135844,0.78088045,0.79649806,0.8160201,0.8316377,0.8511597,0.7418364,0.63641757,0.5270943,0.42167544,0.31235218,0.26940376,0.22255093,0.1756981,0.13274968,0.08589685,0.078088045,0.07418364,0.06637484,0.058566034,0.05075723,0.093705654,0.13665408,0.1756981,0.21864653,0.26159495,0.3240654,0.38263142,0.44119745,0.5036679,0.5622339,0.5231899,0.48805028,0.44900626,0.41386664,0.37482262,0.37872702,0.38653582,0.39044023,0.39434463,0.39824903,0.3435874,0.28502136,0.22645533,0.1717937,0.113227665,0.10541886,0.09761006,0.08980125,0.08199245,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.25378615,0.40605783,0.5583295,0.7106012,0.8628729,0.8941081,0.92924774,0.96048295,0.9917182,1.0268579,1.0307622,1.0346665,1.038571,1.0463798,1.0502841,1.6320401,2.2137961,2.7994564,3.3812122,3.9629683,4.6345253,5.3060827,5.9815445,6.6531014,7.3246584,7.2426662,7.1606736,7.0786815,6.996689,6.910792,7.9337454,8.952794,9.971844,10.990892,12.013845,13.286681,14.56342,15.836256,17.112995,18.38583,18.038338,17.690847,17.343355,16.995863,16.64837,15.844065,15.039758,14.235451,13.431144,12.626837,11.82253,11.018223,10.217821,9.413514,8.6131115,8.628729,8.648251,8.663869,8.683391,8.699008,7.492548,6.2860875,5.0757227,3.8692627,2.6628022,2.2840753,1.9092526,1.5305257,1.1517987,0.77307165,0.74964523,0.7262188,0.698888,0.6754616,0.6481308,0.60518235,0.5583295,0.5153811,0.46852827,0.42557985,0.39434463,0.3631094,0.3357786,0.30454338,0.27330816,0.27330816,0.26940376,0.26940376,0.26549935,0.26159495,0.21083772,0.15617609,0.10541886,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24597734,0.48805028,0.7340276,0.98000497,1.2259823,0.98000497,0.7340276,0.48805028,0.24597734,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.046852827,0.06637484,0.08589685,0.10541886,0.12494087,0.113227665,0.10541886,0.093705654,0.08589685,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.4997635,0.94876975,1.4016805,1.8506867,2.2996929,2.6042364,2.9087796,3.213323,3.521771,3.8263142,5.7785153,7.734621,9.690726,11.6468315,13.599033,13.403813,13.208592,13.013372,12.818152,12.626837,13.177358,13.731783,14.282304,14.836729,15.387249,13.94262,12.497992,11.053363,9.608734,8.164105,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.023426414,0.031235218,0.042948425,0.05075723,0.062470436,0.06637484,0.06637484,0.07027924,0.07418364,0.07418364,0.113227665,0.15617609,0.19522011,0.23426414,0.27330816,0.25378615,0.23035973,0.20693332,0.1835069,0.1639849,0.15617609,0.15227169,0.14836729,0.14055848,0.13665408,0.113227665,0.08589685,0.062470436,0.039044023,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.062470436,0.113227665,0.1639849,0.21083772,0.26159495,0.3670138,0.47243267,0.57785153,0.6832704,0.78868926,0.78868926,0.79259366,0.79649806,0.79649806,0.80040246,0.679366,0.5544251,0.43338865,0.30844778,0.18741131,0.1639849,0.14055848,0.12103647,0.09761006,0.07418364,0.06637484,0.05466163,0.046852827,0.03513962,0.023426414,0.08980125,0.15617609,0.21864653,0.28502136,0.3513962,0.42948425,0.5114767,0.58956474,0.6715572,0.74964523,0.698888,0.6481308,0.60127795,0.5505207,0.4997635,0.5036679,0.5036679,0.5075723,0.5114767,0.5114767,0.44119745,0.3670138,0.29673457,0.22255093,0.14836729,0.14055848,0.12884527,0.12103647,0.10932326,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.13274968,0.21474212,0.29673457,0.37872702,0.46071947,0.5349031,0.60908675,0.679366,0.75354964,0.8238289,0.9136301,1.0034313,1.0932326,1.1869383,1.2767396,1.698415,2.1200905,2.541766,2.9634414,3.3890212,3.8185053,4.2479897,4.677474,5.1069584,5.5364423,5.5169206,5.493494,5.4700675,5.446641,5.423215,6.610153,7.793187,8.980125,10.163159,11.350098,12.751778,14.149553,15.551234,16.94901,18.35069,18.268698,18.19061,18.108618,18.030529,17.948538,17.10909,16.269644,15.430198,14.590752,13.751305,12.829865,11.908427,10.990892,10.069453,9.151918,9.4018,9.655587,9.909373,10.159255,10.413041,9.0386915,7.6682463,6.2938967,4.9234514,3.5491016,3.0415294,2.533957,2.0263848,1.5188124,1.0112402,0.92534333,0.8394465,0.74964523,0.6637484,0.57394713,0.5153811,0.45681506,0.39434463,0.3357786,0.27330816,0.28502136,0.29673457,0.30454338,0.31625658,0.3240654,0.3318742,0.3357786,0.339683,0.3435874,0.3513962,0.28111696,0.21083772,0.14055848,0.07027924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12103647,0.24597734,0.3670138,0.48805028,0.61299115,0.48805028,0.3670138,0.24597734,0.12103647,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.023426414,0.031235218,0.042948425,0.05075723,0.062470436,0.058566034,0.05075723,0.046852827,0.042948425,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.24988174,0.47633708,0.698888,0.92534333,1.1517987,1.3157835,1.4797685,1.6437533,1.8116426,1.9756275,2.951728,3.9317331,4.9078336,5.883934,6.8639393,6.7897553,6.715572,6.6452928,6.571109,6.5008297,7.043542,7.590158,8.136774,8.679486,9.226103,8.488171,7.7541428,7.0201154,6.2860875,5.548156,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.113227665,0.1639849,0.21083772,0.26159495,0.31235218,0.28892577,0.26159495,0.23816854,0.21083772,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.3631094,0.47633708,0.58566034,0.698888,0.81211567,0.80040246,0.78868926,0.77307165,0.76135844,0.74964523,0.61299115,0.47633708,0.3357786,0.19912452,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.5388075,0.63641757,0.737932,0.8394465,0.93705654,0.8745861,0.81211567,0.74964523,0.6871748,0.62470436,0.62470436,0.62470436,0.62470436,0.62470436,0.62470436,0.5388075,0.44900626,0.3631094,0.27330816,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.1756981,0.28892577,0.39824903,0.5114767,0.62470436,0.80040246,0.97610056,1.1517987,1.3235924,1.4992905,1.7608855,2.0263848,2.2879796,2.5495746,2.8111696,2.998581,3.1859922,3.3734035,3.5608149,3.7482262,3.78727,3.8263142,3.8614538,3.900498,3.9356375,5.2865605,6.6374836,7.988407,9.339331,10.686349,12.212971,13.735687,15.262308,16.788929,18.311647,18.499058,18.68647,18.87388,19.061293,19.248703,18.374117,17.49953,16.624945,15.750359,14.875772,13.837202,12.798631,11.763964,10.725393,9.686822,10.174872,10.662923,11.150972,11.639023,12.123169,10.588739,9.050405,7.5120697,5.9737353,4.4393053,3.7989833,3.1625657,2.5261483,1.8858263,1.2494087,1.1010414,0.94876975,0.80040246,0.6481308,0.4997635,0.42557985,0.3513962,0.27330816,0.19912452,0.12494087,0.1756981,0.22645533,0.27330816,0.3240654,0.37482262,0.38653582,0.39824903,0.41386664,0.42557985,0.43729305,0.3513962,0.26159495,0.1756981,0.08589685,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.1756981,0.22645533,0.27330816,0.3240654,0.37482262,0.9136301,1.4485333,1.9873407,2.5261483,3.0610514,3.0376248,3.0141985,2.9868677,2.9634414,2.9361105,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.08980125,0.12884527,0.1717937,0.21083772,0.24988174,0.23035973,0.21083772,0.19131571,0.1717937,0.14836729,0.14055848,0.12884527,0.12103647,0.10932326,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.015617609,0.023426414,0.027330816,0.031235218,0.039044023,0.03513962,0.031235218,0.031235218,0.027330816,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.027330816,0.031235218,0.031235218,0.03513962,0.039044023,0.031235218,0.027330816,0.023426414,0.015617609,0.011713207,0.05075723,0.08589685,0.12494087,0.1639849,0.19912452,0.1639849,0.12884527,0.093705654,0.058566034,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.28892577,0.37872702,0.46852827,0.5583295,0.6481308,0.6442264,0.64032197,0.63641757,0.62860876,0.62470436,0.5700427,0.5153811,0.46071947,0.40605783,0.3513962,0.3279698,0.30454338,0.28111696,0.26159495,0.23816854,0.23035973,0.22255093,0.21474212,0.20693332,0.19912452,0.28892577,0.37482262,0.46071947,0.5505207,0.63641757,0.76526284,0.8941081,1.0190489,1.1478943,1.2767396,1.1908426,1.1049459,1.0190489,0.93315214,0.8511597,0.78478485,0.71841,0.6559396,0.58956474,0.5231899,0.44900626,0.37482262,0.30063897,0.22645533,0.14836729,0.14836729,0.14446288,0.14055848,0.14055848,0.13665408,0.10932326,0.08199245,0.05466163,0.027330816,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.20693332,0.30844778,0.40996224,0.5114767,0.42557985,0.3357786,0.24988174,0.1639849,0.07418364,0.16008049,0.24597734,0.3318742,0.41386664,0.4997635,0.64032197,0.78088045,0.92143893,1.0580931,1.1986516,1.4133936,1.6242313,1.8389735,2.0498111,2.260649,2.4285383,2.592523,2.7565079,2.9243972,3.0883822,3.3148375,3.541293,3.7716527,3.998108,4.224563,5.282656,6.3407493,7.3988423,8.456935,9.511124,11.018223,12.521418,14.028518,15.531713,17.03881,17.31993,17.601046,17.886066,18.167183,18.448301,18.057861,17.663515,17.273075,16.87873,16.48829,15.74255,14.996809,14.251068,13.509232,12.763491,12.677594,12.591698,12.5058,12.423808,12.337912,10.8542385,9.37447,7.890797,6.407124,4.9234514,4.267512,3.611572,2.951728,2.2957885,1.6359446,1.4875772,1.33921,1.1869383,1.038571,0.8862993,0.8433509,0.80430686,0.76135844,0.71841,0.6754616,0.6715572,0.6637484,0.659844,0.6559396,0.6481308,0.59346914,0.5388075,0.48414588,0.42948425,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.14055848,0.1835069,0.22645533,0.26940376,0.31235218,0.74964523,1.1869383,1.6242313,2.0615244,2.4988174,2.4792955,2.4597735,2.4402514,2.4207294,2.4012074,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.06637484,0.09761006,0.12884527,0.15617609,0.18741131,0.1717937,0.15617609,0.14055848,0.12884527,0.113227665,0.10541886,0.09761006,0.08980125,0.08199245,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.03513962,0.046852827,0.05466163,0.06637484,0.07418364,0.07027924,0.06637484,0.058566034,0.05466163,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05466163,0.058566034,0.06637484,0.07027924,0.07418364,0.06637484,0.05466163,0.046852827,0.03513962,0.023426414,0.10151446,0.1756981,0.24988174,0.3240654,0.39824903,0.3318742,0.26159495,0.19131571,0.12103647,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.21864653,0.28502136,0.3513962,0.42167544,0.48805028,0.48805028,0.49195468,0.4958591,0.4958591,0.4997635,0.5270943,0.5544251,0.58175594,0.60908675,0.63641757,0.59346914,0.5466163,0.5036679,0.45681506,0.41386664,0.40996224,0.40605783,0.40605783,0.40215343,0.39824903,0.48805028,0.57394713,0.6637484,0.74964523,0.8394465,0.9917182,1.1478943,1.3040704,1.456342,1.6125181,1.5031948,1.397776,1.2884527,1.183034,1.0737107,0.94486535,0.8160201,0.6832704,0.5544251,0.42557985,0.3631094,0.30063897,0.23816854,0.1756981,0.113227665,0.12103647,0.12884527,0.13665408,0.14055848,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.20693332,0.40996224,0.61689556,0.8199245,1.0268579,0.8355421,0.6481308,0.46071947,0.27330816,0.08589685,0.14446288,0.20302892,0.26159495,0.31625658,0.37482262,0.48024148,0.58566034,0.6910792,0.79649806,0.9019169,1.0619974,1.2259823,1.3860629,1.5500476,1.7140326,1.8545911,1.999054,2.1396124,2.2840753,2.4246337,2.8424048,3.260176,3.677947,4.095718,4.513489,5.278752,6.044015,6.8092775,7.570636,8.335898,9.823476,11.307149,12.790822,14.278399,15.762072,16.140799,16.515621,16.894348,17.273075,17.651802,17.741604,17.831406,17.921206,18.011007,18.10081,17.647898,17.194988,16.742077,16.289165,15.836256,15.180316,14.524376,13.864532,13.208592,12.548749,11.123642,9.694631,8.265619,6.8405128,5.4115014,4.73604,4.056674,3.3812122,2.7018464,2.0263848,1.8741131,1.7257458,1.5734742,1.4251068,1.2767396,1.2650263,1.2533131,1.2455044,1.2337911,1.2259823,1.1635119,1.1049459,1.0463798,0.98390937,0.92534333,0.80430686,0.679366,0.5583295,0.43338865,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.10932326,0.14446288,0.1796025,0.21474212,0.24988174,0.58566034,0.92534333,1.261122,1.6008049,1.9365835,1.9209659,1.9092526,1.893635,1.8780174,1.8623998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.046852827,0.06637484,0.08589685,0.10541886,0.12494087,0.113227665,0.10541886,0.093705654,0.08589685,0.07418364,0.07027924,0.06637484,0.058566034,0.05466163,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.44900626,0.359205,0.26940376,0.1796025,0.08980125,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.05075723,0.06637484,0.08199245,0.09761006,0.113227665,0.10541886,0.09761006,0.08980125,0.08199245,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.08199245,0.08980125,0.09761006,0.10541886,0.113227665,0.09761006,0.08199245,0.06637484,0.05075723,0.039044023,0.14836729,0.26159495,0.37482262,0.48805028,0.60127795,0.4958591,0.39044023,0.28502136,0.1796025,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.14446288,0.19131571,0.23426414,0.28111696,0.3240654,0.3357786,0.3435874,0.3553006,0.3631094,0.37482262,0.48414588,0.59346914,0.7066968,0.8160201,0.92534333,0.8589685,0.78868926,0.7223144,0.6559396,0.58566034,0.58956474,0.59346914,0.59346914,0.59737355,0.60127795,0.6871748,0.77307165,0.8628729,0.94876975,1.038571,1.2181735,1.4016805,1.5851873,1.7686942,1.9482968,1.8194515,1.6906061,1.5617609,1.4290112,1.3001659,1.1049459,0.9097257,0.7145056,0.5192855,0.3240654,0.27330816,0.22645533,0.1756981,0.12494087,0.07418364,0.093705654,0.10932326,0.12884527,0.14446288,0.1639849,0.12884527,0.09761006,0.06637484,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.30844778,0.61689556,0.92143893,1.2298868,1.5383345,1.2494087,0.96438736,0.6754616,0.38653582,0.10151446,0.12884527,0.16008049,0.19131571,0.21864653,0.24988174,0.32016098,0.39044023,0.46071947,0.5309987,0.60127795,0.7106012,0.8238289,0.93705654,1.0502841,1.1635119,1.2806439,1.4016805,1.5227169,1.6437533,1.7608855,2.3699722,2.979059,3.5842414,4.193328,4.7985106,5.270943,5.743376,6.2158084,6.688241,7.1606736,8.628729,10.09288,11.557031,13.021181,14.489237,14.96167,15.434102,15.906535,16.378967,16.8514,17.421442,17.99539,18.569338,19.13938,19.713327,19.553246,19.393166,19.233086,19.073006,18.912924,17.683039,16.453152,15.223265,13.993378,12.763491,11.389141,10.018696,8.644346,7.2739015,5.899552,5.2006636,4.50568,3.8067923,3.1118085,2.4129205,2.260649,2.1122816,1.9639144,1.8116426,1.6632754,1.6867018,1.7062237,1.7296503,1.7530766,1.7765031,1.6593709,1.5461433,1.4290112,1.3157835,1.1986516,1.0112402,0.8199245,0.62860876,0.44119745,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.046852827,0.08980125,0.13665408,0.1796025,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.078088045,0.10541886,0.13274968,0.16008049,0.18741131,0.42557985,0.6637484,0.9019169,1.1361811,1.3743496,1.3665408,1.3548276,1.3431144,1.3353056,1.3235924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.023426414,0.031235218,0.042948425,0.05075723,0.062470436,0.058566034,0.05075723,0.046852827,0.042948425,0.039044023,0.03513962,0.031235218,0.031235218,0.027330816,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.60127795,0.48024148,0.359205,0.23816854,0.12103647,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.07027924,0.08980125,0.10932326,0.12884527,0.14836729,0.14055848,0.12884527,0.12103647,0.10932326,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10932326,0.12103647,0.12884527,0.14055848,0.14836729,0.12884527,0.10932326,0.08980125,0.07027924,0.05075723,0.19912452,0.3513962,0.4997635,0.6481308,0.80040246,0.659844,0.5192855,0.37872702,0.23816854,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.07418364,0.093705654,0.11713207,0.14055848,0.1639849,0.1796025,0.19912452,0.21474212,0.23426414,0.24988174,0.44119745,0.63641757,0.8277333,1.0190489,1.2142692,1.1205635,1.0307622,0.94096094,0.8511597,0.76135844,0.76916724,0.77697605,0.78478485,0.79259366,0.80040246,0.8862993,0.97610056,1.0619974,1.1517987,1.2376955,1.4485333,1.6593709,1.8663043,2.077142,2.2879796,2.135708,1.9834363,1.8311646,1.678893,1.5266213,1.2650263,1.0034313,0.74574083,0.48414588,0.22645533,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.06637484,0.093705654,0.12103647,0.14836729,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.40996224,0.8199245,1.2298868,1.639849,2.0498111,1.6632754,1.2767396,0.8862993,0.4997635,0.113227665,0.113227665,0.11713207,0.12103647,0.12103647,0.12494087,0.16008049,0.19522011,0.23035973,0.26549935,0.30063897,0.3631094,0.42557985,0.48805028,0.5505207,0.61299115,0.7106012,0.80821127,0.9058213,1.0034313,1.1010414,1.8975395,2.6940374,3.49444,4.290938,5.087436,5.267039,5.446641,5.6262436,5.805846,5.989353,7.433982,8.878611,10.323239,11.767868,13.212498,13.778636,14.348679,14.914817,15.480955,16.050997,17.105186,18.159374,19.213564,20.271656,21.325846,21.458595,21.591345,21.724094,21.856844,21.98569,20.18576,18.381926,16.578093,14.778163,12.974329,11.6585455,10.338858,9.023073,7.703386,6.387602,5.6691923,4.950782,4.2362766,3.5178664,2.7994564,2.6510892,2.4988174,2.35045,2.1981785,2.0498111,2.1044729,2.1591344,2.2137961,2.2684577,2.3231194,2.15523,1.9834363,1.815547,1.6437533,1.475864,1.2181735,0.96048295,0.7027924,0.44510186,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.046852827,0.06637484,0.08589685,0.10541886,0.12494087,0.26159495,0.39824903,0.5388075,0.6754616,0.81211567,0.80821127,0.80430686,0.79649806,0.79259366,0.78868926,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,0.74964523,0.60127795,0.44900626,0.30063897,0.14836729,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.24988174,0.43729305,0.62470436,0.81211567,0.999527,0.8238289,0.6481308,0.47633708,0.30063897,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.39824903,0.6754616,0.94876975,1.2259823,1.4992905,1.3860629,1.2767396,1.1635119,1.0502841,0.93705654,0.94876975,0.96438736,0.97610056,0.9878138,0.999527,1.0893283,1.175225,1.261122,1.3509232,1.43682,1.6749885,1.9131571,2.1513257,2.3855898,2.6237583,2.4480603,2.2762666,2.1005683,1.9248703,1.7491722,1.4251068,1.1010414,0.77307165,0.44900626,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5114767,1.0268579,1.5383345,2.0498111,2.5612879,2.0732377,1.5890918,1.1010414,0.61299115,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.13665408,0.21083772,0.28892577,0.3631094,0.43729305,1.4251068,2.4129205,3.4007344,4.388548,5.376362,5.263134,5.1499066,5.036679,4.9234514,4.814128,6.239235,7.6643414,9.089449,10.510651,11.935758,12.599506,13.263254,13.923099,14.586847,15.250595,16.788929,18.32336,19.861694,21.400028,22.938364,23.363943,23.785618,24.211199,24.636778,25.062359,22.688482,20.310701,17.936825,15.562947,13.189071,11.924045,10.662923,9.4018,8.136774,6.8756523,6.13772,5.3997884,4.661856,3.9239242,3.1859922,3.0376248,2.8892577,2.736986,2.5886188,2.436347,2.5261483,2.612045,2.7018464,2.787743,2.87364,2.6510892,2.4246337,2.1981785,1.9756275,1.7491722,1.4251068,1.1010414,0.77307165,0.44900626,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.10151446,0.13665408,0.1756981,0.21083772,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.042948425,0.058566034,0.078088045,0.093705654,0.113227665,0.113227665,0.113227665,0.113227665,0.113227665,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.019522011,0.015617609,0.015617609,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.042948425,0.07418364,0.10151446,0.13274968,0.1639849,0.25769055,0.3513962,0.44900626,0.5427119,0.63641757,0.5114767,0.38263142,0.25378615,0.12884527,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.046852827,0.078088045,0.10932326,0.14055848,0.1756981,0.1678893,0.16008049,0.15227169,0.14446288,0.13665408,0.18741131,0.23816854,0.28892577,0.3357786,0.38653582,0.3513962,0.31235218,0.27330816,0.23816854,0.19912452,0.24207294,0.28502136,0.3279698,0.3709182,0.41386664,0.359205,0.30844778,0.25378615,0.20302892,0.14836729,0.12884527,0.10932326,0.08980125,0.07027924,0.05075723,0.19912452,0.3513962,0.4997635,0.6481308,0.80040246,0.6676528,0.5349031,0.40215343,0.26940376,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.19912452,0.61689556,1.0307622,1.4446288,1.8584955,2.2762666,2.2645533,2.2567444,2.2450314,2.233318,2.2255092,1.9912452,1.756981,1.5188124,1.2845483,1.0502841,1.1010414,1.1517987,1.1986516,1.2494087,1.3001659,1.3235924,1.3431144,1.3665408,1.3899672,1.4133936,1.1986516,0.9878138,0.77307165,0.5622339,0.3513962,0.57785153,0.80430686,1.0307622,1.261122,1.4875772,1.5149081,1.542239,1.5695697,1.5969005,1.6242313,1.5070993,1.3899672,1.2728351,1.1557031,1.038571,1.0893283,1.1361811,1.1869383,1.2376955,1.2884527,1.6632754,2.0380979,2.4129205,2.787743,3.1625657,2.9243972,2.6862288,2.4480603,2.2137961,1.9756275,1.6593709,1.33921,1.0229534,0.7066968,0.38653582,0.3474918,0.30844778,0.26940376,0.22645533,0.18741131,0.1796025,0.1717937,0.1639849,0.15617609,0.14836729,0.14446288,0.14055848,0.13665408,0.12884527,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.40996224,0.8199245,1.2298868,1.639849,2.0498111,1.6593709,1.2689307,0.8784905,0.48805028,0.10151446,0.1678893,0.23426414,0.30063897,0.3709182,0.43729305,0.3513962,0.26159495,0.1756981,0.08589685,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.3709182,0.60127795,0.8355421,1.0659018,1.3001659,2.0029583,2.7057507,3.408543,4.1113358,4.814128,4.6969957,4.5837684,4.466636,4.3534083,4.2362766,5.4154058,6.590631,7.7697606,8.94889,10.124115,10.77615,11.424281,12.076316,12.724447,13.376482,15.000713,16.624945,18.249176,19.873407,21.501543,22.434696,23.371752,24.304905,25.24196,26.175114,23.953508,21.735807,19.514202,17.296501,15.074897,13.645885,12.216875,10.783959,9.354948,7.9259367,7.2426662,6.559396,5.8761253,5.196759,4.513489,4.251894,3.9942036,3.7326086,3.4710135,3.213323,3.1391394,3.06886,2.9946766,2.9243972,2.8502135,2.7408905,2.631567,2.5183394,2.4090161,2.2996929,1.9639144,1.6242313,1.2884527,0.94876975,0.61299115,0.5036679,0.39434463,0.28111696,0.1717937,0.062470436,0.08980125,0.11713207,0.14446288,0.1717937,0.19912452,0.27330816,0.3513962,0.42557985,0.4997635,0.57394713,0.47243267,0.3709182,0.26940376,0.1639849,0.062470436,0.06637484,0.07418364,0.078088045,0.08199245,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12884527,0.26159495,0.39044023,0.5192855,0.6481308,0.5192855,0.39044023,0.26159495,0.12884527,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.08980125,0.13665408,0.1796025,0.22645533,0.23035973,0.23426414,0.23816854,0.24597734,0.24988174,0.26159495,0.27330816,0.28892577,0.30063897,0.31235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.08589685,0.12103647,0.15617609,0.19131571,0.22645533,0.22645533,0.22645533,0.22645533,0.22645533,0.22645533,0.19912452,0.1756981,0.14836729,0.12494087,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.046852827,0.039044023,0.03513962,0.031235218,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.058566034,0.093705654,0.12884527,0.1639849,0.19912452,0.26549935,0.3318742,0.39434463,0.46071947,0.5231899,0.42167544,0.31625658,0.21083772,0.10541886,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.078088045,0.12884527,0.1835069,0.23426414,0.28892577,0.27330816,0.25769055,0.24207294,0.22645533,0.21083772,0.28892577,0.3631094,0.43729305,0.5114767,0.58566034,0.5231899,0.46071947,0.39824903,0.3357786,0.27330816,0.359205,0.44510186,0.5309987,0.61689556,0.698888,0.58175594,0.46462387,0.3474918,0.23035973,0.113227665,0.09761006,0.08199245,0.06637484,0.05075723,0.039044023,0.14836729,0.26159495,0.37482262,0.48805028,0.60127795,0.5114767,0.42167544,0.3318742,0.23816854,0.14836729,0.19912452,0.24988174,0.30063897,0.3513962,0.39824903,1.2298868,2.0615244,2.8892577,3.7208953,4.548629,4.5291066,4.5095844,4.4900627,4.4705405,4.4510183,3.978586,3.5100577,3.0415294,2.5690966,2.1005683,2.1981785,2.2996929,2.4012074,2.4988174,2.6003318,2.6432803,2.690133,2.7330816,2.7799344,2.8267872,2.3738766,1.9248703,1.475864,1.0268579,0.57394713,0.75354964,0.93315214,1.116659,1.2962615,1.475864,1.6437533,1.8116426,1.9756275,2.1435168,2.3114061,2.0654287,1.8194515,1.5695697,1.3235924,1.0737107,1.0893283,1.1010414,1.1127546,1.1244678,1.1361811,1.6515622,2.1630387,2.6745155,3.1859922,3.7013733,3.4007344,3.1000953,2.7994564,2.4988174,2.1981785,1.8897307,1.5812829,1.2689307,0.96048295,0.6481308,0.59346914,0.5388075,0.48414588,0.42948425,0.37482262,0.3240654,0.26940376,0.21864653,0.1639849,0.113227665,0.14055848,0.1678893,0.19522011,0.22255093,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.30844778,0.61689556,0.92143893,1.2298868,1.5383345,1.2455044,0.95267415,0.659844,0.3670138,0.07418364,0.23426414,0.39434463,0.5544251,0.7145056,0.8745861,0.698888,0.5231899,0.3513962,0.1756981,0.0,0.042948425,0.08589685,0.12884527,0.1717937,0.21083772,0.60127795,0.9917182,1.3821584,1.7725986,2.1630387,2.5808098,2.998581,3.416352,3.8341231,4.251894,4.1308575,4.0137253,3.8965936,3.7794614,3.6623292,4.591577,5.520825,6.453977,7.3832245,8.312472,8.94889,9.589212,10.22563,10.862047,11.498465,13.212498,14.92653,16.636658,18.35069,20.06082,21.509352,22.953981,24.39861,25.843239,27.287867,25.222439,23.15701,21.091581,19.026152,16.960724,15.363823,13.766922,12.170022,10.573121,8.976221,8.347612,7.719003,7.094299,6.46569,5.8370814,5.466163,5.099149,4.728231,4.357313,3.9863946,3.7560349,3.521771,3.2914112,3.057147,2.8267872,2.8306916,2.8345962,2.8385005,2.8463092,2.8502135,2.4988174,2.1513257,1.7999294,1.4485333,1.1010414,0.9058213,0.7106012,0.5153811,0.32016098,0.12494087,0.1796025,0.23426414,0.28892577,0.3435874,0.39824903,0.5505207,0.698888,0.8511597,0.999527,1.1517987,0.94486535,0.7418364,0.5349031,0.3318742,0.12494087,0.13665408,0.14446288,0.15617609,0.1639849,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19912452,0.39434463,0.59346914,0.78868926,0.9878138,0.78868926,0.59346914,0.39434463,0.19912452,0.0,0.046852827,0.08980125,0.13665408,0.1796025,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.078088045,0.15617609,0.23426414,0.30844778,0.38653582,0.359205,0.3318742,0.30454338,0.27721256,0.24988174,0.27330816,0.30063897,0.3240654,0.3513962,0.37482262,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.12884527,0.1796025,0.23426414,0.28502136,0.3357786,0.3357786,0.3357786,0.3357786,0.3357786,0.3357786,0.30063897,0.26159495,0.22645533,0.18741131,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.078088045,0.11713207,0.15617609,0.19912452,0.23816854,0.27330816,0.30844778,0.3435874,0.37872702,0.41386664,0.3318742,0.24597734,0.1639849,0.08199245,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.10932326,0.1835069,0.25378615,0.3279698,0.39824903,0.37872702,0.3553006,0.3318742,0.30844778,0.28892577,0.38653582,0.48805028,0.58566034,0.6871748,0.78868926,0.698888,0.61299115,0.5231899,0.43729305,0.3513962,0.47633708,0.60518235,0.7340276,0.8589685,0.9878138,0.80430686,0.62079996,0.44119745,0.25769055,0.07418364,0.06637484,0.05466163,0.046852827,0.03513962,0.023426414,0.10151446,0.1756981,0.24988174,0.3240654,0.39824903,0.3513962,0.30454338,0.25769055,0.21083772,0.1639849,0.24988174,0.3357786,0.42557985,0.5114767,0.60127795,1.8467822,3.0883822,4.3338866,5.579391,6.824895,6.79366,6.7663293,6.735094,6.703859,6.676528,5.969831,5.263134,4.560342,3.853645,3.1508527,3.2992198,3.4514916,3.5998588,3.7482262,3.900498,3.9668727,4.0332475,4.1035266,4.169902,4.2362766,3.5491016,2.8619268,2.174752,1.4875772,0.80040246,0.93315214,1.0659018,1.1986516,1.3314011,1.4641509,1.7686942,2.077142,2.3855898,2.6940374,2.998581,2.6237583,2.2450314,1.8663043,1.4914817,1.1127546,1.0893283,1.0619974,1.038571,1.0112402,0.9878138,1.6359446,2.2879796,2.9361105,3.5881457,4.2362766,3.873167,3.513962,3.1508527,2.787743,2.4246337,2.1239948,1.8194515,1.5188124,1.2142692,0.9136301,0.8433509,0.77307165,0.7027924,0.63251317,0.5622339,0.46462387,0.3670138,0.26940376,0.1717937,0.07418364,0.13665408,0.19522011,0.25378615,0.31625658,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.20693332,0.40996224,0.61689556,0.8199245,1.0268579,0.8316377,0.63641757,0.44119745,0.24597734,0.05075723,0.30063897,0.5544251,0.80821127,1.0580931,1.3118792,1.0502841,0.78868926,0.5231899,0.26159495,0.0,0.058566034,0.113227665,0.1717937,0.23035973,0.28892577,0.8355421,1.3821584,1.9287747,2.4792955,3.0259118,3.1586614,3.2914112,3.4241607,3.5569105,3.6857557,3.5686235,3.4475873,3.3265507,3.2094188,3.0883822,3.7716527,4.4510183,5.134289,5.8175592,6.5008297,7.125534,7.7502384,8.374943,8.999647,9.6243515,11.424281,13.224211,15.024139,16.82407,18.623999,20.580105,22.53621,24.48841,26.444517,28.400621,26.49137,24.578213,22.668959,20.759706,18.850454,17.085665,15.320874,13.556085,11.791295,10.0265045,9.452558,8.878611,8.308568,7.734621,7.1606736,6.6843367,6.2040954,5.7238536,5.2436123,4.7633705,4.369026,3.978586,3.5842414,3.193801,2.7994564,2.920493,3.0415294,3.1586614,3.279698,3.4007344,3.0376248,2.6745155,2.3114061,1.9482968,1.5890918,1.3079748,1.0268579,0.74574083,0.46852827,0.18741131,0.26940376,0.3513962,0.43338865,0.5192855,0.60127795,0.8238289,1.0502841,1.2767396,1.4992905,1.7257458,1.4172981,1.1088502,0.80430686,0.4958591,0.18741131,0.20302892,0.21864653,0.23426414,0.24597734,0.26159495,0.21083772,0.15617609,0.10541886,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26549935,0.5309987,0.79649806,1.0580931,1.3235924,1.0580931,0.79649806,0.5309987,0.26549935,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10932326,0.21864653,0.3318742,0.44119745,0.5505207,0.48805028,0.42948425,0.3709182,0.30844778,0.24988174,0.28892577,0.3240654,0.3631094,0.39824903,0.43729305,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.1717937,0.23816854,0.30844778,0.37872702,0.44900626,0.44900626,0.44900626,0.44900626,0.44900626,0.44900626,0.39824903,0.3513962,0.30063897,0.24988174,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.093705654,0.14055848,0.1835069,0.23035973,0.27330816,0.28111696,0.28502136,0.28892577,0.29673457,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.14055848,0.23426414,0.3279698,0.42167544,0.5114767,0.48414588,0.45291066,0.42167544,0.39434463,0.3631094,0.48805028,0.61299115,0.737932,0.8628729,0.9878138,0.8745861,0.76135844,0.6481308,0.5388075,0.42557985,0.59346914,0.76526284,0.93315214,1.1049459,1.2767396,1.0268579,0.78088045,0.5309987,0.28502136,0.039044023,0.031235218,0.027330816,0.023426414,0.015617609,0.011713207,0.05075723,0.08589685,0.12494087,0.1639849,0.19912452,0.19522011,0.19131571,0.1835069,0.1796025,0.1756981,0.30063897,0.42557985,0.5505207,0.6754616,0.80040246,2.4597735,4.1191444,5.7785153,7.4417906,9.101162,9.058213,9.019169,8.980125,8.941081,8.898132,7.9610763,7.0201154,6.0791545,5.138193,4.2011366,4.4002614,4.5993857,4.7985106,5.001539,5.2006636,5.290465,5.380266,5.4700675,5.559869,5.64967,4.7243266,3.7989833,2.87364,1.9482968,1.0268579,1.1088502,1.1947471,1.2806439,1.3665408,1.4485333,1.8975395,2.3465457,2.7916477,3.240654,3.6857557,3.1781836,2.6706111,2.1630387,1.6593709,1.1517987,1.0893283,1.0268579,0.96438736,0.9019169,0.8394465,1.6242313,2.4129205,3.2016098,3.9863946,4.775084,4.349504,3.9239242,3.4983444,3.076669,2.6510892,2.3543546,2.0615244,1.7647898,1.4680552,1.175225,1.0893283,1.0034313,0.92143893,0.8355421,0.74964523,0.60908675,0.46462387,0.3240654,0.1796025,0.039044023,0.12884527,0.22255093,0.31625658,0.40605783,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.20693332,0.30844778,0.40996224,0.5114767,0.41386664,0.31625658,0.21864653,0.12103647,0.023426414,0.3709182,0.7145056,1.0580931,1.4055848,1.7491722,1.4016805,1.0502841,0.698888,0.3513962,0.0,0.07418364,0.14446288,0.21864653,0.28892577,0.3631094,1.0659018,1.7725986,2.4792955,3.182088,3.8887846,3.736513,3.5842414,3.4280653,3.2757936,3.1235218,3.0024853,2.8814487,2.7565079,2.6354716,2.514435,2.9478238,3.3812122,3.8185053,4.251894,4.689187,5.298274,5.911265,6.524256,7.137247,7.7502384,9.636065,11.525795,13.411622,15.3013525,17.18718,19.650856,22.118439,24.582117,27.045794,29.513376,27.756395,26.003319,24.246338,22.493261,20.73628,18.8036,16.870922,14.938243,13.005564,11.076789,10.557504,10.0382185,9.522837,9.0035515,8.488171,7.898606,7.309041,6.715572,6.126007,5.5364423,4.985922,4.4314966,3.8809757,3.3265507,2.77603,3.0102942,3.2445583,3.4788225,3.7130866,3.951255,3.5764325,3.2016098,2.8267872,2.4480603,2.0732377,1.7101282,1.3431144,0.98000497,0.61689556,0.24988174,0.359205,0.46852827,0.58175594,0.6910792,0.80040246,1.1010414,1.4016805,1.698415,1.999054,2.2996929,1.8897307,1.4797685,1.0698062,0.659844,0.24988174,0.26940376,0.28892577,0.30844778,0.3318742,0.3513962,0.28111696,0.21083772,0.14055848,0.07027924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3318742,0.6637484,0.9956226,1.3314011,1.6632754,1.3314011,0.9956226,0.6637484,0.3318742,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14055848,0.28502136,0.42557985,0.5700427,0.7106012,0.62079996,0.5270943,0.43338865,0.3435874,0.24988174,0.30063897,0.3513962,0.39824903,0.44900626,0.4997635,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.21083772,0.30063897,0.38653582,0.47633708,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.4997635,0.43729305,0.37482262,0.31235218,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.113227665,0.1639849,0.21083772,0.26159495,0.31235218,0.28892577,0.26159495,0.23816854,0.21083772,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.1756981,0.28892577,0.39824903,0.5114767,0.62470436,0.58566034,0.5505207,0.5114767,0.47633708,0.43729305,0.58566034,0.737932,0.8862993,1.038571,1.1869383,1.0502841,0.9136301,0.77307165,0.63641757,0.4997635,0.7106012,0.92534333,1.1361811,1.3509232,1.5617609,1.2494087,0.93705654,0.62470436,0.31235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.3513962,0.5114767,0.6754616,0.8394465,0.999527,3.076669,5.1499066,7.223144,9.300286,11.373524,11.326671,11.275913,11.225157,11.174399,11.123642,9.948417,8.773191,7.601871,6.426646,5.251421,5.5013027,5.7511845,6.001066,6.250948,6.5008297,6.6140575,6.7233806,6.8366084,6.949836,7.0630636,5.899552,4.73604,3.5764325,2.4129205,1.2494087,1.2884527,1.3235924,1.3626363,1.4016805,1.43682,2.0263848,2.612045,3.2016098,3.78727,4.376835,3.736513,3.1000953,2.463678,1.8233559,1.1869383,1.0893283,0.9878138,0.8862993,0.78868926,0.6871748,1.6125181,2.5378613,3.4632049,4.388548,5.3138914,4.825841,4.337791,3.8497405,3.3616903,2.87364,2.5886188,2.2996929,2.0107672,1.7257458,1.43682,1.33921,1.2376955,1.1361811,1.038571,0.93705654,0.74964523,0.5622339,0.37482262,0.18741131,0.0,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.43729305,0.8745861,1.3118792,1.7491722,2.1864653,1.7491722,1.3118792,0.8745861,0.43729305,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,1.3001659,2.1630387,3.0259118,3.8887846,4.7516575,4.3143644,3.873167,3.435874,2.998581,2.5612879,2.436347,2.3114061,2.1864653,2.0615244,1.9365835,2.1239948,2.3114061,2.4988174,2.6862288,2.87364,3.474918,4.0761957,4.6735697,5.2748475,5.8761253,7.8517528,9.823476,11.799104,13.774731,15.750359,18.725513,21.700668,24.675823,27.650976,30.626131,29.025326,27.424522,25.823717,24.226816,22.62601,20.525442,18.424873,16.324306,14.223738,12.123169,11.66245,11.20173,10.737106,10.276386,9.811763,9.112875,8.413987,7.7111945,7.012306,6.3134184,5.5989127,4.8883114,4.173806,3.4632049,2.7486992,3.1000953,3.4514916,3.7989833,4.1503797,4.5017757,4.1113358,3.7247996,3.338264,2.951728,2.5612879,2.1122816,1.6632754,1.2142692,0.76135844,0.31235218,0.44900626,0.58566034,0.7262188,0.8628729,0.999527,1.3743496,1.7491722,2.1239948,2.4988174,2.87364,2.3621633,1.8506867,1.33921,0.8238289,0.31235218,0.3357786,0.3631094,0.38653582,0.41386664,0.43729305,0.3513962,0.26159495,0.1756981,0.08589685,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.39824903,0.80040246,1.1986516,1.6008049,1.999054,1.6008049,1.1986516,0.80040246,0.39824903,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1756981,0.3513962,0.5231899,0.698888,0.8745861,0.74964523,0.62470436,0.4997635,0.37482262,0.24988174,0.31235218,0.37482262,0.43729305,0.4997635,0.5622339,0.23816854,0.21083772,0.1835069,0.15617609,0.12884527,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.046852827,0.046852827,0.042948425,0.039044023,0.039044023,0.046852827,0.05075723,0.058566034,0.06637484,0.07418364,0.06637484,0.05466163,0.046852827,0.03513962,0.023426414,0.058566034,0.093705654,0.12884527,0.1639849,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.15617609,0.19912452,0.23816854,0.28111696,0.3240654,0.37482262,0.42557985,0.47633708,0.5231899,0.57394713,0.6442264,0.7145056,0.78478485,0.8550641,0.92534333,0.8511597,0.77307165,0.698888,0.62470436,0.5505207,0.48024148,0.40996224,0.339683,0.26940376,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.058566034,0.06637484,0.07418364,0.078088045,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.14836729,0.19912452,0.24988174,0.30063897,0.3513962,0.31625658,0.28111696,0.24597734,0.21083772,0.1756981,0.30844778,0.44510186,0.58175594,0.7145056,0.8511597,0.71841,0.58956474,0.46071947,0.3318742,0.19912452,0.30454338,0.40996224,0.5153811,0.62079996,0.7262188,0.7106012,0.698888,0.6871748,0.6754616,0.6637484,0.75354964,0.8472553,0.94096094,1.0307622,1.1244678,1.0815194,1.038571,0.9956226,0.95657855,0.9136301,1.0698062,1.2259823,1.3860629,1.542239,1.698415,1.4836729,1.2650263,1.0463798,0.8316377,0.61299115,0.64032197,0.6676528,0.6949836,0.7223144,0.74964523,0.94876975,1.1517987,1.3509232,1.5500476,1.7491722,1.5617609,1.3704453,1.1791295,0.9917182,0.80040246,1.1674163,1.53443,1.901444,2.2684577,2.639376,4.0137253,5.3919797,6.7702336,8.148487,9.526741,9.425227,9.323712,9.226103,9.124588,9.023073,8.093826,7.1606736,6.2275214,5.2943697,4.3612175,4.564246,4.7672753,4.970304,5.173333,5.376362,5.4583545,5.5403466,5.6223392,5.704332,5.786324,4.841459,3.892689,2.9439192,1.999054,1.0502841,1.077615,1.1049459,1.1322767,1.1596074,1.1869383,1.8389735,2.4871042,3.1391394,3.78727,4.4393053,4.1503797,3.8614538,3.5764325,3.2875066,2.998581,2.9322062,2.8658314,2.7994564,2.7291772,2.6628022,3.2172275,3.7716527,4.3260775,4.884407,5.4388323,4.903929,4.3729305,3.8419318,3.3070288,2.77603,2.4831998,2.1903696,1.8975395,1.6047094,1.3118792,1.2415999,1.1713207,1.1010414,1.0307622,0.96438736,0.77307165,0.58566034,0.39824903,0.21083772,0.023426414,0.14446288,0.26549935,0.38653582,0.5036679,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10932326,0.093705654,0.078088045,0.06637484,0.05075723,0.058566034,0.06637484,0.07418364,0.078088045,0.08589685,0.30454338,0.5231899,0.7418364,0.95657855,1.175225,1.0424755,0.9097257,0.77697605,0.6442264,0.5114767,1.0268579,1.542239,2.05762,2.5730011,3.0883822,2.9361105,2.7838387,2.631567,2.4792955,2.3231194,2.241127,2.15523,2.069333,1.9834363,1.901444,2.522244,3.1469483,3.767748,4.388548,5.0132523,4.7087092,4.4041657,4.095718,3.7911747,3.4866312,3.2211318,2.9556324,2.6940374,2.4285383,2.1630387,2.2489357,2.330928,2.416825,2.5027218,2.5886188,3.018103,3.4514916,3.8848803,4.318269,4.7516575,6.4110284,8.074304,9.737579,11.400854,13.06413,15.9104395,18.756748,21.606962,24.453272,27.29958,26.549934,25.80029,25.050644,24.300999,23.551353,21.923218,20.295082,18.666946,17.03881,15.410676,14.641508,13.872341,13.103174,12.334006,11.560935,10.764437,9.967939,9.171441,8.371038,7.57454,6.824895,6.0752497,5.3256044,4.575959,3.8263142,3.9434462,4.0605783,4.1777105,4.2948427,4.4119744,4.068387,3.7287042,3.3851168,3.0415294,2.7018464,2.3231194,1.9443923,1.5656652,1.1908426,0.81211567,0.8160201,0.8160201,0.8199245,0.8238289,0.8238289,1.1361811,1.4485333,1.7608855,2.0732377,2.3855898,1.9834363,1.5773785,1.1713207,0.76916724,0.3631094,0.359205,0.359205,0.3553006,0.3513962,0.3513962,0.42167544,0.49195468,0.5583295,0.62860876,0.698888,0.8667773,1.0307622,1.1947471,1.358732,1.5266213,1.4680552,1.4094892,1.3509232,1.2962615,1.2376955,1.0151446,0.79259366,0.5700427,0.3474918,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.32016098,0.64032197,0.96048295,1.2806439,1.6008049,1.2806439,0.96048295,0.64032197,0.32016098,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.15617609,0.30844778,0.46462387,0.62079996,0.77307165,0.6715572,0.5661383,0.46071947,0.3553006,0.24988174,0.30063897,0.3553006,0.40605783,0.46071947,0.5114767,0.47633708,0.42167544,0.3631094,0.30844778,0.25378615,0.19912452,0.1796025,0.16008049,0.14055848,0.12103647,0.10151446,0.093705654,0.08980125,0.08589685,0.078088045,0.07418364,0.08980125,0.10541886,0.12103647,0.13665408,0.14836729,0.12884527,0.10932326,0.08980125,0.07027924,0.05075723,0.07027924,0.08980125,0.10932326,0.12884527,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.08980125,0.13665408,0.1796025,0.22645533,0.30844778,0.39434463,0.48024148,0.5661383,0.6481308,0.7262188,0.80040246,0.8745861,0.94876975,1.0268579,1.077615,1.1283722,1.183034,1.2337911,1.2884527,1.1361811,0.9878138,0.8394465,0.6871748,0.5388075,0.46071947,0.38263142,0.30454338,0.22645533,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.13665408,0.12884527,0.12103647,0.113227665,0.10932326,0.10151446,0.113227665,0.12884527,0.14446288,0.16008049,0.1756981,0.14836729,0.12494087,0.10151446,0.07418364,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.18741131,0.23816854,0.28892577,0.3357786,0.38653582,0.3435874,0.29673457,0.25378615,0.20693332,0.1639849,0.46852827,0.77697605,1.0854238,1.3938715,1.698415,1.4290112,1.1557031,0.8823949,0.60908675,0.3357786,0.43338865,0.5309987,0.62860876,0.7262188,0.8238289,0.8394465,0.8511597,0.8628729,0.8745861,0.8862993,0.92143893,0.95657855,0.9917182,1.0268579,1.0619974,1.116659,1.1674163,1.2181735,1.2728351,1.3235924,1.4290112,1.5305257,1.6320401,1.7335546,1.8389735,1.7140326,1.5929961,1.4680552,1.3470187,1.2259823,1.2806439,1.3353056,1.3899672,1.4446288,1.4992905,1.901444,2.2996929,2.7018464,3.1000953,3.4983444,3.0805733,2.6667068,2.2489357,1.8311646,1.4133936,1.9834363,2.5573835,3.1313305,3.7013733,4.2753205,4.9546866,5.6340523,6.3134184,6.996689,7.676055,7.523783,7.375416,7.223144,7.0747766,6.9264097,6.2353306,5.5442514,4.853172,4.165997,3.474918,3.631094,3.7833657,3.9395418,4.095718,4.251894,4.3026514,4.3534083,4.40807,4.4588275,4.513489,3.7794614,3.049338,2.3153105,1.5812829,0.8511597,0.8667773,0.8862993,0.9019169,0.92143893,0.93705654,1.6515622,2.3621633,3.076669,3.78727,4.5017757,4.564246,4.6267166,4.689187,4.7516575,4.814128,4.7789884,4.743849,4.7087092,4.6735697,4.6384296,4.8219366,5.009348,5.192855,5.376362,5.563773,4.985922,4.40807,3.8302186,3.252367,2.6745155,2.377781,2.0810463,1.7843118,1.4836729,1.1869383,1.1478943,1.1088502,1.0659018,1.0268579,0.9878138,0.80040246,0.61299115,0.42557985,0.23816854,0.05075723,0.1639849,0.28111696,0.39434463,0.5114767,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.21864653,0.19131571,0.16008049,0.12884527,0.10151446,0.113227665,0.12884527,0.14446288,0.16008049,0.1756981,0.60908675,1.0463798,1.4797685,1.9131571,2.35045,2.084951,1.8194515,1.5539521,1.2884527,1.0268579,1.6164225,2.2098918,2.803361,3.39683,3.9863946,4.1191444,4.251894,4.3846436,4.5173936,4.650143,4.3924527,4.134762,3.8770714,3.619381,3.3616903,3.7443218,4.126953,4.5095844,4.892216,5.2748475,5.1030536,4.93126,4.755562,4.5837684,4.4119744,4.0059166,3.6037633,3.1977055,2.7916477,2.3855898,2.3699722,2.3543546,2.3348327,2.3192148,2.2996929,2.5651922,2.8306916,3.096191,3.3616903,3.6232853,4.9742084,6.3251314,7.676055,9.023073,10.373997,13.095366,15.816733,18.534197,21.255566,23.97303,24.074545,24.17606,24.273668,24.375183,24.476698,23.320995,22.16529,21.009588,19.853886,18.698183,17.620567,16.546856,15.469242,14.391626,13.314012,12.415999,11.521891,10.627783,9.733675,8.835662,8.050878,7.262188,6.473499,5.688714,4.900025,4.786797,4.6696653,4.5564375,4.4393053,4.3260775,4.029343,3.7287042,3.4319696,3.135235,2.8385005,2.533957,2.2294137,1.9209659,1.6164225,1.3118792,1.1791295,1.0463798,0.9136301,0.78088045,0.6481308,0.9019169,1.1517987,1.4016805,1.6515622,1.901444,1.6008049,1.3040704,1.0073358,0.7106012,0.41386664,0.38263142,0.3513962,0.3240654,0.29283017,0.26159495,0.49195468,0.71841,0.94486535,1.1713207,1.4016805,1.7296503,2.0615244,2.3894942,2.7213683,3.049338,2.9361105,2.8189783,2.7057507,2.5886188,2.475391,2.018576,1.5617609,1.1010414,0.6442264,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23816854,0.48024148,0.71841,0.96048295,1.1986516,0.96048295,0.71841,0.48024148,0.23816854,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.13665408,0.26940376,0.40605783,0.5388075,0.6754616,0.58956474,0.5036679,0.42167544,0.3357786,0.24988174,0.29283017,0.3357786,0.37872702,0.42167544,0.46071947,0.7106012,0.62860876,0.5466163,0.46462387,0.38263142,0.30063897,0.26940376,0.23816854,0.21083772,0.1796025,0.14836729,0.14055848,0.13665408,0.12884527,0.12103647,0.113227665,0.13665408,0.15617609,0.1796025,0.20302892,0.22645533,0.19522011,0.1639849,0.13665408,0.10541886,0.07418364,0.078088045,0.08589685,0.08980125,0.093705654,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06637484,0.13665408,0.20302892,0.26940376,0.3357786,0.46462387,0.59346914,0.71841,0.8472553,0.97610056,1.0737107,1.175225,1.2767396,1.3743496,1.475864,1.5110037,1.5461433,1.5812829,1.6164225,1.6515622,1.4251068,1.1986516,0.97610056,0.74964523,0.5231899,0.44119745,0.3553006,0.26940376,0.1835069,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.1756981,0.1717937,0.1639849,0.16008049,0.15617609,0.14836729,0.1717937,0.19522011,0.21864653,0.23816854,0.26159495,0.22645533,0.18741131,0.14836729,0.113227665,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.22645533,0.27330816,0.3240654,0.37482262,0.42557985,0.3709182,0.31625658,0.26159495,0.20693332,0.14836729,0.62860876,1.1088502,1.5890918,2.069333,2.5495746,2.135708,1.7218413,1.3040704,0.8902037,0.47633708,0.5661383,0.6559396,0.74574083,0.8355421,0.92534333,0.96438736,0.999527,1.038571,1.0737107,1.1127546,1.0893283,1.0659018,1.0463798,1.0229534,0.999527,1.1478943,1.2962615,1.4407244,1.5890918,1.737459,1.7843118,1.8311646,1.8819219,1.9287747,1.9756275,1.9482968,1.9209659,1.893635,1.8663043,1.8389735,1.9209659,2.0029583,2.084951,2.1669433,2.2489357,2.8502135,3.4514916,4.0488653,4.650143,5.251421,4.60329,3.959064,3.3148375,2.6706111,2.0263848,2.803361,3.5803368,4.357313,5.134289,5.911265,5.8956475,5.8761253,5.860508,5.840986,5.825368,5.6262436,5.423215,5.22409,5.024966,4.825841,4.376835,3.9317331,3.4827268,3.0337205,2.5886188,2.6940374,2.803361,2.9087796,3.018103,3.1235218,3.1469483,3.1703746,3.193801,3.213323,3.2367494,2.7213683,2.2020829,1.6867018,1.1674163,0.6481308,0.6559396,0.6637484,0.6715572,0.679366,0.6871748,1.4641509,2.2372224,3.0141985,3.78727,4.564246,4.9742084,5.388075,5.801942,6.211904,6.6257706,6.621866,6.621866,6.617962,6.6140575,6.6140575,6.426646,6.2431393,6.055728,5.872221,5.688714,5.0640097,4.4432096,3.8185053,3.1977055,2.5769055,2.2723622,1.9717231,1.6671798,1.3665408,1.0619974,1.0541886,1.0424755,1.0307622,1.0229534,1.0112402,0.8238289,0.63641757,0.44900626,0.26159495,0.07418364,0.1835069,0.29673457,0.40605783,0.5153811,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.3318742,0.28502136,0.23816854,0.19522011,0.14836729,0.1717937,0.19522011,0.21864653,0.23816854,0.26159495,0.9136301,1.5656652,2.2216048,2.87364,3.5256753,3.1274261,2.7291772,2.330928,1.9365835,1.5383345,2.2059872,2.8775444,3.5491016,4.2167544,4.8883114,5.3060827,5.7238536,6.141625,6.559396,6.9732623,6.5437784,6.114294,5.6848097,5.2553253,4.825841,4.9663997,5.1108627,5.251421,5.395884,5.5364423,5.4973984,5.4583545,5.4193106,5.376362,5.337318,4.7907014,4.2479897,3.7013733,3.1586614,2.612045,2.4910088,2.3738766,2.25284,2.1318035,2.0107672,2.1083772,2.2059872,2.3035975,2.4012074,2.4988174,3.5373883,4.575959,5.610626,6.649197,7.687768,10.280292,12.872814,15.465338,18.057861,20.650383,21.599154,22.551826,23.500597,24.449368,25.398136,24.718771,24.0355,23.35223,22.668959,21.98569,20.60353,19.217468,17.831406,16.449247,15.063184,14.0714655,13.075843,12.084125,11.092407,10.100689,9.276859,8.449126,7.6252975,6.801469,5.9737353,5.6262436,5.278752,4.93126,4.5837684,4.2362766,3.9863946,3.7326086,3.4788225,3.2289407,2.9751544,2.7408905,2.5105307,2.2762666,2.0459068,1.8116426,1.5461433,1.2767396,1.0112402,0.7418364,0.47633708,0.6637484,0.8511597,1.038571,1.2259823,1.4133936,1.2220778,1.0307622,0.8433509,0.6520352,0.46071947,0.40605783,0.3474918,0.28892577,0.23426414,0.1756981,0.5583295,0.94486535,1.3314011,1.7140326,2.1005683,2.5964274,3.0883822,3.5842414,4.0801005,4.575959,4.4041657,4.2284675,4.056674,3.8848803,3.7130866,3.018103,2.3270237,1.6359446,0.94096094,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16008049,0.32016098,0.48024148,0.64032197,0.80040246,0.64032197,0.48024148,0.32016098,0.16008049,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.113227665,0.23035973,0.3435874,0.46071947,0.57394713,0.5114767,0.44510186,0.37872702,0.31625658,0.24988174,0.28111696,0.31625658,0.3474918,0.37872702,0.41386664,0.94876975,0.8394465,0.7301232,0.62079996,0.5114767,0.39824903,0.359205,0.32016098,0.28111696,0.23816854,0.19912452,0.19131571,0.1796025,0.1717937,0.16008049,0.14836729,0.1796025,0.21083772,0.23816854,0.26940376,0.30063897,0.26159495,0.21864653,0.1796025,0.14055848,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08980125,0.1796025,0.26940376,0.359205,0.44900626,0.62079996,0.78868926,0.96048295,1.1283722,1.3001659,1.4251068,1.5500476,1.6749885,1.7999294,1.9248703,1.9443923,1.9600099,1.9756275,1.9951496,2.0107672,1.7140326,1.4133936,1.1127546,0.81211567,0.5114767,0.42167544,0.3279698,0.23426414,0.14055848,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.062470436,0.10151446,0.13665408,0.1756981,0.21083772,0.21083772,0.20693332,0.20693332,0.20302892,0.19912452,0.23035973,0.26159495,0.28892577,0.32016098,0.3513962,0.30063897,0.24988174,0.19912452,0.14836729,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.042948425,0.08589685,0.12884527,0.1717937,0.21083772,0.26159495,0.31235218,0.3631094,0.41386664,0.46071947,0.39824903,0.3318742,0.26940376,0.20302892,0.13665408,0.78868926,1.4407244,2.096664,2.7486992,3.4007344,2.8424048,2.2840753,1.7257458,1.1713207,0.61299115,0.6949836,0.77697605,0.8589685,0.94096094,1.0268579,1.0893283,1.1517987,1.2142692,1.2767396,1.33921,1.2572175,1.1791295,1.097137,1.0190489,0.93705654,1.1791295,1.4212024,1.6632754,1.9092526,2.1513257,2.1435168,2.135708,2.1278992,2.1200905,2.1122816,2.1786566,2.2489357,2.3153105,2.3816853,2.4480603,2.5612879,2.6706111,2.7799344,2.8892577,2.998581,3.7989833,4.5993857,5.3997884,6.2001905,7.000593,6.126007,5.2553253,4.380739,3.5100577,2.639376,3.619381,4.60329,5.5832953,6.5672045,7.551114,6.8366084,6.1181984,5.4036927,4.689187,3.9746814,3.7247996,3.474918,3.2250361,2.9751544,2.7252727,2.5183394,2.3153105,2.1083772,1.9053483,1.698415,1.7608855,1.8194515,1.8819219,1.9404879,1.999054,1.9912452,1.9834363,1.9756275,1.9717231,1.9639144,1.6593709,1.358732,1.0541886,0.75354964,0.44900626,0.44900626,0.44510186,0.44119745,0.44119745,0.43729305,1.2767396,2.1122816,2.951728,3.78727,4.6267166,5.388075,6.1494336,6.910792,7.676055,8.437413,8.468649,8.495979,8.527214,8.55845,8.58578,8.031356,7.47693,6.9225054,6.36808,5.813655,5.1460023,4.478349,3.8106966,3.1430438,2.475391,2.1669433,1.8584955,1.5539521,1.2455044,0.93705654,0.95657855,0.97610056,0.9956226,1.0190489,1.038571,0.8511597,0.6637484,0.47633708,0.28892577,0.10151446,0.20693332,0.30844778,0.41386664,0.5192855,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.44119745,0.37872702,0.32016098,0.26159495,0.19912452,0.23035973,0.26159495,0.28892577,0.32016098,0.3513962,1.2181735,2.0888553,2.959537,3.8302186,4.7009,4.169902,3.638903,3.1118085,2.5808098,2.0498111,2.7994564,3.5451972,4.290938,5.040583,5.786324,6.4891167,7.191909,7.8947015,8.597494,9.300286,8.699008,8.093826,7.492548,6.89127,6.2860875,6.1884775,6.0908675,5.9932575,5.8956475,5.801942,5.891743,5.985449,6.0791545,6.168956,6.262661,5.579391,4.892216,4.2089458,3.521771,2.8385005,2.6159496,2.3933985,2.1708477,1.9482968,1.7257458,1.6554666,1.5851873,1.5149081,1.4446288,1.3743496,2.1005683,2.8267872,3.5491016,4.2753205,5.001539,7.465217,9.928895,12.396477,14.860155,17.323833,19.123762,20.92369,22.723621,24.52355,26.32348,26.116547,25.905708,25.694872,25.484034,25.273195,23.58259,21.891983,20.197474,18.506866,16.812357,15.723028,14.633699,13.544372,12.4511385,11.361811,10.498938,9.636065,8.773191,7.914223,7.0513506,6.4695945,5.891743,5.309987,4.728231,4.1503797,3.9434462,3.736513,3.5256753,3.3187418,3.1118085,2.951728,2.7916477,2.631567,2.4714866,2.3114061,1.9092526,1.5070993,1.1049459,0.7027924,0.30063897,0.42557985,0.5505207,0.6754616,0.80040246,0.92534333,0.8433509,0.76135844,0.679366,0.59346914,0.5114767,0.42557985,0.3435874,0.25769055,0.1717937,0.08589685,0.62860876,1.1713207,1.7140326,2.2567444,2.7994564,3.4593005,4.1191444,4.7789884,5.4388323,6.098676,5.8683167,5.6418614,5.4115014,5.181142,4.950782,4.0215344,3.096191,2.1669433,1.2415999,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,0.32016098,0.23816854,0.16008049,0.078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.093705654,0.19131571,0.28502136,0.37872702,0.47633708,0.42948425,0.38653582,0.339683,0.29673457,0.24988174,0.27330816,0.29673457,0.31625658,0.339683,0.3631094,1.1869383,1.0502841,0.9136301,0.77307165,0.63641757,0.4997635,0.44900626,0.39824903,0.3513962,0.30063897,0.24988174,0.23816854,0.22645533,0.21083772,0.19912452,0.18741131,0.22645533,0.26159495,0.30063897,0.3357786,0.37482262,0.3240654,0.27330816,0.22645533,0.1756981,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.113227665,0.22645533,0.3357786,0.44900626,0.5622339,0.77307165,0.9878138,1.1986516,1.4133936,1.6242313,1.7765031,1.9248703,2.0732377,2.2255092,2.3738766,2.3738766,2.3738766,2.3738766,2.3738766,2.3738766,1.999054,1.6242313,1.2494087,0.8745861,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.28892577,0.3240654,0.3631094,0.39824903,0.43729305,0.37482262,0.31235218,0.24988174,0.18741131,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.30063897,0.3513962,0.39824903,0.44900626,0.4997635,0.42557985,0.3513962,0.27330816,0.19912452,0.12494087,0.94876975,1.7765031,2.6003318,3.4241607,4.251894,3.5491016,2.8502135,2.1513257,1.4485333,0.74964523,0.8238289,0.9019169,0.97610056,1.0502841,1.1244678,1.2142692,1.3001659,1.3860629,1.475864,1.5617609,1.4251068,1.2884527,1.1517987,1.0112402,0.8745861,1.2142692,1.5500476,1.8858263,2.2255092,2.5612879,2.4988174,2.436347,2.3738766,2.3114061,2.2489357,2.4129205,2.5769055,2.736986,2.900971,3.0610514,3.2016098,3.338264,3.474918,3.611572,3.7482262,4.7516575,5.7511845,6.7507114,7.7502384,8.749765,7.648724,6.551587,5.4505453,4.349504,3.2484627,4.4393053,5.6262436,6.813182,8.00012,9.187058,7.773665,6.364176,4.950782,3.5373883,2.1239948,1.8233559,1.5266213,1.2259823,0.92534333,0.62470436,0.6637484,0.698888,0.737932,0.77307165,0.81211567,0.8238289,0.8394465,0.8511597,0.8628729,0.8745861,0.8394465,0.80040246,0.76135844,0.7262188,0.6871748,0.60127795,0.5114767,0.42557985,0.3357786,0.24988174,0.23816854,0.22645533,0.21083772,0.19912452,0.18741131,1.0893283,1.9873407,2.8892577,3.78727,4.689187,5.7980375,6.910792,8.023546,9.136301,10.249056,10.311526,10.373997,10.436467,10.498938,10.561408,9.636065,8.710721,7.7892823,6.8639393,5.938596,5.22409,4.513489,3.7989833,3.0883822,2.3738766,2.0615244,1.7491722,1.43682,1.1244678,0.81211567,0.8628729,0.9136301,0.96438736,1.0112402,1.0619974,0.8745861,0.6871748,0.4997635,0.31235218,0.12494087,0.22645533,0.3240654,0.42557985,0.5231899,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.0,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,0.5505207,0.47633708,0.39824903,0.3240654,0.24988174,0.28892577,0.3240654,0.3631094,0.39824903,0.43729305,1.5266213,2.612045,3.7013733,4.786797,5.8761253,5.212377,4.548629,3.8887846,3.2250361,2.5612879,3.3890212,4.21285,5.036679,5.8644123,6.688241,7.676055,8.663869,9.651682,10.6355915,11.623405,10.850334,10.073358,9.300286,8.52331,7.7502384,7.4105554,7.0747766,6.7389984,6.3993154,6.0635366,6.2860875,6.5125427,6.7389984,6.9615493,7.1880045,6.364176,5.5364423,4.7126136,3.8887846,3.0610514,2.736986,2.4129205,2.0888553,1.7608855,1.43682,1.1986516,0.96438736,0.7262188,0.48805028,0.24988174,0.6637484,1.0737107,1.4875772,1.901444,2.3114061,4.650143,6.98888,9.323712,11.66245,14.001186,16.64837,19.29946,21.95055,24.601639,27.248823,27.514322,27.775917,28.037512,28.299107,28.560703,26.56165,24.562595,22.563541,20.560583,18.56153,17.37459,16.187653,15.000713,13.813775,12.626837,11.72492,10.826907,9.924991,9.023073,8.125061,7.3129454,6.5008297,5.688714,4.8765984,4.0605783,3.900498,3.736513,3.5764325,3.4124475,3.2484627,3.1625657,3.076669,2.9868677,2.900971,2.8111696,2.2762666,1.737459,1.1986516,0.6637484,0.12494087,0.18741131,0.24988174,0.31235218,0.37482262,0.43729305,0.46071947,0.48805028,0.5114767,0.5388075,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.698888,1.4016805,2.1005683,2.7994564,3.4983444,4.3260775,5.1499066,5.9737353,6.801469,7.6252975,7.336372,7.0513506,6.7624245,6.473499,6.1884775,5.024966,3.8614538,2.7018464,1.5383345,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.3513962,0.3240654,0.30063897,0.27330816,0.24988174,0.26159495,0.27330816,0.28892577,0.30063897,0.31235218,0.94876975,0.8394465,0.7301232,0.62079996,0.5114767,0.39824903,0.359205,0.32016098,0.28111696,0.23816854,0.19912452,0.19131571,0.1796025,0.1717937,0.16008049,0.14836729,0.19912452,0.24597734,0.29283017,0.339683,0.38653582,0.359205,0.3318742,0.30454338,0.27721256,0.24988174,0.23816854,0.22645533,0.21083772,0.19912452,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.07418364,0.13274968,0.19131571,0.25378615,0.31235218,0.3318742,0.3513962,0.3709182,0.39434463,0.41386664,0.359205,0.30844778,0.25378615,0.20302892,0.14836729,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.13665408,0.24988174,0.3631094,0.47633708,0.58566034,0.80430686,1.0229534,1.2415999,1.456342,1.6749885,1.7413634,1.8116426,1.8780174,1.9443923,2.0107672,1.9912452,1.9678187,1.9443923,1.9209659,1.901444,1.6008049,1.3001659,0.999527,0.698888,0.39824903,0.32016098,0.23816854,0.16008049,0.078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.046852827,0.039044023,0.03513962,0.031235218,0.023426414,0.093705654,0.16008049,0.22645533,0.29673457,0.3631094,0.30063897,0.23816854,0.1756981,0.113227665,0.05075723,0.078088045,0.10932326,0.14055848,0.1717937,0.19912452,0.23816854,0.28111696,0.32016098,0.359205,0.39824903,0.4958591,0.59346914,0.6910792,0.78868926,0.8862993,0.8862993,0.8862993,0.8862993,0.8862993,0.8862993,0.8394465,0.79259366,0.74574083,0.698888,0.6481308,0.61689556,0.58175594,0.5466163,0.5114767,0.47633708,0.4958591,0.5153811,0.5349031,0.5544251,0.57394713,0.5075723,0.44119745,0.3709182,0.30454338,0.23816854,0.9136301,1.5890918,2.260649,2.9361105,3.611572,3.1469483,2.67842,2.2098918,1.7413634,1.2767396,1.4290112,1.5812829,1.7335546,1.8858263,2.0380979,2.1981785,2.3621633,2.5261483,2.6862288,2.8502135,2.893162,2.9400148,2.9868677,3.0298162,3.076669,3.1235218,3.174279,3.2250361,3.2757936,3.3265507,3.2640803,3.2055142,3.1469483,3.084478,3.0259118,3.0649557,3.1039999,3.1469483,3.1859922,3.2250361,3.3187418,3.416352,3.5100577,3.6037633,3.7013733,4.548629,5.3997884,6.250948,7.098203,7.9493628,6.9537406,5.958118,4.9663997,3.970777,2.9751544,3.9629683,4.950782,5.938596,6.9264097,7.914223,6.9225054,5.930787,4.942973,3.951255,2.9634414,2.6862288,2.4090161,2.1318035,1.8506867,1.5734742,1.5305257,1.4836729,1.4407244,1.3938715,1.3509232,1.3314011,1.3157835,1.2962615,1.2806439,1.261122,1.1596074,1.0580931,0.95657855,0.8511597,0.74964523,0.7066968,0.6637484,0.62079996,0.58175594,0.5388075,0.698888,0.8589685,1.0190489,1.1791295,1.33921,2.2216048,3.1079042,3.9942036,4.8765984,5.7628975,6.575013,7.387129,8.1992445,9.01136,9.823476,9.8195715,9.815667,9.811763,9.803954,9.80005,9.0035515,8.203149,7.406651,6.610153,5.813655,5.22409,4.630621,4.041056,3.4514916,2.8619268,2.5066261,2.1474214,1.7882162,1.4329157,1.0737107,1.0893283,1.1049459,1.1205635,1.1361811,1.1517987,0.96829176,0.78478485,0.60127795,0.42167544,0.23816854,0.29283017,0.3474918,0.40215343,0.45681506,0.5114767,0.45681506,0.40215343,0.3474918,0.29283017,0.23816854,0.39434463,0.5466163,0.7027924,0.8589685,1.0112402,0.94096094,0.8667773,0.79649806,0.7223144,0.6481308,0.98390937,1.319688,1.6554666,1.9912452,2.3231194,3.1391394,3.951255,4.7633705,5.575486,6.387602,5.688714,4.985922,4.2870336,3.5881457,2.8892577,3.6349986,4.380739,5.1303844,5.8761253,6.6257706,7.480835,8.335898,9.190963,10.046027,10.901091,10.09288,9.284669,8.476458,7.6682463,6.8639393,6.6687193,6.473499,6.278279,6.083059,5.8878384,6.0713453,6.2587566,6.4422636,6.6257706,6.813182,6.1572423,5.5013027,4.8492675,4.193328,3.5373883,3.213323,2.8892577,2.5612879,2.2372224,1.9131571,1.6437533,1.3782539,1.1088502,0.8433509,0.57394713,0.8394465,1.1049459,1.3704453,1.6359446,1.901444,3.7833657,5.6652875,7.5472097,9.4291315,11.311053,13.509232,15.7035055,17.89778,20.092054,22.286327,22.840754,23.391273,23.9457,24.49622,25.050644,23.926178,22.801708,21.673336,20.548868,19.4244,18.35069,17.27698,16.199366,15.125654,14.051944,13.134409,12.220779,11.303245,10.389614,9.475985,8.574067,7.6682463,6.7663293,5.8644123,4.9624953,4.829746,4.6969957,4.564246,4.4314966,4.298747,4.041056,3.7794614,3.521771,3.260176,2.998581,2.463678,1.9287747,1.3938715,0.8589685,0.3240654,0.3474918,0.3709182,0.39434463,0.41386664,0.43729305,0.44119745,0.44119745,0.44510186,0.44900626,0.44900626,0.359205,0.26940376,0.1796025,0.08980125,0.0,0.5700427,1.1400855,1.7101282,2.280171,2.8502135,4.0918136,5.3295093,6.571109,7.8088045,9.050405,8.542832,8.03526,7.5276875,7.0201154,6.5125427,5.3334136,4.154284,2.97125,1.7921207,0.61299115,0.48805028,0.3670138,0.24597734,0.12103647,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14446288,0.21864653,0.28892577,0.3631094,0.59737355,0.8316377,1.0659018,1.3040704,1.5383345,1.2337911,0.93315214,0.62860876,0.3279698,0.023426414,0.023426414,0.019522011,0.015617609,0.015617609,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.06637484,0.12884527,0.19522011,0.26159495,0.3240654,0.30063897,0.28111696,0.25769055,0.23426414,0.21083772,0.22255093,0.23426414,0.24207294,0.25378615,0.26159495,0.7106012,0.62860876,0.5466163,0.46462387,0.38263142,0.30063897,0.26940376,0.23816854,0.21083772,0.1796025,0.14836729,0.14055848,0.13665408,0.12884527,0.12103647,0.113227665,0.1717937,0.22645533,0.28502136,0.3435874,0.39824903,0.39434463,0.39044023,0.38653582,0.37872702,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.14446288,0.26549935,0.38653582,0.5036679,0.62470436,0.6520352,0.679366,0.7066968,0.7340276,0.76135844,0.6715572,0.57785153,0.48414588,0.39434463,0.30063897,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.1639849,0.27330816,0.38653582,0.4997635,0.61299115,0.8355421,1.0580931,1.2806439,1.5031948,1.7257458,1.7101282,1.6945106,1.678893,1.6632754,1.6515622,1.6047094,1.5617609,1.5149081,1.4680552,1.4251068,1.1986516,0.97610056,0.74964523,0.5231899,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.1835069,0.32016098,0.45681506,0.58956474,0.7262188,0.60127795,0.47633708,0.3513962,0.22645533,0.10151446,0.10932326,0.12103647,0.12884527,0.14055848,0.14836729,0.23035973,0.30844778,0.39044023,0.46852827,0.5505207,0.7066968,0.8667773,1.0229534,1.1791295,1.33921,1.4016805,1.4641509,1.5266213,1.5890918,1.6515622,1.5812829,1.5110037,1.4407244,1.3704453,1.3001659,1.1791295,1.0580931,0.94096094,0.8199245,0.698888,0.6910792,0.679366,0.6715572,0.659844,0.6481308,0.58956474,0.5309987,0.46852827,0.40996224,0.3513962,0.8745861,1.4016805,1.9248703,2.4480603,2.9751544,2.7408905,2.5066261,2.2684577,2.0341935,1.7999294,2.0302892,2.260649,2.4910088,2.7213683,2.951728,3.1859922,3.4241607,3.6623292,3.900498,4.138666,4.365122,4.591577,4.8219366,5.0483923,5.2748475,5.036679,4.7985106,4.564246,4.3260775,4.087909,4.029343,3.970777,3.9161155,3.8575494,3.7989833,3.716991,3.6349986,3.5530062,3.4710135,3.3890212,3.4397783,3.49444,3.5451972,3.5959544,3.6506162,4.349504,5.0483923,5.7511845,6.4500723,7.1489606,6.2587566,5.368553,4.478349,3.5881457,2.7018464,3.4866312,4.2753205,5.0640097,5.8487945,6.6374836,6.0713453,5.5013027,4.9351645,4.369026,3.7989833,3.5451972,3.2914112,3.0337205,2.7799344,2.5261483,2.397303,2.2684577,2.1435168,2.0146716,1.8858263,1.8389735,1.7921207,1.7452679,1.698415,1.6515622,1.4836729,1.3157835,1.1478943,0.98000497,0.81211567,0.8160201,0.8160201,0.8199245,0.8238289,0.8238289,1.1557031,1.4914817,1.8233559,2.15523,2.4871042,3.357786,4.2284675,5.099149,5.9659266,6.8366084,7.348085,7.8634663,8.374943,8.886419,9.4018,9.327617,9.253433,9.183154,9.108971,9.0386915,8.367134,7.6955767,7.027924,6.356367,5.688714,5.2201858,4.7516575,4.283129,3.8185053,3.349977,2.9478238,2.5456703,2.1435168,1.7413634,1.33921,1.3157835,1.2962615,1.2767396,1.2572175,1.2376955,1.0580931,0.8823949,0.7066968,0.5270943,0.3513962,0.359205,0.3709182,0.37872702,0.39044023,0.39824903,0.41386664,0.42948425,0.44510186,0.46071947,0.47633708,0.659844,0.8433509,1.0307622,1.2142692,1.4016805,1.3314011,1.261122,1.1908426,1.1205635,1.0502841,1.6827974,2.3153105,2.9478238,3.5803368,4.21285,4.7516575,5.2865605,5.825368,6.364176,6.899079,6.1611466,5.423215,4.689187,3.951255,3.213323,3.8809757,4.552533,5.22409,5.891743,6.5633,7.2856145,8.007929,8.730244,9.452558,10.174872,9.335425,8.495979,7.656533,6.813182,5.9737353,5.9229784,5.8683167,5.8175592,5.7668023,5.7121406,5.8566036,6.001066,6.1494336,6.2938967,6.4383593,5.9542136,5.466163,4.9820175,4.4978714,4.0137253,3.6857557,3.3616903,3.0376248,2.7135596,2.3855898,2.0888553,1.7921207,1.4953861,1.1986516,0.9019169,1.0190489,1.1361811,1.2533131,1.3704453,1.4875772,2.9165885,4.3416953,5.7707067,7.195813,8.624825,10.366188,12.103647,13.845011,15.586374,17.323833,18.167183,19.010534,19.853886,20.693333,21.536682,21.2868,21.036919,20.787037,20.537155,20.287273,19.326792,18.362404,17.40192,16.437534,15.473146,14.543899,13.614651,12.685403,11.756155,10.826907,9.8312845,8.839567,7.8478484,6.8561306,5.8644123,5.758993,5.657479,5.5559645,5.45445,5.349031,4.9156423,4.4861584,4.0527697,3.619381,3.1859922,2.6549935,2.1239948,1.5890918,1.0580931,0.5231899,0.5075723,0.48805028,0.47243267,0.45681506,0.43729305,0.41777104,0.39824903,0.37872702,0.359205,0.3357786,0.26940376,0.20302892,0.13665408,0.06637484,0.0,0.44119745,0.8784905,1.319688,1.7608855,2.1981785,3.853645,5.5091114,7.164578,8.8200445,10.475512,9.749292,9.019169,8.292951,7.5667315,6.8366084,5.6418614,4.4432096,3.2445583,2.0459068,0.8511597,0.679366,0.5114767,0.339683,0.1717937,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.0,0.0,0.0,0.0,0.0,0.14446288,0.28892577,0.43338865,0.58175594,0.7262188,1.1947471,1.6632754,2.135708,2.6042364,3.076669,2.4714866,1.8663043,1.261122,0.6559396,0.05075723,0.046852827,0.039044023,0.03513962,0.031235218,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.05466163,0.10932326,0.1639849,0.21864653,0.27330816,0.25378615,0.23426414,0.21474212,0.19522011,0.1756981,0.1835069,0.19131571,0.19912452,0.20693332,0.21083772,0.47633708,0.42167544,0.3631094,0.30844778,0.25378615,0.19912452,0.1796025,0.16008049,0.14055848,0.12103647,0.10151446,0.093705654,0.08980125,0.08589685,0.078088045,0.07418364,0.14055848,0.21083772,0.27721256,0.3435874,0.41386664,0.42948425,0.44900626,0.46462387,0.48414588,0.4997635,0.5114767,0.5231899,0.5388075,0.5505207,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.21864653,0.39824903,0.57785153,0.75745404,0.93705654,0.97219616,1.0073358,1.0424755,1.077615,1.1127546,0.98000497,0.8472553,0.7145056,0.58175594,0.44900626,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.18741131,0.30063897,0.41386664,0.5231899,0.63641757,0.8667773,1.0932326,1.319688,1.5461433,1.7765031,1.678893,1.5812829,1.4836729,1.3860629,1.2884527,1.2181735,1.1517987,1.0854238,1.0190489,0.94876975,0.80040246,0.6481308,0.4997635,0.3513962,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.13665408,0.12103647,0.10541886,0.08980125,0.07418364,0.27721256,0.48024148,0.6832704,0.8862993,1.0893283,0.9019169,0.7106012,0.5231899,0.3357786,0.14836729,0.14055848,0.12884527,0.12103647,0.10932326,0.10151446,0.21864653,0.339683,0.46071947,0.58175594,0.698888,0.91753453,1.1361811,1.3509232,1.5695697,1.7882162,1.9131571,2.0380979,2.1630387,2.2879796,2.4129205,2.3192148,2.2294137,2.135708,2.0420024,1.9482968,1.7452679,1.5383345,1.3353056,1.1283722,0.92534333,0.8862993,0.8433509,0.80430686,0.76526284,0.7262188,0.6715572,0.62079996,0.5661383,0.5153811,0.46071947,0.8394465,1.2142692,1.5890918,1.9639144,2.338737,2.3348327,2.330928,2.330928,2.3270237,2.3231194,2.631567,2.9400148,3.2484627,3.5569105,3.8614538,4.173806,4.4861584,4.7985106,5.1108627,5.423215,5.833177,6.2431393,6.6531014,7.0630636,7.47693,6.949836,6.426646,5.899552,5.376362,4.8492675,4.794606,4.7399445,4.6852827,4.630621,4.575959,4.369026,4.165997,3.959064,3.7560349,3.5491016,3.5608149,3.5686235,3.5803368,3.5881457,3.5998588,4.1503797,4.7009,5.251421,5.801942,6.348558,5.563773,4.7789884,3.9942036,3.2094188,2.4246337,3.0141985,3.5998588,4.1894236,4.775084,5.3607445,5.2162814,5.0718184,4.927356,4.7828927,4.6384296,4.4041657,4.173806,3.9395418,3.7091823,3.474918,3.2640803,3.0532427,2.8463092,2.6354716,2.4246337,2.3465457,2.2684577,2.194274,2.1161861,2.0380979,1.8038338,1.5734742,1.33921,1.1088502,0.8745861,0.92143893,0.96829176,1.0190489,1.0659018,1.1127546,1.6164225,2.1239948,2.6276627,3.1313305,3.638903,4.493967,5.349031,6.2040954,7.0591593,7.914223,8.125061,8.335898,8.550641,8.761478,8.976221,8.835662,8.695104,8.554545,8.413987,8.273428,7.7307167,7.191909,6.649197,6.1064854,5.563773,5.2162814,4.872694,4.5291066,4.181615,3.8380275,3.3890212,2.9439192,2.494913,2.0459068,1.6008049,1.5461433,1.4914817,1.43682,1.3782539,1.3235924,1.1517987,0.98000497,0.80821127,0.63641757,0.46071947,0.42557985,0.39434463,0.359205,0.3240654,0.28892577,0.3709182,0.45681506,0.5427119,0.62860876,0.7106012,0.92924774,1.1439898,1.358732,1.5734742,1.7882162,1.7218413,1.6515622,1.5851873,1.5188124,1.4485333,2.3816853,3.310933,4.240181,5.169429,6.098676,6.364176,6.6257706,6.8873653,7.1489606,7.4105554,6.6374836,5.8644123,5.087436,4.3143644,3.5373883,4.1308575,4.7243266,5.3138914,5.9073606,6.5008297,7.0903945,7.6799593,8.269524,8.859089,9.448653,8.577971,7.703386,6.832704,5.958118,5.087436,5.1772375,5.267039,5.35684,5.446641,5.5364423,5.6418614,5.74728,5.852699,5.958118,6.0635366,5.74728,5.4310236,5.1186714,4.802415,4.4861584,4.1620927,3.8380275,3.513962,3.1859922,2.8619268,2.533957,2.2059872,1.8819219,1.5539521,1.2259823,1.1947471,1.1635119,1.1361811,1.1049459,1.0737107,2.0459068,3.018103,3.9942036,4.9663997,5.938596,7.223144,8.507692,9.792241,11.076789,12.361338,13.493614,14.625891,15.758167,16.894348,18.026625,18.651329,19.276033,19.900738,20.525442,21.150146,20.298986,19.451733,18.600573,17.749413,16.898252,15.953387,15.008522,14.063657,13.118792,12.173926,11.092407,10.010887,8.929368,7.843944,6.7624245,6.688241,6.617962,6.5437784,6.473499,6.3993154,5.794133,5.1889505,4.5837684,3.978586,3.3734035,2.8463092,2.3153105,1.7843118,1.2533131,0.7262188,0.6676528,0.60908675,0.5544251,0.4958591,0.43729305,0.39434463,0.3513962,0.30844778,0.26940376,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.30844778,0.62079996,0.92924774,1.2415999,1.5500476,3.619381,5.688714,7.7619514,9.8312845,11.900618,10.951848,10.003078,9.058213,8.109444,7.1606736,5.9464045,4.732136,3.5178664,2.3035975,1.0893283,0.8706817,0.6520352,0.43338865,0.21864653,0.0,0.0,0.0,0.0,0.0,0.0,0.113227665,0.22645533,0.3357786,0.44900626,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.05075723,0.10541886,0.15617609,0.21083772,0.26159495,0.21083772,0.15617609,0.10541886,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.21864653,0.43338865,0.6520352,0.8706817,1.0893283,1.7921207,2.4988174,3.2016098,3.9083066,4.6110992,3.7052777,2.7994564,1.8897307,0.98390937,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.046852827,0.08980125,0.13665408,0.1796025,0.22645533,0.20693332,0.19131571,0.1717937,0.15617609,0.13665408,0.14055848,0.14836729,0.15227169,0.15617609,0.1639849,0.23816854,0.21083772,0.1835069,0.15617609,0.12884527,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.046852827,0.046852827,0.042948425,0.039044023,0.039044023,0.113227665,0.19131571,0.26940376,0.3474918,0.42557985,0.46462387,0.5036679,0.5466163,0.58566034,0.62470436,0.6481308,0.6754616,0.698888,0.7262188,0.74964523,0.60127795,0.44900626,0.30063897,0.14836729,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.28892577,0.5309987,0.76916724,1.0112402,1.2494087,1.2923572,1.3353056,1.3782539,1.4212024,1.4641509,1.2884527,1.116659,0.94486535,0.77307165,0.60127795,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.21083772,0.3240654,0.43729305,0.5505207,0.6637484,0.8941081,1.1283722,1.358732,1.5929961,1.8233559,1.6437533,1.4641509,1.2845483,1.1049459,0.92534333,0.8355421,0.74574083,0.6559396,0.5661383,0.47633708,0.39824903,0.3240654,0.24988174,0.1756981,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.1796025,0.16008049,0.14055848,0.12103647,0.10151446,0.3709182,0.64032197,0.9097257,1.1791295,1.4485333,1.1986516,0.94876975,0.698888,0.44900626,0.19912452,0.1717937,0.14055848,0.10932326,0.078088045,0.05075723,0.21083772,0.3709182,0.5309987,0.6910792,0.8511597,1.1283722,1.4055848,1.6827974,1.9600099,2.2372224,2.4246337,2.612045,2.7994564,2.9868677,3.174279,3.0610514,2.9439192,2.8306916,2.7135596,2.6003318,2.3114061,2.018576,1.7296503,1.4407244,1.1517987,1.0815194,1.0112402,0.94096094,0.8706817,0.80040246,0.75354964,0.7106012,0.6637484,0.62079996,0.57394713,0.80040246,1.0268579,1.2494087,1.475864,1.698415,1.9287747,2.1591344,2.3894942,2.619854,2.8502135,3.2367494,3.619381,4.0059166,4.388548,4.775084,5.1616197,5.548156,5.938596,6.3251314,6.7116675,7.3051367,7.898606,8.488171,9.081639,9.675109,8.862993,8.050878,7.238762,6.426646,5.610626,5.559869,5.5091114,5.45445,5.4036927,5.349031,5.0210614,4.6930914,4.369026,4.041056,3.7130866,3.6818514,3.6467118,3.6154766,3.5842414,3.5491016,3.951255,4.349504,4.7516575,5.1499066,5.548156,4.8687897,4.1894236,3.5100577,2.8306916,2.1513257,2.5378613,2.9243972,3.310933,3.7013733,4.087909,4.365122,4.6423345,4.919547,5.196759,5.473972,5.263134,5.056201,4.845363,4.6345253,4.423688,4.1308575,3.8419318,3.5491016,3.2562714,2.9634414,2.854118,2.7486992,2.639376,2.533957,2.4246337,2.1278992,1.8311646,1.53443,1.2337911,0.93705654,1.0307622,1.1205635,1.2142692,1.3079748,1.4016805,2.077142,2.7565079,3.4319696,4.1113358,4.786797,5.6262436,6.46569,7.309041,8.148487,8.987934,8.898132,8.812236,8.726339,8.636538,8.550641,8.343708,8.136774,7.9259367,7.719003,7.5120697,7.098203,6.6843367,6.266566,5.852699,5.4388323,5.2162814,4.9937305,4.7711797,4.548629,4.3260775,3.8341231,3.338264,2.8463092,2.3543546,1.8623998,1.7725986,1.6827974,1.5929961,1.5031948,1.4133936,1.2455044,1.077615,0.9097257,0.7418364,0.57394713,0.4958591,0.41386664,0.3357786,0.25378615,0.1756981,0.3318742,0.48414588,0.64032197,0.79649806,0.94876975,1.1947471,1.4407244,1.6867018,1.9287747,2.174752,2.1083772,2.0459068,1.979532,1.9131571,1.8506867,3.076669,4.3065557,5.532538,6.75852,7.988407,7.9766936,7.9610763,7.9493628,7.9376497,7.9259367,7.113821,6.3017054,5.4856853,4.6735697,3.8614538,4.376835,4.892216,5.407597,5.9229784,6.4383593,6.8951745,7.3519893,7.8088045,8.265619,8.726339,7.8205175,6.914696,6.008875,5.1030536,4.2011366,4.4314966,4.6657605,4.8961205,5.1303844,5.3607445,5.4271193,5.493494,5.5559645,5.6223392,5.688714,5.5442514,5.395884,5.251421,5.1069584,4.9624953,4.6384296,4.3143644,3.9863946,3.6623292,3.338264,2.979059,2.6237583,2.2645533,1.9092526,1.5500476,1.3743496,1.1947471,1.0190489,0.8394465,0.6637484,1.1791295,1.698415,2.2137961,2.7330816,3.2484627,4.0801005,4.911738,5.7394714,6.571109,7.3988423,8.823949,10.2451515,11.666354,13.091461,14.512663,16.011953,17.511244,19.014439,20.51373,22.01302,21.275087,20.537155,19.799223,19.061293,18.32336,17.366781,16.406298,15.445815,14.4853325,13.524849,12.353529,11.178304,10.006983,8.835662,7.6643414,7.621393,7.578445,7.535496,7.492548,7.4495993,6.6726236,5.8956475,5.1186714,4.3416953,3.5608149,3.0337205,2.5066261,1.979532,1.4524376,0.92534333,0.8277333,0.7301232,0.63251317,0.5349031,0.43729305,0.3709182,0.30844778,0.24207294,0.1756981,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.1796025,0.359205,0.5388075,0.71841,0.9019169,3.3851168,5.8683167,8.355421,10.838621,13.325725,12.158309,10.990892,9.823476,8.65606,7.4886436,6.2548523,5.0210614,3.7911747,2.5573835,1.3235924,1.0580931,0.79649806,0.5309987,0.26549935,0.0,0.0,0.0,0.0,0.0,0.0,0.14836729,0.30063897,0.44900626,0.60127795,0.74964523,0.60127795,0.44900626,0.30063897,0.14836729,0.0,0.07027924,0.14055848,0.21083772,0.28111696,0.3513962,0.28111696,0.21083772,0.14055848,0.07027924,0.0,0.0,0.0,0.0,0.0,0.0,0.28892577,0.58175594,0.8706817,1.1596074,1.4485333,2.3894942,3.330455,4.271416,5.2084727,6.1494336,4.939069,3.7287042,2.5183394,1.3118792,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.16008049,0.14446288,0.12884527,0.113227665,0.10151446,0.10151446,0.10541886,0.10932326,0.10932326,0.113227665,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.4997635,0.5622339,0.62470436,0.6871748,0.74964523,0.78868926,0.8238289,0.8628729,0.9019169,0.93705654,0.74964523,0.5622339,0.37482262,0.18741131,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.3631094,0.6637484,0.96438736,1.261122,1.5617609,1.6125181,1.6632754,1.7140326,1.7608855,1.8116426,1.6008049,1.3860629,1.175225,0.96438736,0.74964523,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.23816854,0.3513962,0.46071947,0.57394713,0.6871748,0.92534333,1.1635119,1.4016805,1.6359446,1.8741131,1.6125181,1.3509232,1.0893283,0.8238289,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.22645533,0.19912452,0.1756981,0.14836729,0.12494087,0.46071947,0.80040246,1.1361811,1.475864,1.8116426,1.4992905,1.1869383,0.8745861,0.5622339,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.19912452,0.39824903,0.60127795,0.80040246,0.999527,1.33921,1.6749885,2.0107672,2.35045,2.6862288,2.9361105,3.1859922,3.435874,3.6857557,3.9356375,3.7989833,3.6623292,3.5256753,3.3890212,3.2484627,2.87364,2.4988174,2.1239948,1.7491722,1.3743496,1.2767396,1.175225,1.0737107,0.97610056,0.8745861,0.8394465,0.80040246,0.76135844,0.7262188,0.6871748,0.76135844,0.8394465,0.9136301,0.9878138,1.0619974,1.5266213,1.9873407,2.4519646,2.912684,3.3734035,3.8380275,4.298747,4.7633705,5.22409,5.688714,6.1494336,6.6140575,7.0747766,7.5394006,8.00012,8.773191,9.550168,10.323239,11.100216,11.873287,10.77615,9.675109,8.574067,7.47693,6.375889,6.3251314,6.2743745,6.223617,6.1767645,6.126007,5.6730967,5.22409,4.775084,4.3260775,3.873167,3.7989833,3.7247996,3.6506162,3.5764325,3.4983444,3.7482262,3.998108,4.251894,4.5017757,4.7516575,4.173806,3.5998588,3.0259118,2.4480603,1.8741131,2.0615244,2.2489357,2.436347,2.6237583,2.8111696,3.513962,4.21285,4.911738,5.610626,6.3134184,6.126007,5.938596,5.7511845,5.563773,5.376362,5.001539,4.6267166,4.251894,3.873167,3.4983444,3.3616903,3.2250361,3.0883822,2.951728,2.8111696,2.4480603,2.0888553,1.7257458,1.3626363,0.999527,1.1361811,1.2767396,1.4133936,1.5500476,1.6867018,2.5378613,3.3890212,4.2362766,5.087436,5.938596,6.7624245,7.5862536,8.413987,9.237816,10.061645,9.675109,9.288573,8.898132,8.511597,8.125061,7.8517528,7.57454,7.3012323,7.0240197,6.7507114,6.461786,6.1767645,5.8878384,5.5989127,5.3138914,5.212377,5.1108627,5.0132523,4.911738,4.814128,4.2753205,3.736513,3.2016098,2.6628022,2.1239948,1.999054,1.8741131,1.7491722,1.6242313,1.4992905,1.33921,1.175225,1.0112402,0.8511597,0.6871748,0.5622339,0.43729305,0.31235218,0.18741131,0.062470436,0.28892577,0.5114767,0.737932,0.96438736,1.1869383,1.4641509,1.737459,2.0107672,2.2879796,2.5612879,2.4988174,2.436347,2.3738766,2.3114061,2.2489357,3.775557,5.298274,6.824895,8.351517,9.874233,9.589212,9.300286,9.01136,8.726339,8.437413,7.5862536,6.7389984,5.8878384,5.036679,4.1894236,4.6267166,5.0640097,5.5013027,5.938596,6.375889,6.699954,7.0240197,7.348085,7.676055,8.00012,7.0630636,6.126007,5.1889505,4.251894,3.310933,3.6857557,4.0605783,4.4393053,4.814128,5.1889505,5.212377,5.2358036,5.263134,5.2865605,5.3138914,5.337318,5.3607445,5.388075,5.4115014,5.4388323,5.1108627,4.786797,4.462732,4.138666,3.8106966,3.4241607,3.0376248,2.6510892,2.260649,1.8741131,1.5500476,1.2259823,0.9019169,0.57394713,0.24988174,0.31235218,0.37482262,0.43729305,0.4997635,0.5622339,0.93705654,1.3118792,1.6867018,2.0615244,2.436347,4.1503797,5.860508,7.57454,9.288573,10.998701,13.376482,15.750359,18.124235,20.498112,22.875893,22.251188,21.626484,21.00178,20.37317,19.748466,18.77627,17.800169,16.82407,15.851873,14.875772,13.610746,12.349625,11.088503,9.823476,8.562354,8.550641,8.538928,8.52331,8.511597,8.499884,7.551114,6.5984397,5.64967,4.7009,3.7482262,3.2250361,2.7018464,2.174752,1.6515622,1.1244678,0.9878138,0.8511597,0.7106012,0.57394713,0.43729305,0.3513962,0.26159495,0.1756981,0.08589685,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,3.1508527,6.0518236,8.94889,11.849861,14.750832,13.360865,11.974802,10.588739,9.198771,7.812709,6.5633,5.3138914,4.0605783,2.8111696,1.5617609,1.2494087,0.93705654,0.62470436,0.31235218,0.0,0.0,0.0,0.0,0.0,0.0,0.18741131,0.37482262,0.5622339,0.74964523,0.93705654,0.74964523,0.5622339,0.37482262,0.18741131,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.3513962,0.26159495,0.1756981,0.08589685,0.0,0.0,0.0,0.0,0.0,0.0,0.3631094,0.7262188,1.0893283,1.4485333,1.8116426,2.9868677,4.1620927,5.337318,6.5125427,7.687768,6.1767645,4.661856,3.1508527,1.6359446,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.113227665,0.19912452,0.28892577,0.37482262,0.46071947,0.5192855,0.57394713,0.62860876,0.6832704,0.737932,0.78478485,0.8316377,0.8784905,0.92924774,0.97610056,0.79649806,0.62079996,0.44119745,0.26549935,0.08589685,0.08199245,0.078088045,0.07418364,0.06637484,0.062470436,0.3279698,0.59346914,0.8589685,1.1205635,1.3860629,1.4407244,1.4992905,1.5539521,1.6086137,1.6632754,1.4719596,1.2806439,1.0932326,0.9019169,0.7106012,0.60908675,0.5075723,0.40605783,0.30063897,0.19912452,0.1835069,0.1639849,0.14836729,0.12884527,0.113227665,0.22255093,0.3318742,0.44119745,0.5544251,0.6637484,0.8550641,1.0463798,1.2415999,1.4329157,1.6242313,1.3938715,1.1596074,0.92924774,0.6949836,0.46071947,0.39434463,0.3240654,0.25378615,0.1835069,0.113227665,0.113227665,0.113227665,0.113227665,0.113227665,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.07027924,0.14055848,0.21083772,0.28111696,0.3513962,0.3553006,0.359205,0.3631094,0.3709182,0.37482262,0.59737355,0.8199245,1.0424755,1.2650263,1.4875772,1.261122,1.038571,0.81211567,0.58566034,0.3631094,0.46071947,0.5583295,0.6559396,0.75354964,0.8511597,1.175225,1.4992905,1.8233559,2.1513257,2.475391,3.1313305,3.7911747,4.447114,5.1069584,5.7628975,5.6535745,5.548156,5.4388323,5.3334136,5.22409,5.1069584,4.989826,4.872694,4.755562,4.6384296,4.3338866,4.0332475,3.7287042,3.4280653,3.1235218,2.998581,2.87364,2.7486992,2.6237583,2.4988174,2.5730011,2.6432803,2.717464,2.7916477,2.8619268,2.7682211,2.6706111,2.5769055,2.4831998,2.3855898,2.8619268,3.3343596,3.8067923,4.279225,4.7516575,5.35684,5.958118,6.5633,7.168483,7.773665,7.918128,8.058686,8.203149,8.343708,8.488171,9.120684,9.757101,10.393518,11.0260315,11.66245,10.596548,9.526741,8.460839,7.3910336,6.3251314,6.348558,6.36808,6.3915067,6.4149327,6.4383593,6.028397,5.6223392,5.2162814,4.806319,4.4002614,4.3534083,4.31046,4.263607,4.220659,4.173806,4.6735697,5.173333,5.6730967,6.1767645,6.676528,5.891743,5.1108627,4.3260775,3.5451972,2.7643168,2.8385005,2.912684,2.9868677,3.0610514,3.1391394,3.6076677,4.0761957,4.548629,5.017157,5.4856853,5.677001,5.8683167,6.055728,6.2470436,6.4383593,5.743376,5.0483923,4.3534083,3.6584249,2.9634414,2.9868677,3.0141985,3.0376248,3.0610514,3.0883822,2.8775444,2.6667068,2.455869,2.2489357,2.0380979,1.9404879,1.8428779,1.7452679,1.6476578,1.5500476,2.194274,2.8345962,3.4788225,4.1191444,4.7633705,5.481781,6.196286,6.914696,7.633106,8.351517,8.0040245,7.660437,7.3168497,6.969358,6.6257706,6.5359693,6.446168,6.356367,6.266566,6.1767645,6.0752497,5.9737353,5.8761253,5.774611,5.6730967,5.708236,5.7394714,5.7707067,5.805846,5.8370814,5.2358036,4.6384296,4.037152,3.435874,2.8385005,2.6159496,2.3933985,2.1708477,1.9482968,1.7257458,1.4953861,1.2650263,1.0346665,0.80430686,0.57394713,0.48805028,0.39824903,0.31235218,0.22645533,0.13665408,0.3435874,0.5466163,0.75354964,0.95657855,1.1635119,1.358732,1.5539521,1.7491722,1.9443923,2.135708,2.3855898,2.631567,2.8814487,3.1274261,3.3734035,4.9234514,6.4695945,8.015738,9.565785,11.111929,11.381332,11.6468315,11.916236,12.181735,12.4511385,10.795672,9.140205,7.4847393,5.8292727,4.173806,4.4197836,4.6657605,4.911738,5.153811,5.3997884,5.6379566,5.8761253,6.114294,6.348558,6.5867267,5.8487945,5.1108627,4.376835,3.638903,2.900971,3.5686235,4.240181,4.911738,5.579391,6.250948,6.1884775,6.126007,6.0635366,6.001066,5.938596,5.969831,6.001066,6.036206,6.067441,6.098676,5.7511845,5.4036927,5.056201,4.7087092,4.3612175,4.165997,3.970777,3.7794614,3.5842414,3.3890212,2.9439192,2.5027218,2.0615244,1.6164225,1.175225,1.0346665,0.8941081,0.75354964,0.61689556,0.47633708,0.93315214,1.3899672,1.8467822,2.3035975,2.7643168,3.998108,5.2318993,6.46569,7.703386,8.937177,11.037745,13.138313,15.238882,17.335546,19.436115,19.311174,19.186234,19.061293,18.936352,18.81141,18.424873,18.038338,17.651802,17.261362,16.874826,15.590279,14.30573,13.021181,11.736633,10.44818,10.139732,9.8312845,9.518932,9.2104845,8.898132,8.078208,7.2582836,6.4383593,5.618435,4.7985106,4.2440853,3.6857557,3.1274261,2.5690966,2.0107672,1.7843118,1.5578566,1.3314011,1.1010414,0.8745861,0.7066968,0.5349031,0.3631094,0.19522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,2.6628022,4.950782,7.238762,9.526741,11.810817,10.951848,10.09288,9.2339115,8.371038,7.5120697,6.4305506,5.3529353,4.271416,3.193801,2.1122816,1.7452679,1.3782539,1.0112402,0.6442264,0.27330816,0.26159495,0.24597734,0.23035973,0.21474212,0.19912452,0.339683,0.48024148,0.62079996,0.76135844,0.9019169,0.71841,0.5388075,0.359205,0.1796025,0.0,0.07027924,0.14055848,0.21083772,0.28111696,0.3513962,0.3553006,0.359205,0.3631094,0.3709182,0.37482262,0.49195468,0.60518235,0.71841,0.8355421,0.94876975,1.3860629,1.8233559,2.260649,2.7018464,3.1391394,4.0059166,4.872694,5.7394714,6.606249,7.47693,6.055728,4.6384296,3.2211318,1.8038338,0.38653582,0.32016098,0.25378615,0.1835069,0.11713207,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.10151446,0.093705654,0.08199245,0.07418364,0.062470436,0.06637484,0.07418364,0.078088045,0.08199245,0.08589685,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.13665408,0.22645533,0.31235218,0.39824903,0.48805028,0.5349031,0.58175594,0.62860876,0.679366,0.7262188,0.78088045,0.8394465,0.8980125,0.95657855,1.0112402,0.8433509,0.679366,0.5114767,0.3435874,0.1756981,0.15227169,0.12884527,0.10932326,0.08589685,0.062470436,0.29283017,0.5231899,0.75354964,0.98390937,1.2142692,1.2728351,1.3314011,1.3938715,1.4524376,1.5110037,1.3431144,1.1791295,1.0112402,0.8433509,0.6754616,0.59346914,0.5153811,0.43338865,0.3553006,0.27330816,0.23816854,0.20693332,0.1717937,0.13665408,0.10151446,0.20693332,0.31625658,0.42167544,0.5309987,0.63641757,0.78478485,0.93315214,1.0815194,1.2259823,1.3743496,1.1713207,0.96829176,0.76916724,0.5661383,0.3631094,0.3357786,0.30844778,0.28111696,0.25378615,0.22645533,0.22645533,0.22645533,0.22645533,0.22645533,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.08980125,0.1796025,0.26940376,0.359205,0.44900626,0.48414588,0.5192855,0.5544251,0.58956474,0.62470436,0.7340276,0.8394465,0.94876975,1.0541886,1.1635119,1.0268579,0.8862993,0.74964523,0.61299115,0.47633708,0.71841,0.96438736,1.2103647,1.456342,1.698415,2.1513257,2.6003318,3.049338,3.4983444,3.951255,4.927356,5.903456,6.883461,7.859562,8.835662,8.371038,7.9064145,7.4417906,6.9771667,6.5125427,6.4149327,6.3173227,6.2197127,6.1221027,6.0244927,5.794133,5.563773,5.3334136,5.1069584,4.8765984,4.7243266,4.575959,4.423688,4.2753205,4.126953,4.3065557,4.4900627,4.6735697,4.853172,5.036679,4.7711797,4.50568,4.2440853,3.978586,3.7130866,4.193328,4.677474,5.1616197,5.6418614,6.126007,6.871748,7.621393,8.367134,9.116779,9.86252,9.686822,9.507219,9.331521,9.151918,8.976221,9.468176,9.964035,10.459893,10.955752,11.4516115,10.416945,9.378374,8.343708,7.309041,6.2743745,6.36808,6.46569,6.559396,6.6531014,6.7507114,6.3836975,6.0205884,5.6535745,5.290465,4.9234514,4.911738,4.8961205,4.8805027,4.8648853,4.8492675,5.5989127,6.348558,7.098203,7.8517528,8.601398,7.60968,6.621866,5.630148,4.6384296,3.6506162,3.611572,3.5764325,3.5373883,3.4983444,3.4632049,3.7013733,3.9434462,4.181615,4.423688,4.661856,5.2318993,5.7980375,6.364176,6.9342184,7.5003567,6.4852123,5.4700675,4.454923,3.4397783,2.4246337,2.612045,2.7994564,2.9868677,3.174279,3.3616903,3.3031244,3.2484627,3.1898966,3.1313305,3.076669,2.7408905,2.4090161,2.077142,1.7452679,1.4133936,1.8467822,2.2840753,2.717464,3.1508527,3.5881457,4.1972322,4.806319,5.4193106,6.028397,6.6374836,6.336845,6.0323014,5.7316628,5.4271193,5.12648,5.2201858,5.3138914,5.4115014,5.505207,5.5989127,5.688714,5.774611,5.8644123,5.950309,6.036206,6.2040954,6.36808,6.532065,6.6960497,6.8639393,6.2001905,5.5364423,4.8765984,4.21285,3.5491016,3.2289407,2.9087796,2.5886188,2.2684577,1.9482968,1.6515622,1.3548276,1.0580931,0.76135844,0.46071947,0.41386664,0.3631094,0.31235218,0.26159495,0.21083772,0.39824903,0.58175594,0.76916724,0.95267415,1.1361811,1.2533131,1.3665408,1.4836729,1.5969005,1.7140326,2.2684577,2.8267872,3.3851168,3.9434462,4.5017757,6.0713453,7.6409154,9.2104845,10.780055,12.349625,13.173453,13.993378,14.817206,15.641035,16.46096,14.001186,11.541413,9.081639,6.621866,4.1620927,4.2167544,4.267512,4.318269,4.3729305,4.423688,4.575959,4.7243266,4.8765984,5.024966,5.173333,4.6384296,4.0996222,3.5608149,3.0259118,2.4871042,3.4514916,4.415879,5.3841705,6.348558,7.3129454,7.1606736,7.012306,6.8639393,6.7116675,6.5633,6.602344,6.6413884,6.6843367,6.7233806,6.7624245,6.3915067,6.0205884,5.6535745,5.282656,4.911738,4.911738,4.9078336,4.903929,4.903929,4.900025,4.3416953,3.7794614,3.2211318,2.6588979,2.1005683,1.756981,1.4133936,1.0737107,0.7301232,0.38653582,0.92924774,1.4680552,2.0068626,2.5456703,3.0883822,3.8458362,4.60329,5.3607445,6.1181984,6.8756523,8.699008,10.526268,12.349625,14.176885,16.00024,16.375063,16.749886,17.124708,17.49953,17.874353,18.073479,18.276506,18.475632,18.674755,18.87388,17.565907,16.261835,14.95386,13.645885,12.337912,11.728825,11.123642,10.514555,9.909373,9.300286,8.609207,7.918128,7.230953,6.5398736,5.8487945,5.2592297,4.6696653,4.0801005,3.4905357,2.900971,2.5808098,2.2645533,1.9482968,1.6281357,1.3118792,1.0580931,0.80821127,0.5544251,0.30063897,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,2.174752,3.8497405,5.5247293,7.1997175,8.874706,8.542832,8.210958,7.8790836,7.5433054,7.211431,6.3017054,5.3919797,4.482254,3.5725281,2.6628022,2.241127,1.8194515,1.3938715,0.97219616,0.5505207,0.5192855,0.49195468,0.46071947,0.42948425,0.39824903,0.49195468,0.58566034,0.679366,0.76916724,0.8628729,0.6910792,0.5192855,0.3435874,0.1717937,0.0,0.05075723,0.10541886,0.15617609,0.21083772,0.26159495,0.359205,0.45681506,0.5544251,0.6520352,0.74964523,0.98000497,1.2103647,1.4407244,1.6710842,1.901444,2.4129205,2.9243972,3.435874,3.951255,4.462732,5.0210614,5.5832953,6.141625,6.703859,7.262188,5.938596,4.618908,3.2953155,1.9717231,0.6481308,0.5270943,0.40605783,0.28111696,0.16008049,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.093705654,0.08589685,0.078088045,0.07027924,0.062470436,0.07418364,0.08199245,0.093705654,0.10151446,0.113227665,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.1639849,0.24988174,0.3357786,0.42557985,0.5114767,0.5544251,0.59346914,0.63251317,0.6715572,0.7106012,0.78088045,0.8472553,0.9136301,0.98390937,1.0502841,0.8941081,0.7340276,0.57785153,0.42167544,0.26159495,0.22255093,0.1835069,0.14055848,0.10151446,0.062470436,0.25769055,0.45291066,0.6481308,0.8433509,1.038571,1.1010414,1.1674163,1.2337911,1.2962615,1.3626363,1.2181735,1.0737107,0.92924774,0.78088045,0.63641757,0.58175594,0.5231899,0.46462387,0.40605783,0.3513962,0.29673457,0.24597734,0.19131571,0.14055848,0.08589685,0.19131571,0.29673457,0.40215343,0.5075723,0.61299115,0.7145056,0.8160201,0.92143893,1.0229534,1.1244678,0.95267415,0.78088045,0.60908675,0.43338865,0.26159495,0.27721256,0.29283017,0.30844778,0.3240654,0.3357786,0.3357786,0.3357786,0.3357786,0.3357786,0.3357786,0.26940376,0.20302892,0.13665408,0.06637484,0.0,0.0,0.0,0.0,0.0,0.0,0.10932326,0.21864653,0.3318742,0.44119745,0.5505207,0.61689556,0.679366,0.74574083,0.80821127,0.8745861,0.8667773,0.8589685,0.8511597,0.8433509,0.8394465,0.78868926,0.737932,0.6871748,0.63641757,0.58566034,0.98000497,1.3743496,1.7647898,2.1591344,2.5495746,3.1235218,3.7013733,4.2753205,4.8492675,5.423215,6.7233806,8.019642,9.315904,10.61607,11.912332,11.088503,10.268578,9.444749,8.62092,7.800996,7.7229075,7.6448197,7.5667315,7.4886436,7.4105554,7.2543793,7.098203,6.9381227,6.7819467,6.6257706,6.4500723,6.2743745,6.098676,5.9268827,5.7511845,6.044015,6.336845,6.6257706,6.918601,7.211431,6.7780423,6.3407493,5.9073606,5.473972,5.036679,5.5286336,6.0205884,6.5164475,7.008402,7.5003567,8.39056,9.280765,10.170968,11.061172,11.951375,11.4516115,10.955752,10.455989,9.96013,9.464272,9.815667,10.170968,10.526268,10.881569,11.23687,10.2334385,9.2339115,8.23048,7.2270484,6.223617,6.3915067,6.559396,6.727285,6.8951745,7.0630636,6.7389984,6.4188375,6.094772,5.7707067,5.4505453,5.466163,5.481781,5.493494,5.5091114,5.5247293,6.524256,7.523783,8.52331,9.526741,10.526268,9.327617,8.128965,6.9342184,5.735567,4.5369153,4.388548,4.2362766,4.087909,3.9356375,3.78727,3.7989833,3.8067923,3.8185053,3.8263142,3.8380275,4.7828927,5.727758,6.6726236,7.617489,8.562354,7.2270484,5.891743,4.5564375,3.2211318,1.8858263,2.2372224,2.5886188,2.9361105,3.2875066,3.638903,3.7326086,3.8263142,3.9239242,4.01763,4.1113358,3.5451972,2.979059,2.4090161,1.8428779,1.2767396,1.5031948,1.7296503,1.9561055,2.1864653,2.4129205,2.9165885,3.416352,3.9200199,4.423688,4.9234514,4.6657605,4.4041657,4.1464753,3.8848803,3.6232853,3.9044023,4.185519,4.466636,4.743849,5.024966,5.298274,5.575486,5.8487945,6.126007,6.3993154,6.6960497,6.996689,7.2934237,7.590158,7.8868923,7.1606736,6.4383593,5.7121406,4.985922,4.263607,3.8458362,3.4280653,3.0102942,2.592523,2.174752,1.8116426,1.4446288,1.0815194,0.7145056,0.3513962,0.3357786,0.3240654,0.31235218,0.30063897,0.28892577,0.45291066,0.61689556,0.78088045,0.94876975,1.1127546,1.1478943,1.183034,1.2181735,1.2533131,1.2884527,2.15523,3.0220075,3.8887846,4.755562,5.6262436,7.2192397,8.8083315,10.401327,11.994324,13.58732,14.965574,16.343828,17.718178,19.096432,20.474686,17.210606,13.946525,10.67854,7.4144597,4.1503797,4.009821,3.8692627,3.7287042,3.5881457,3.4514916,3.513962,3.5764325,3.638903,3.7013733,3.7638438,3.4241607,3.0883822,2.7486992,2.4129205,2.0732377,3.3343596,4.5954814,5.8566036,7.113821,8.374943,8.136774,7.898606,7.6643414,7.426173,7.1880045,7.2348576,7.28171,7.328563,7.37932,7.426173,7.0318284,6.6413884,6.2470436,5.8566036,5.462259,5.6535745,5.840986,6.0323014,6.223617,6.4110284,5.735567,5.056201,4.380739,3.7013733,3.0259118,2.4792955,1.9365835,1.3899672,0.8433509,0.30063897,0.92143893,1.5461433,2.1669433,2.7916477,3.4124475,3.6935644,3.970777,4.251894,4.533011,4.814128,6.364176,7.914223,9.464272,11.014318,12.564366,13.438952,14.313539,15.188125,16.062712,16.937298,17.725986,18.51077,19.29946,20.08815,20.876839,19.545437,18.214037,16.88654,15.555139,14.223738,13.32182,12.415999,11.510178,10.604357,9.698535,9.140205,8.581876,8.019642,7.461313,6.899079,6.278279,5.6535745,5.0327744,4.40807,3.78727,3.3812122,2.97125,2.5651922,2.1591344,1.7491722,1.4133936,1.0815194,0.74574083,0.40996224,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.12494087,0.24988174,0.37482262,0.4997635,0.62470436,1.6867018,2.7486992,3.8106966,4.8765984,5.938596,6.133816,6.329036,6.524256,6.715572,6.910792,6.17286,5.4310236,4.6930914,3.951255,3.213323,2.7330816,2.2567444,1.7804074,1.3040704,0.8238289,0.78088045,0.7340276,0.6910792,0.6442264,0.60127795,0.6442264,0.6910792,0.7340276,0.78088045,0.8238289,0.659844,0.4958591,0.3318742,0.1639849,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.3631094,0.5544251,0.74574083,0.93315214,1.1244678,1.4719596,1.815547,2.1591344,2.5066261,2.8502135,3.435874,4.025439,4.6110992,5.2006636,5.786324,6.04011,6.2938967,6.5437784,6.7975645,7.0513506,5.8214636,4.5954814,3.3655949,2.1396124,0.9136301,0.7340276,0.5583295,0.37872702,0.20302892,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.08199245,0.078088045,0.07418364,0.06637484,0.062470436,0.078088045,0.093705654,0.10932326,0.12103647,0.13665408,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.18741131,0.27330816,0.3631094,0.44900626,0.5388075,0.5700427,0.60127795,0.63641757,0.6676528,0.698888,0.77697605,0.8550641,0.93315214,1.0112402,1.0893283,0.94096094,0.79259366,0.6442264,0.4958591,0.3513962,0.29283017,0.23426414,0.1756981,0.12103647,0.062470436,0.22255093,0.38263142,0.5427119,0.7027924,0.8628729,0.93315214,1.0034313,1.0737107,1.1439898,1.2142692,1.0893283,0.96829176,0.8433509,0.7223144,0.60127795,0.5661383,0.5309987,0.4958591,0.46071947,0.42557985,0.3553006,0.28502136,0.21474212,0.14446288,0.07418364,0.1756981,0.28111696,0.38263142,0.48414588,0.58566034,0.6442264,0.7027924,0.76135844,0.8160201,0.8745861,0.7340276,0.58956474,0.44900626,0.30454338,0.1639849,0.21864653,0.27721256,0.3357786,0.39434463,0.44900626,0.44900626,0.44900626,0.44900626,0.44900626,0.44900626,0.359205,0.26940376,0.1796025,0.08980125,0.0,0.0,0.0,0.0,0.0,0.0,0.12884527,0.26159495,0.39044023,0.5192855,0.6481308,0.74574083,0.8394465,0.93315214,1.0307622,1.1244678,1.0034313,0.8784905,0.75745404,0.63641757,0.5114767,0.5505207,0.58566034,0.62470436,0.6637484,0.698888,1.2415999,1.7804074,2.3192148,2.8619268,3.4007344,4.0996222,4.7985106,5.5013027,6.2001905,6.899079,8.519405,10.135828,11.752251,13.368673,14.989,13.805966,12.626837,11.447707,10.268578,9.089449,9.030883,8.972317,8.913751,8.859089,8.800523,8.714626,8.628729,8.546737,8.460839,8.374943,8.175818,7.9766936,7.773665,7.57454,7.375416,7.7775693,8.179723,8.581876,8.98403,9.386183,8.781001,8.175818,7.570636,6.969358,6.364176,6.8639393,7.367607,7.871275,8.371038,8.874706,9.909373,10.940135,11.970898,13.005564,14.036326,13.220306,12.404286,11.584361,10.768341,9.948417,10.163159,10.381805,10.596548,10.81129,11.0260315,10.053836,9.085544,8.113348,7.1450562,6.1767645,6.4149327,6.6531014,6.8951745,7.1333427,7.375416,7.094299,6.813182,6.5359693,6.2548523,5.9737353,6.0205884,6.0635366,6.1103897,6.153338,6.2001905,7.4495993,8.699008,9.948417,11.20173,12.4511385,11.045554,9.639969,8.234385,6.8287997,5.423215,5.1616197,4.900025,4.6384296,4.376835,4.1113358,3.892689,3.6740425,3.4514916,3.232845,3.0141985,4.3338866,5.657479,6.9810715,8.300759,9.6243515,7.968885,6.3134184,4.661856,3.0063896,1.3509232,1.8623998,2.3738766,2.8892577,3.4007344,3.912211,4.1581883,4.40807,4.6540475,4.903929,5.1499066,4.3455997,3.5451972,2.7408905,1.9404879,1.1361811,1.1557031,1.1791295,1.1986516,1.2181735,1.2376955,1.6320401,2.0263848,2.4207294,2.8189783,3.213323,2.9946766,2.77603,2.5612879,2.3426414,2.1239948,2.5886188,3.0532427,3.521771,3.9863946,4.4510183,4.911738,5.376362,5.8370814,6.3017054,6.7624245,7.191909,7.621393,8.050878,8.484266,8.913751,8.125061,7.336372,6.551587,5.7628975,4.9742084,4.4588275,3.9434462,3.4280653,2.9165885,2.4012074,1.9678187,1.53443,1.1010414,0.6715572,0.23816854,0.26159495,0.28892577,0.31235218,0.3357786,0.3631094,0.5075723,0.6520352,0.79649806,0.94096094,1.0893283,1.0424755,0.9956226,0.95267415,0.9058213,0.8628729,2.0380979,3.2172275,4.396357,5.571582,6.7507114,8.36323,9.979652,11.596075,13.208592,14.825015,16.757694,18.690374,20.623053,22.555733,24.48841,20.416119,16.347733,12.2793455,8.207053,4.138666,3.8067923,3.4710135,3.1391394,2.8072653,2.475391,2.4480603,2.4246337,2.4012074,2.3738766,2.35045,2.2137961,2.0732377,1.9365835,1.7999294,1.6632754,3.2172275,4.7711797,6.329036,7.882988,9.43694,9.112875,8.78881,8.460839,8.136774,7.812709,7.8673706,7.9220324,7.9766936,8.031356,8.086017,7.6721506,7.2582836,6.844417,6.426646,6.012779,6.395411,6.7780423,7.1606736,7.5433054,7.9259367,7.1294384,6.336845,5.5403466,4.743849,3.951255,3.2016098,2.455869,1.7062237,0.96048295,0.21083772,0.91753453,1.6242313,2.3270237,3.0337205,3.736513,3.541293,3.3421683,3.1430438,2.9478238,2.7486992,4.025439,5.298274,6.575013,7.8517528,9.124588,10.498938,11.873287,13.251541,14.625891,16.00024,17.37459,18.74894,20.12329,21.501543,22.875893,21.521065,20.170141,18.81922,17.464392,16.113468,14.9109125,13.708356,12.5058,11.303245,10.100689,9.671205,9.24172,8.8083315,8.378847,7.9493628,7.2934237,6.6413884,5.985449,5.3295093,4.6735697,4.1777105,3.6818514,3.182088,2.6862288,2.1864653,1.7686942,1.3509232,0.93315214,0.5192855,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.14836729,0.30063897,0.44900626,0.60127795,0.74964523,1.1986516,1.6515622,2.1005683,2.5495746,2.998581,3.7208953,4.4432096,5.169429,5.891743,6.6140575,6.044015,5.473972,4.903929,4.3338866,3.7638438,3.2289407,2.697942,2.1630387,1.6320401,1.1010414,1.038571,0.98000497,0.92143893,0.8589685,0.80040246,0.79649806,0.79649806,0.79259366,0.78868926,0.78868926,0.62860876,0.47243267,0.31625658,0.15617609,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.3709182,0.6520352,0.93315214,1.2181735,1.4992905,1.9600099,2.4207294,2.8814487,3.338264,3.7989833,4.462732,5.12648,5.786324,6.4500723,7.113821,7.0591593,7.000593,6.9459314,6.89127,6.8366084,5.704332,4.572055,3.4397783,2.3075018,1.175225,0.94096094,0.7106012,0.47633708,0.24597734,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.07418364,0.07027924,0.06637484,0.06637484,0.062470436,0.08199245,0.10151446,0.12103647,0.14055848,0.1639849,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.21083772,0.30063897,0.38653582,0.47633708,0.5622339,0.58566034,0.61299115,0.63641757,0.6637484,0.6871748,0.77307165,0.8628729,0.94876975,1.038571,1.1244678,0.9878138,0.8511597,0.7106012,0.57394713,0.43729305,0.3631094,0.28892577,0.21083772,0.13665408,0.062470436,0.18741131,0.31235218,0.43729305,0.5622339,0.6871748,0.76135844,0.8394465,0.9136301,0.9878138,1.0619974,0.96438736,0.8628729,0.76135844,0.6637484,0.5622339,0.5505207,0.5388075,0.5231899,0.5114767,0.4997635,0.41386664,0.3240654,0.23816854,0.14836729,0.062470436,0.1639849,0.26159495,0.3631094,0.46071947,0.5622339,0.57394713,0.58566034,0.60127795,0.61299115,0.62470436,0.5114767,0.39824903,0.28892577,0.1756981,0.062470436,0.1639849,0.26159495,0.3631094,0.46071947,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.0,0.0,0.0,0.0,0.0,0.14836729,0.30063897,0.44900626,0.60127795,0.74964523,0.8745861,0.999527,1.1244678,1.2494087,1.3743496,1.1361811,0.9019169,0.6637484,0.42557985,0.18741131,0.31235218,0.43729305,0.5622339,0.6871748,0.81211567,1.4992905,2.1864653,2.87364,3.5608149,4.251894,5.0757227,5.899552,6.7233806,7.551114,8.374943,10.311526,12.24811,14.188598,16.125181,18.061766,16.52343,14.989,13.450665,11.912332,10.373997,10.338858,10.299813,10.260769,10.22563,10.186585,10.174872,10.163159,10.151445,10.135828,10.124115,9.901564,9.675109,9.448653,9.226103,8.999647,9.511124,10.0265045,10.537982,11.0494585,11.560935,10.787864,10.010887,9.237816,8.460839,7.687768,8.1992445,8.710721,9.226103,9.737579,10.249056,11.424281,12.599506,13.774731,14.949956,16.125181,14.989,13.848915,12.712734,11.576552,10.436467,10.510651,10.588739,10.662923,10.737106,10.81129,9.874233,8.937177,8.00012,7.0630636,6.126007,6.4383593,6.7507114,7.0630636,7.375416,7.687768,7.4495993,7.211431,6.9732623,6.7389984,6.5008297,6.575013,6.649197,6.7233806,6.801469,6.8756523,8.374943,9.874233,11.373524,12.8767185,14.376009,12.763491,11.150972,9.538455,7.9259367,6.3134184,5.938596,5.563773,5.1889505,4.814128,4.4393053,3.9863946,3.5373883,3.0883822,2.639376,2.1864653,3.8887846,5.5871997,7.2856145,8.987934,10.686349,8.710721,6.7389984,4.7633705,2.787743,0.81211567,1.4875772,2.1630387,2.8385005,3.513962,4.1894236,4.5876727,4.985922,5.388075,5.786324,6.1884775,5.1499066,4.1113358,3.076669,2.0380979,0.999527,0.81211567,0.62470436,0.43729305,0.24988174,0.062470436,0.3513962,0.63641757,0.92534333,1.2142692,1.4992905,1.3235924,1.1517987,0.97610056,0.80040246,0.62470436,1.2767396,1.9248703,2.5769055,3.2250361,3.873167,4.5252023,5.173333,5.825368,6.473499,7.125534,7.687768,8.250002,8.812236,9.37447,9.936704,9.089449,8.238289,7.387129,6.5359693,5.688714,5.0757227,4.462732,3.8497405,3.2367494,2.6237583,2.1239948,1.6242313,1.1244678,0.62470436,0.12494087,0.18741131,0.24988174,0.31235218,0.37482262,0.43729305,0.5622339,0.6871748,0.81211567,0.93705654,1.0619974,0.93705654,0.81211567,0.6871748,0.5622339,0.43729305,1.9248703,3.4124475,4.900025,6.387602,7.8751793,9.511124,11.150972,12.786918,14.426766,16.062712,18.549814,21.036919,23.524023,26.011127,28.498232,23.625538,18.74894,13.8762455,8.999647,4.123049,3.5998588,3.076669,2.5495746,2.0263848,1.4992905,1.3860629,1.2767396,1.1635119,1.0502841,0.93705654,0.999527,1.0619974,1.1244678,1.1869383,1.2494087,3.1000953,4.950782,6.801469,8.648251,10.498938,10.088976,9.675109,9.261242,8.85128,8.437413,8.499884,8.562354,8.624825,8.687295,8.749765,8.312472,7.8751793,7.437886,7.000593,6.5633,7.137247,7.7111945,8.289046,8.862993,9.43694,8.52331,7.6135845,6.699954,5.786324,4.8765984,3.9239242,2.9751544,2.0263848,1.0737107,0.12494087,0.9136301,1.698415,2.4871042,3.2757936,4.0605783,3.3890212,2.7135596,2.0380979,1.3626363,0.6871748,1.6867018,2.6862288,3.6857557,4.689187,5.688714,7.562827,9.43694,11.311053,13.189071,15.063184,17.023193,18.987108,20.951023,22.911032,24.874947,23.500597,22.126247,20.751898,19.373644,17.999294,16.500004,15.000713,13.501423,11.998228,10.498938,10.198298,9.901564,9.600925,9.300286,8.999647,8.312472,7.6252975,6.9381227,6.250948,5.563773,4.9742084,4.388548,3.7989833,3.213323,2.6237583,2.1239948,1.6242313,1.1244678,0.62470436,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.1756981,0.3513962,0.5231899,0.698888,0.8745861,0.7106012,0.5505207,0.38653582,0.22645533,0.062470436,1.3118792,2.5612879,3.8106966,5.0640097,6.3134184,5.911265,5.5130157,5.1108627,4.7126136,4.3143644,3.7247996,3.1391394,2.5495746,1.9639144,1.3743496,1.3001659,1.2259823,1.1517987,1.0737107,0.999527,0.94876975,0.9019169,0.8511597,0.80040246,0.74964523,0.60127795,0.44900626,0.30063897,0.14836729,0.0,0.0,0.0,0.0,0.0,0.0,0.37482262,0.74964523,1.1244678,1.4992905,1.8741131,2.4519646,3.0259118,3.5998588,4.173806,4.7516575,5.4856853,6.223617,6.9615493,7.699481,8.437413,8.074304,7.7111945,7.348085,6.98888,6.6257706,5.5871997,4.548629,3.513962,2.475391,1.43682,1.1517987,0.8628729,0.57394713,0.28892577,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.31235218,0.30063897,0.28892577,0.27330816,0.26159495,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,0.07027924,0.078088045,0.08589685,0.093705654,0.10151446,0.18741131,0.27330816,0.3631094,0.44900626,0.5388075,0.57785153,0.61689556,0.6559396,0.698888,0.737932,0.76916724,0.80430686,0.8355421,0.8667773,0.9019169,0.78868926,0.679366,0.5700427,0.46071947,0.3513962,0.28892577,0.23035973,0.1717937,0.10932326,0.05075723,0.14836729,0.24988174,0.3513962,0.44900626,0.5505207,0.62860876,0.7066968,0.78088045,0.8589685,0.93705654,0.8511597,0.76135844,0.6754616,0.58566034,0.4997635,0.48024148,0.46071947,0.44119745,0.42167544,0.39824903,0.3318742,0.26159495,0.19131571,0.12103647,0.05075723,0.15617609,0.26549935,0.3709182,0.48024148,0.58566034,0.60127795,0.61299115,0.62470436,0.63641757,0.6481308,0.659844,0.6715572,0.679366,0.6910792,0.698888,0.7106012,0.7262188,0.737932,0.74964523,0.76135844,0.7027924,0.6442264,0.58175594,0.5231899,0.46071947,0.3709182,0.27721256,0.1835069,0.093705654,0.0,0.0,0.0,0.0,0.0,0.0,0.12103647,0.23816854,0.359205,0.48024148,0.60127795,0.698888,0.80040246,0.9019169,0.999527,1.1010414,0.9097257,0.71841,0.5309987,0.339683,0.14836729,0.24988174,0.3513962,0.44900626,0.5505207,0.6481308,1.1986516,1.7491722,2.2996929,2.8502135,3.4007344,4.0605783,4.7243266,5.388075,6.0518236,6.7116675,8.441318,10.170968,11.900618,13.634172,15.363823,14.297921,13.232019,12.166118,11.10412,10.0382185,10.194394,10.350571,10.510651,10.666827,10.826907,11.287627,11.748346,12.212971,12.67369,13.138313,12.911859,12.681499,12.455043,12.228588,11.998228,12.228588,12.458947,12.689307,12.919667,13.150026,12.466757,11.779582,11.096312,10.409137,9.725866,9.686822,9.651682,9.612638,9.573594,9.538455,10.331048,11.127546,11.924045,12.716639,13.513136,12.681499,11.845957,11.014318,10.182681,9.351044,9.331521,9.315904,9.296382,9.280765,9.261242,8.609207,7.9532676,7.297328,6.6413884,5.989353,6.1494336,6.3134184,6.473499,6.6374836,6.801469,6.5984397,6.3993154,6.2001905,6.001066,5.7980375,5.8683167,5.9346914,6.001066,6.0713453,6.13772,7.601871,9.066022,10.534078,11.998228,13.462379,12.130978,10.795672,9.464272,8.13287,6.801469,6.551587,6.3017054,6.0518236,5.801942,5.548156,5.0601053,4.5681505,4.0801005,3.5881457,3.1000953,4.4041657,5.708236,7.016211,8.320281,9.6243515,7.918128,6.211904,4.5017757,2.795552,1.0893283,1.5969005,2.1005683,2.6081407,3.1157131,3.6232853,3.9239242,4.224563,4.5252023,4.825841,5.12648,4.271416,3.416352,2.5612879,1.7062237,0.8511597,0.7145056,0.58175594,0.44510186,0.30844778,0.1756981,0.41777104,0.659844,0.9019169,1.1439898,1.3860629,1.2494087,1.1127546,0.97610056,0.8394465,0.698888,1.2103647,1.7218413,2.2294137,2.7408905,3.2484627,3.802888,4.3534083,4.9078336,5.4583545,6.012779,6.461786,6.910792,7.363703,7.812709,8.261715,7.5550184,6.8483214,6.141625,5.4310236,4.7243266,4.2089458,3.6935644,3.1781836,2.6667068,2.1513257,1.7530766,1.358732,0.96438736,0.5700427,0.1756981,0.31625658,0.46071947,0.60127795,0.74574083,0.8862993,0.98390937,1.077615,1.1713207,1.2689307,1.3626363,1.7491722,2.1318035,2.5183394,2.900971,3.2875066,4.185519,5.083532,5.9815445,6.8756523,7.773665,8.94889,10.124115,11.29934,12.4745655,13.64979,15.719124,17.788456,19.861694,21.931028,24.00036,20.209187,16.421915,12.630741,8.839567,5.0483923,4.50568,3.959064,3.416352,2.8697357,2.3231194,2.096664,1.8702087,1.6437533,1.4133936,1.1869383,1.2142692,1.2376955,1.261122,1.2884527,1.3118792,2.7643168,4.2167544,5.6691923,7.1216297,8.574067,8.6131115,8.648251,8.687295,8.726339,8.761478,8.85128,8.937177,9.023073,9.112875,9.198771,9.081639,8.964508,8.847376,8.730244,8.6131115,8.636538,8.65606,8.679486,8.702912,8.726339,8.023546,7.320754,6.617962,5.9151692,5.212377,4.380739,3.5530062,2.7213683,1.893635,1.0619974,1.5812829,2.096664,2.6159496,3.1313305,3.6506162,3.0649557,2.4792955,1.893635,1.3118792,0.7262188,1.5188124,2.3114061,3.1039999,3.8965936,4.689187,6.211904,7.7385254,9.261242,10.787864,12.31058,13.981665,15.652749,17.323833,18.991013,20.662096,19.908546,19.151093,18.397543,17.643993,16.88654,15.992432,15.098324,14.204215,13.306203,12.412095,11.861574,11.311053,10.764437,10.213917,9.663396,8.890324,8.117252,7.3441806,6.571109,5.801942,5.309987,4.8219366,4.3299823,3.8419318,3.349977,2.7643168,2.174752,1.5890918,0.999527,0.41386664,0.5544251,0.698888,0.8394465,0.98390937,1.1244678,1.6242313,2.1200905,2.6159496,3.1157131,3.611572,3.1118085,2.612045,2.1122816,1.6125181,1.1127546,2.4871042,3.8614538,5.2358036,6.6140575,7.988407,7.629202,7.266093,6.9068875,6.547683,6.1884775,5.579391,4.9663997,4.357313,3.7482262,3.1391394,2.7799344,2.4207294,2.0654287,1.7062237,1.3509232,1.2884527,1.2298868,1.1713207,1.1088502,1.0502841,0.8550641,0.659844,0.46462387,0.26940376,0.07418364,0.14055848,0.21083772,0.27721256,0.3435874,0.41386664,0.62860876,0.8472553,1.0659018,1.2806439,1.4992905,2.0732377,2.6432803,3.2172275,3.7911747,4.3612175,4.9468775,5.5286336,6.1103897,6.6921453,7.2739015,6.9732623,6.6687193,6.36808,6.0635366,5.7628975,4.860981,3.9629683,3.0610514,2.1630387,1.261122,1.0112402,0.75745404,0.5036679,0.25378615,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.058566034,0.058566034,0.05466163,0.05075723,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.1756981,0.37482262,0.39824903,0.42557985,0.44900626,0.47633708,0.4997635,0.42557985,0.3513962,0.27330816,0.19912452,0.12494087,0.113227665,0.10541886,0.093705654,0.08589685,0.07418364,0.1639849,0.24988174,0.3357786,0.42557985,0.5114767,0.5661383,0.62079996,0.679366,0.7340276,0.78868926,0.76526284,0.7418364,0.71841,0.698888,0.6754616,0.59346914,0.5114767,0.42557985,0.3435874,0.26159495,0.21864653,0.1717937,0.12884527,0.08199245,0.039044023,0.113227665,0.18741131,0.26159495,0.3357786,0.41386664,0.49195468,0.57394713,0.6520352,0.7340276,0.81211567,0.737932,0.6637484,0.58566034,0.5114767,0.43729305,0.40996224,0.38263142,0.3553006,0.3279698,0.30063897,0.24597734,0.19522011,0.14055848,0.08980125,0.039044023,0.15227169,0.26940376,0.38263142,0.4958591,0.61299115,0.62470436,0.63641757,0.6481308,0.6637484,0.6754616,0.80821127,0.94096094,1.0737107,1.2064602,1.33921,1.261122,1.1869383,1.1127546,1.038571,0.96438736,0.8433509,0.7223144,0.60127795,0.48414588,0.3631094,0.28892577,0.21864653,0.14446288,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.08980125,0.1796025,0.26940376,0.359205,0.44900626,0.5231899,0.60127795,0.6754616,0.74964523,0.8238289,0.6832704,0.5388075,0.39824903,0.25378615,0.113227665,0.18741131,0.26159495,0.3357786,0.41386664,0.48805028,0.9019169,1.3118792,1.7257458,2.135708,2.5495746,3.049338,3.5491016,4.0488653,4.548629,5.0483923,6.571109,8.093826,9.616543,11.139259,12.661977,12.068507,11.478943,10.885473,10.292005,9.698535,10.053836,10.405232,10.756628,11.111929,11.4633255,12.400381,13.337439,14.274494,15.211552,16.148607,15.918248,15.6917925,15.461433,15.231073,15.000713,14.946052,14.895294,14.840633,14.789876,14.739119,14.141745,13.548276,12.950902,12.357433,11.763964,11.174399,10.588739,9.999174,9.413514,8.823949,9.24172,9.655587,10.069453,10.48332,10.901091,10.373997,9.846903,9.315904,8.78881,8.261715,8.152391,8.043069,7.9337454,7.824422,7.7111945,7.3402762,6.969358,6.5945354,6.223617,5.8487945,5.8644123,5.8761253,5.8878384,5.899552,5.911265,5.7511845,5.5871997,5.423215,5.263134,5.099149,5.1616197,5.2201858,5.278752,5.3412223,5.3997884,6.8287997,8.261715,9.690726,11.119738,12.548749,11.498465,10.444276,9.393991,8.339804,7.2856145,7.1606736,7.0357327,6.910792,6.785851,6.66091,6.133816,5.602817,5.0718184,4.5408196,4.0137253,4.9234514,5.833177,6.7429028,7.6526284,8.562354,7.1216297,5.6809053,4.2440853,2.803361,1.3626363,1.7023194,2.0420024,2.3816853,2.7213683,3.0610514,3.2640803,3.4632049,3.6623292,3.8614538,4.0605783,3.3890212,2.717464,2.0459068,1.3743496,0.698888,0.61689556,0.5349031,0.45291066,0.3709182,0.28892577,0.48414588,0.6832704,0.8784905,1.077615,1.2767396,1.175225,1.0737107,0.97610056,0.8745861,0.77307165,1.1439898,1.5149081,1.8858263,2.2567444,2.6237583,3.0805733,3.533484,3.9902992,4.4432096,4.900025,5.2358036,5.575486,5.911265,6.250948,6.5867267,6.0205884,5.4583545,4.892216,4.3260775,3.7638438,3.3460727,2.9283018,2.5105307,2.0927596,1.6749885,1.3860629,1.0932326,0.80430686,0.5153811,0.22645533,0.44900626,0.6715572,0.8941081,1.116659,1.33921,1.4016805,1.4680552,1.53443,1.5969005,1.6632754,2.5573835,3.4514916,4.3455997,5.2436123,6.13772,6.446168,6.7507114,7.0591593,7.367607,7.676055,8.386656,9.101162,9.811763,10.526268,11.23687,12.888432,14.543899,16.195461,17.847023,19.498585,16.796738,14.090988,11.385237,8.679486,5.9737353,5.4115014,4.845363,4.279225,3.7130866,3.1508527,2.8072653,2.463678,2.1239948,1.7804074,1.43682,1.4251068,1.4133936,1.4016805,1.3860629,1.3743496,2.4285383,3.4866312,4.5408196,5.5950084,6.649197,7.137247,7.6252975,8.113348,8.601398,9.089449,9.198771,9.311999,9.425227,9.538455,9.651682,9.850807,10.053836,10.256865,10.459893,10.662923,10.131924,9.600925,9.073831,8.542832,8.011833,7.519879,7.027924,6.5359693,6.044015,5.548156,4.841459,4.1308575,3.4202564,2.7096553,1.999054,2.2489357,2.494913,2.7408905,2.9907722,3.2367494,2.7408905,2.2489357,1.7530766,1.2572175,0.76135844,1.3470187,1.9326792,2.5183394,3.1039999,3.6857557,4.860981,6.036206,7.211431,8.386656,9.561881,10.940135,12.318389,13.696643,15.070992,16.449247,16.316498,16.179844,16.043188,15.9104395,15.773785,15.484859,15.195933,14.903104,14.614178,14.325252,13.524849,12.724447,11.924045,11.123642,10.323239,9.468176,8.609207,7.7541428,6.8951745,6.036206,5.645766,5.251421,4.860981,4.466636,4.0761957,3.4007344,2.7252727,2.0498111,1.3743496,0.698888,1.0112402,1.319688,1.6281357,1.9404879,2.2489357,3.06886,3.8887846,4.7087092,5.5286336,6.348558,5.5130157,4.6735697,3.8380275,2.998581,2.1630387,3.6623292,5.1616197,6.66091,8.164105,9.663396,9.343235,9.023073,8.702912,8.382751,8.062591,7.4300776,6.7975645,6.165051,5.532538,4.900025,4.2597027,3.619381,2.979059,2.338737,1.698415,1.6281357,1.5617609,1.4914817,1.4212024,1.3509232,1.1088502,0.8706817,0.62860876,0.39044023,0.14836729,0.28502136,0.42167544,0.5544251,0.6910792,0.8238289,0.8862993,0.94486535,1.0034313,1.0659018,1.1244678,1.6945106,2.2645533,2.8345962,3.4046388,3.9746814,4.4041657,4.829746,5.2592297,5.6848097,6.114294,5.8683167,5.6262436,5.3841705,5.142098,4.900025,4.138666,3.3734035,2.612045,1.8506867,1.0893283,0.8706817,0.6520352,0.43338865,0.21864653,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.058566034,0.05075723,0.046852827,0.042948425,0.039044023,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.43729305,0.4997635,0.5622339,0.62470436,0.6871748,0.74964523,0.63641757,0.5231899,0.41386664,0.30063897,0.18741131,0.16008049,0.13274968,0.10541886,0.078088045,0.05075723,0.13665408,0.22645533,0.31235218,0.39824903,0.48805028,0.5583295,0.62860876,0.698888,0.76916724,0.8394465,0.76135844,0.6832704,0.60518235,0.5270943,0.44900626,0.39434463,0.339683,0.28502136,0.23035973,0.1756981,0.14446288,0.113227665,0.08589685,0.05466163,0.023426414,0.07418364,0.12494087,0.1756981,0.22645533,0.27330816,0.359205,0.44119745,0.5231899,0.60518235,0.6871748,0.62470436,0.5622339,0.4997635,0.43729305,0.37482262,0.339683,0.30454338,0.26940376,0.23426414,0.19912452,0.1639849,0.12884527,0.093705654,0.058566034,0.023426414,0.14836729,0.26940376,0.39434463,0.5153811,0.63641757,0.6481308,0.6637484,0.6754616,0.6871748,0.698888,0.95657855,1.2103647,1.4641509,1.7218413,1.9756275,1.8116426,1.6515622,1.4875772,1.3235924,1.1635119,0.98390937,0.80430686,0.62079996,0.44119745,0.26159495,0.21083772,0.15617609,0.10541886,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.3513962,0.39824903,0.44900626,0.4997635,0.5505207,0.45681506,0.359205,0.26549935,0.1717937,0.07418364,0.12494087,0.1756981,0.22645533,0.27330816,0.3240654,0.60127795,0.8745861,1.1517987,1.4251068,1.698415,2.0380979,2.3738766,2.7135596,3.049338,3.3890212,4.7009,6.016684,7.3324676,8.648251,9.964035,9.8429985,9.721962,9.600925,9.483793,9.362757,9.909373,10.455989,11.00651,11.553126,12.099743,13.513136,14.92653,16.33602,17.749413,19.162806,18.928543,18.698183,18.463919,18.233559,17.999294,17.663515,17.331642,16.995863,16.660084,16.324306,15.820638,15.313066,14.809398,14.30573,13.798158,12.661977,11.525795,10.38571,9.249529,8.113348,8.148487,8.183627,8.218767,8.253906,8.289046,8.066495,7.843944,7.621393,7.3988423,7.1762915,6.9732623,6.7702336,6.5672045,6.364176,6.1611466,6.0713453,5.9815445,5.891743,5.801942,5.7121406,5.575486,5.4388323,5.298274,5.1616197,5.024966,4.900025,4.775084,4.650143,4.5252023,4.4002614,4.4510183,4.50568,4.5564375,4.6110992,4.661856,6.055728,7.453504,8.847376,10.241247,11.639023,10.865952,10.09288,9.319808,8.546737,7.773665,7.773665,7.773665,7.773665,7.773665,7.773665,7.2036223,6.6335793,6.0635366,5.493494,4.9234514,5.4388323,5.9542136,6.4695945,6.984976,7.5003567,6.329036,5.153811,3.9824903,2.8111696,1.6359446,1.8116426,1.9834363,2.15523,2.3270237,2.4988174,2.6003318,2.7018464,2.7994564,2.900971,2.998581,2.5105307,2.018576,1.5305257,1.038571,0.5505207,0.5192855,0.48805028,0.46071947,0.42948425,0.39824903,0.5544251,0.7066968,0.8589685,1.0112402,1.1635119,1.1010414,1.038571,0.97610056,0.9136301,0.8511597,1.0815194,1.3118792,1.5383345,1.7686942,1.999054,2.358259,2.7135596,3.0727646,3.4280653,3.78727,4.0137253,4.2362766,4.462732,4.689187,4.911738,4.4900627,4.068387,3.6467118,3.2211318,2.7994564,2.4792955,2.1591344,1.8389735,1.5188124,1.1986516,1.0151446,0.8316377,0.6442264,0.46071947,0.27330816,0.57785153,0.8784905,1.183034,1.4836729,1.7882162,1.8233559,1.8584955,1.893635,1.9287747,1.9639144,3.3655949,4.7711797,6.1767645,7.5823493,8.987934,8.706817,8.421796,8.140678,7.8556576,7.57454,7.824422,8.074304,8.324185,8.574067,8.823949,10.061645,11.295436,12.529227,13.766922,15.000713,13.380386,11.760059,10.139732,8.519405,6.899079,6.3134184,5.7316628,5.1460023,4.560342,3.9746814,3.5178664,3.0610514,2.6042364,2.1435168,1.6867018,1.6359446,1.5890918,1.5383345,1.4875772,1.43682,2.096664,2.7526035,3.408543,4.068387,4.7243266,5.661383,6.5984397,7.5394006,8.476458,9.413514,9.550168,9.686822,9.823476,9.964035,10.100689,10.6238785,11.143164,11.666354,12.189544,12.712734,11.631214,10.545791,9.464272,8.382751,7.3012323,7.016211,6.735094,6.453977,6.168956,5.8878384,5.298274,4.7087092,4.1191444,3.5256753,2.9361105,2.9165885,2.893162,2.8697357,2.8463092,2.8267872,2.4207294,2.0146716,1.6086137,1.2064602,0.80040246,1.1791295,1.5539521,1.9326792,2.3114061,2.6862288,3.513962,4.337791,5.1616197,5.989353,6.813182,7.898606,8.98403,10.069453,11.150972,12.236397,12.724447,13.208592,13.692739,14.176885,14.661031,14.977287,15.293544,15.605896,15.9221525,16.238409,15.188125,14.13784,13.087557,12.037272,10.986988,10.046027,9.101162,8.160201,7.2192397,6.2743745,5.9815445,5.6848097,5.388075,5.095245,4.7985106,4.037152,3.2757936,2.5105307,1.7491722,0.9878138,1.4641509,1.9443923,2.4207294,2.8970666,3.3734035,4.5173936,5.661383,6.801469,7.9454584,9.085544,7.914223,6.7389984,5.563773,4.388548,3.213323,4.8375545,6.461786,8.086017,9.714153,11.338385,11.057267,10.77615,10.498938,10.217821,9.936704,9.280765,8.628729,7.9727893,7.3168497,6.66091,5.7394714,4.8180323,3.8965936,2.97125,2.0498111,1.9717231,1.8897307,1.8116426,1.7296503,1.6515622,1.3665408,1.0815194,0.79649806,0.5114767,0.22645533,0.42557985,0.62860876,0.8316377,1.0346665,1.2376955,1.1400855,1.0424755,0.94486535,0.8472553,0.74964523,1.3157835,1.8858263,2.4519646,3.018103,3.5881457,3.8614538,4.1308575,4.4041657,4.677474,4.950782,4.7672753,4.5837684,4.4041657,4.220659,4.037152,3.4124475,2.787743,2.1630387,1.5383345,0.9136301,0.7301232,0.5466163,0.3631094,0.1835069,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05466163,0.046852827,0.039044023,0.031235218,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.4997635,0.60127795,0.698888,0.80040246,0.9019169,0.999527,0.8511597,0.698888,0.5505207,0.39824903,0.24988174,0.20693332,0.16008049,0.113227665,0.07027924,0.023426414,0.113227665,0.19912452,0.28892577,0.37482262,0.46071947,0.5466163,0.63251317,0.71841,0.80430686,0.8862993,0.75354964,0.62079996,0.48805028,0.359205,0.22645533,0.19912452,0.1717937,0.14055848,0.113227665,0.08589685,0.07418364,0.058566034,0.042948425,0.027330816,0.011713207,0.039044023,0.062470436,0.08589685,0.113227665,0.13665408,0.22255093,0.30844778,0.39434463,0.47633708,0.5622339,0.5114767,0.46071947,0.41386664,0.3631094,0.31235218,0.26940376,0.22645533,0.1835069,0.14055848,0.10151446,0.08199245,0.06637484,0.046852827,0.031235218,0.011713207,0.14055848,0.27330816,0.40215343,0.5309987,0.6637484,0.6754616,0.6871748,0.698888,0.7106012,0.7262188,1.1010414,1.4797685,1.8584955,2.233318,2.612045,2.3621633,2.1122816,1.8623998,1.6125181,1.3626363,1.1205635,0.8823949,0.6442264,0.40215343,0.1639849,0.12884527,0.09761006,0.06637484,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.1756981,0.19912452,0.22645533,0.24988174,0.27330816,0.22645533,0.1796025,0.13274968,0.08589685,0.039044023,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.30063897,0.43729305,0.57394713,0.7106012,0.8511597,1.0268579,1.1986516,1.3743496,1.5500476,1.7257458,2.8306916,3.9395418,5.0483923,6.153338,7.262188,7.6135845,7.968885,8.320281,8.671678,9.023073,9.768814,10.510651,11.252487,11.994324,12.73616,14.625891,16.511717,18.401447,20.287273,22.1731,21.938837,21.704573,21.470308,21.236044,21.00178,20.38098,19.764084,19.147188,18.530293,17.913397,17.495626,17.08176,16.667892,16.254026,15.836256,14.149553,12.4628525,10.77615,9.085544,7.3988423,7.055255,6.7116675,6.364176,6.0205884,5.6730967,5.758993,5.840986,5.9229784,6.0049706,6.086963,5.794133,5.4973984,5.2006636,4.9078336,4.6110992,4.806319,4.997635,5.1889505,5.3841705,5.575486,5.2865605,5.001539,4.7126136,4.423688,4.138666,4.0488653,3.9629683,3.873167,3.78727,3.7013733,3.7443218,3.7911747,3.8341231,3.8809757,3.9239242,5.2865605,6.6452928,8.0040245,9.366661,10.725393,10.2334385,9.741484,9.245625,8.75367,8.261715,8.386656,8.511597,8.636538,8.761478,8.886419,8.277332,7.6682463,7.0591593,6.446168,5.8370814,5.958118,6.0791545,6.196286,6.3173227,6.4383593,5.532538,4.6267166,3.7208953,2.8189783,1.9131571,1.9170616,1.9209659,1.9287747,1.9326792,1.9365835,1.9365835,1.9365835,1.9365835,1.9365835,1.9365835,1.6281357,1.3235924,1.0151446,0.7066968,0.39824903,0.42167544,0.44510186,0.46852827,0.48805028,0.5114767,0.62079996,0.7262188,0.8355421,0.94096094,1.0502841,1.0268579,0.999527,0.97610056,0.94876975,0.92534333,1.0151446,1.1049459,1.1947471,1.2845483,1.3743496,1.6359446,1.893635,2.15523,2.416825,2.6745155,2.787743,2.900971,3.0141985,3.1235218,3.2367494,2.9556324,2.67842,2.397303,2.1161861,1.8389735,1.6164225,1.3938715,1.1713207,0.94876975,0.7262188,0.6442264,0.5661383,0.48414588,0.40605783,0.3240654,0.7066968,1.0893283,1.4719596,1.8545911,2.2372224,2.241127,2.2489357,2.25284,2.2567444,2.260649,4.1777105,6.0908675,8.007929,9.921086,11.838148,10.963562,10.09288,9.218294,8.347612,7.47693,7.262188,7.0513506,6.8366084,6.6257706,6.4110284,7.230953,8.046973,8.866898,9.682918,10.498938,9.964035,9.4291315,8.894228,8.359325,7.824422,7.2192397,6.6140575,6.008875,5.4036927,4.7985106,4.2284675,3.6545205,3.0805733,2.5105307,1.9365835,1.8506867,1.7608855,1.6749885,1.5890918,1.4992905,1.7608855,2.018576,2.280171,2.541766,2.7994564,4.1894236,5.575486,6.9615493,8.351517,9.737579,9.901564,10.061645,10.22563,10.38571,10.549695,11.393045,12.236397,13.075843,13.919194,14.762545,13.1266,11.490656,9.858616,8.2226715,6.5867267,6.5164475,6.4422636,6.36808,6.297801,6.223617,5.755089,5.2865605,4.814128,4.3455997,3.873167,3.5842414,3.2914112,2.998581,2.7057507,2.4129205,2.096664,1.7843118,1.4680552,1.1517987,0.8394465,1.0073358,1.1791295,1.3470187,1.5188124,1.6867018,2.1630387,2.639376,3.1118085,3.5881457,4.0605783,4.853172,5.645766,6.4383593,7.230953,8.023546,9.128492,10.2334385,11.338385,12.44333,13.548276,14.469715,15.391153,16.30869,17.230127,18.151566,16.8514,15.551234,14.251068,12.950902,11.650736,10.6238785,9.593117,8.566258,7.5394006,6.5125427,6.3134184,6.1181984,5.919074,5.7238536,5.5247293,4.6735697,3.8263142,2.9751544,2.1239948,1.2767396,1.9209659,2.5651922,3.2094188,3.853645,4.5017757,5.9659266,7.4300776,8.894228,10.358379,11.826434,10.311526,8.800523,7.2856145,5.774611,4.263607,6.012779,7.7619514,9.511124,11.2642,13.013372,12.771299,12.533132,12.291059,12.05289,11.810817,11.135355,10.455989,9.780528,9.101162,8.4257,7.2192397,6.016684,4.8102236,3.6037633,2.4012074,2.3114061,2.2216048,2.1318035,2.0380979,1.9482968,1.620327,1.2884527,0.96048295,0.62860876,0.30063897,0.5700427,0.8394465,1.1088502,1.3782539,1.6515622,1.3938715,1.1400855,0.8862993,0.62860876,0.37482262,0.94096094,1.5031948,2.069333,2.6354716,3.2016098,3.3187418,3.435874,3.5530062,3.6701381,3.78727,3.6662338,3.541293,3.4202564,3.2992198,3.174279,2.6862288,2.1981785,1.7140326,1.2259823,0.737932,0.58956474,0.44119745,0.29673457,0.14836729,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.042948425,0.031235218,0.023426414,0.011713207,0.039044023,0.062470436,0.08589685,0.113227665,0.13665408,0.5622339,0.698888,0.8394465,0.97610056,1.1127546,1.2494087,1.0619974,0.8745861,0.6871748,0.4997635,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.5388075,0.63641757,0.737932,0.8394465,0.93705654,0.74964523,0.5622339,0.37482262,0.18741131,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.39824903,0.3631094,0.3240654,0.28892577,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.13665408,0.27330816,0.41386664,0.5505207,0.6871748,0.698888,0.7106012,0.7262188,0.737932,0.74964523,1.2494087,1.7491722,2.2489357,2.7486992,3.2484627,2.912684,2.5769055,2.2372224,1.901444,1.5617609,1.261122,0.96438736,0.6637484,0.3631094,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.96438736,1.8623998,2.7643168,3.6623292,4.564246,5.388075,6.211904,7.0357327,7.8634663,8.687295,9.6243515,10.561408,11.498465,12.439425,13.376482,15.738646,18.10081,20.462973,22.825136,25.1873,24.949131,24.710962,24.476698,24.23853,24.00036,23.098444,22.200432,21.298513,20.400501,19.498585,19.174519,18.850454,18.526388,18.19842,17.874353,15.637131,13.399908,11.162686,8.925464,6.688241,5.9620223,5.2358036,4.513489,3.78727,3.0610514,3.4514916,3.8380275,4.224563,4.6110992,5.001539,4.6110992,4.224563,3.8380275,3.4514916,3.0610514,3.5373883,4.0137253,4.4861584,4.9624953,5.4388323,5.001539,4.564246,4.123049,3.6857557,3.2484627,3.2016098,3.1508527,3.1000953,3.049338,2.998581,3.0376248,3.076669,3.1118085,3.1508527,3.1859922,4.513489,5.8370814,7.1606736,8.488171,9.811763,9.600925,9.386183,9.175345,8.960603,8.749765,8.999647,9.249529,9.499411,9.749292,9.999174,9.351044,8.699008,8.050878,7.3988423,6.7507114,6.473499,6.2001905,5.9268827,5.64967,5.376362,4.73604,4.0996222,3.4632049,2.8267872,2.1864653,2.0263848,1.8623998,1.698415,1.5383345,1.3743496,1.2767396,1.175225,1.0737107,0.97610056,0.8745861,0.74964523,0.62470436,0.4997635,0.37482262,0.24988174,0.3240654,0.39824903,0.47633708,0.5505207,0.62470436,0.6871748,0.74964523,0.81211567,0.8745861,0.93705654,0.94876975,0.96438736,0.97610056,0.9878138,0.999527,0.94876975,0.9019169,0.8511597,0.80040246,0.74964523,0.9136301,1.0737107,1.2376955,1.4016805,1.5617609,1.5617609,1.5617609,1.5617609,1.5617609,1.5617609,1.4251068,1.2884527,1.1517987,1.0112402,0.8745861,0.74964523,0.62470436,0.4997635,0.37482262,0.24988174,0.27330816,0.30063897,0.3240654,0.3513962,0.37482262,0.8355421,1.3001659,1.7608855,2.2255092,2.6862288,2.6628022,2.639376,2.612045,2.5886188,2.5612879,4.985922,7.4105554,9.839094,12.263727,14.688361,13.224211,11.763964,10.299813,8.835662,7.375416,6.699954,6.0244927,5.349031,4.6735697,3.998108,4.4002614,4.7985106,5.2006636,5.5989127,6.001066,6.551587,7.098203,7.648724,8.1992445,8.749765,8.125061,7.5003567,6.8756523,6.250948,5.6262436,4.939069,4.251894,3.5608149,2.87364,2.1864653,2.0615244,1.9365835,1.8116426,1.6867018,1.5617609,1.4251068,1.2884527,1.1517987,1.0112402,0.8745861,2.7135596,4.548629,6.387602,8.226576,10.061645,10.249056,10.436467,10.6238785,10.81129,10.998701,12.162213,13.325725,14.489237,15.648844,16.812357,14.625891,12.439425,10.249056,8.062591,5.8761253,6.012779,6.1494336,6.2860875,6.426646,6.5633,6.211904,5.8644123,5.5130157,5.1616197,4.814128,4.251894,3.6857557,3.1235218,2.5612879,1.999054,1.7765031,1.5500476,1.3235924,1.1010414,0.8745861,0.8394465,0.80040246,0.76135844,0.7262188,0.6871748,0.81211567,0.93705654,1.0619974,1.1869383,1.3118792,1.8116426,2.3114061,2.8111696,3.310933,3.8106966,5.5364423,7.262188,8.987934,10.71368,12.439425,13.962143,15.488764,17.01148,18.538101,20.06082,18.51077,16.960724,15.410676,13.860628,12.31058,11.20173,10.088976,8.976221,7.8634663,6.7507114,6.649197,6.551587,6.4500723,6.348558,6.250948,5.3138914,4.376835,3.435874,2.4988174,1.5617609,2.3738766,3.1859922,3.998108,4.814128,5.6262436,7.4144597,9.198771,10.986988,12.775204,14.56342,12.712734,10.862047,9.01136,7.1606736,5.3138914,7.1880045,9.062118,10.936231,12.814248,14.688361,14.489237,14.286208,14.087084,13.887959,13.688834,12.986042,12.287154,11.588266,10.889378,10.186585,8.699008,7.211431,5.7238536,4.2362766,2.7486992,2.6510892,2.5495746,2.4480603,2.35045,2.2489357,1.8741131,1.4992905,1.1244678,0.74964523,0.37482262,0.7106012,1.0502841,1.3860629,1.7257458,2.0615244,1.6515622,1.2376955,0.8238289,0.41386664,0.0,0.5622339,1.1244678,1.6867018,2.2489357,2.8111696,2.77603,2.736986,2.7018464,2.6628022,2.6237583,2.5612879,2.4988174,2.436347,2.3738766,2.3114061,1.9639144,1.6125181,1.261122,0.9136301,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.58566034,0.6715572,0.75354964,0.8355421,0.91753453,0.999527,0.8941081,0.78868926,0.6832704,0.58175594,0.47633708,0.42167544,0.3631094,0.30844778,0.25378615,0.19912452,0.23426414,0.26549935,0.29673457,0.3318742,0.3631094,0.48414588,0.60127795,0.7223144,0.8433509,0.96438736,0.79649806,0.62860876,0.46071947,0.29283017,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07027924,0.14055848,0.21083772,0.28111696,0.3513962,0.32016098,0.28892577,0.26159495,0.23035973,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.12103647,0.23816854,0.359205,0.48024148,0.60127795,0.61689556,0.62860876,0.6442264,0.659844,0.6754616,1.0932326,1.5110037,1.9287747,2.3465457,2.7643168,2.533957,2.3035975,2.0732377,1.8428779,1.6125181,1.3626363,1.1127546,0.8628729,0.61299115,0.3631094,0.3513962,0.3357786,0.3240654,0.31235218,0.30063897,0.28892577,0.27330816,0.26159495,0.24988174,0.23816854,0.3240654,0.41386664,0.4997635,0.58566034,0.6754616,0.62470436,0.57394713,0.5231899,0.47633708,0.42557985,0.3709182,0.31625658,0.26159495,0.20693332,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.8511597,1.6047094,2.358259,3.1118085,3.8614538,4.513489,5.165524,5.8214636,6.473499,7.125534,8.011833,8.898132,9.788337,10.674636,11.560935,13.716166,15.867491,18.018816,20.174046,22.325373,22.177006,22.028637,21.884174,21.735807,21.58744,20.482494,19.377548,18.272602,17.167656,16.062712,15.894821,15.726933,15.559043,15.391153,15.223265,13.341343,11.45942,9.577498,7.6955767,5.813655,5.2318993,4.6540475,4.0722914,3.4905357,2.912684,3.2914112,3.6662338,4.044961,4.423688,4.7985106,4.591577,4.380739,4.169902,3.959064,3.7482262,3.951255,4.1503797,4.349504,4.548629,4.7516575,4.322173,3.8965936,3.4671092,3.0415294,2.612045,2.6588979,2.7057507,2.7565079,2.803361,2.8502135,2.9243972,2.9946766,3.06886,3.1391394,3.213323,4.322173,5.4310236,6.5437784,7.6526284,8.761478,8.538928,8.312472,8.086017,7.8634663,7.6370106,7.957172,8.277332,8.597494,8.917655,9.237816,9.0386915,8.843472,8.644346,8.449126,8.250002,7.9064145,7.558923,7.2153354,6.871748,6.524256,6.016684,5.505207,4.9937305,4.4861584,3.9746814,3.9434462,3.9161155,3.8848803,3.853645,3.8263142,3.7716527,3.7208953,3.6662338,3.6154766,3.5608149,3.3538816,3.1469483,2.9400148,2.7330816,2.5261483,2.463678,2.4012074,2.338737,2.2762666,2.2137961,2.1278992,2.0420024,1.9561055,1.8741131,1.7882162,1.737459,1.6867018,1.6359446,1.5890918,1.5383345,1.4485333,1.358732,1.2689307,1.1791295,1.0893283,1.2962615,1.5031948,1.7101282,1.9170616,2.1239948,2.3114061,2.494913,2.67842,2.8658314,3.049338,3.0298162,3.0102942,2.9907722,2.97125,2.951728,2.6823244,2.416825,2.1474214,1.8819219,1.6125181,1.4212024,1.2259823,1.0346665,0.8433509,0.6481308,1.0815194,1.5149081,1.9482968,2.3816853,2.8111696,2.8463092,2.8775444,2.9087796,2.9439192,2.9751544,4.8492675,6.7233806,8.601398,10.475512,12.349625,11.357906,10.366188,9.370565,8.378847,7.387129,6.844417,6.297801,5.7511845,5.2084727,4.661856,4.8687897,5.0718184,5.278752,5.481781,5.688714,6.2040954,6.715572,7.230953,7.746334,8.261715,7.719003,7.1762915,6.6335793,6.0908675,5.548156,4.958591,4.369026,3.7794614,3.1898966,2.6003318,2.5495746,2.4988174,2.4519646,2.4012074,2.35045,2.2918842,2.2294137,2.1708477,2.1083772,2.0498111,3.5256753,5.001539,6.473499,7.9493628,9.425227,9.479889,9.534551,9.589212,9.643873,9.698535,10.932326,12.166118,13.396004,14.629795,15.863586,14.090988,12.322293,10.553599,8.781001,7.012306,7.0240197,7.0357327,7.0513506,7.0630636,7.0747766,6.621866,6.168956,5.716045,5.263134,4.814128,4.3260775,3.8380275,3.349977,2.8619268,2.3738766,2.135708,1.901444,1.6632754,1.4251068,1.1869383,1.0737107,0.96438736,0.8511597,0.737932,0.62470436,0.7262188,0.8238289,0.92534333,1.0268579,1.1244678,1.6164225,2.1044729,2.5964274,3.084478,3.5764325,4.9234514,6.2743745,7.6252975,8.976221,10.323239,11.580457,12.83377,14.090988,15.344301,16.601519,15.605896,14.614178,13.622459,12.630741,11.639023,10.826907,10.018696,9.20658,8.398369,7.5862536,7.445695,7.309041,7.168483,7.027924,6.8873653,5.985449,5.083532,4.181615,3.2757936,2.3738766,3.0883822,3.7989833,4.513489,5.22409,5.938596,7.3168497,8.691199,10.069453,11.447707,12.825961,11.510178,10.194394,8.878611,7.5667315,6.250948,7.47693,8.706817,9.932799,11.158782,12.388668,13.200784,14.016804,14.832824,15.648844,16.46096,14.996809,13.528754,12.0606985,10.592644,9.124588,8.253906,7.3832245,6.5164475,5.645766,4.775084,4.357313,3.9395418,3.521771,3.1039999,2.6862288,2.5534792,2.4207294,2.2918842,2.1591344,2.0263848,2.0146716,2.0068626,1.9951496,1.9834363,1.9756275,2.0068626,2.0341935,2.0654287,2.096664,2.1239948,2.174752,2.2255092,2.2762666,2.3231194,2.3738766,2.3192148,2.2645533,2.2098918,2.15523,2.1005683,2.0615244,2.0263848,1.9873407,1.9482968,1.9131571,1.7921207,1.6710842,1.5539521,1.4329157,1.3118792,1.1400855,0.96829176,0.79649806,0.62079996,0.44900626,0.3670138,0.28502136,0.20302892,0.12103647,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.078088045,0.15617609,0.23426414,0.30844778,0.38653582,0.30844778,0.23426414,0.15617609,0.078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.06637484,0.05466163,0.046852827,0.03513962,0.023426414,0.039044023,0.05466163,0.07027924,0.08589685,0.10151446,0.61299115,0.64032197,0.6676528,0.6949836,0.7223144,0.74964523,0.7262188,0.7066968,0.6832704,0.659844,0.63641757,0.58956474,0.5427119,0.4958591,0.44900626,0.39824903,0.37872702,0.3553006,0.3318742,0.30844778,0.28892577,0.42557985,0.5661383,0.7066968,0.8472553,0.9878138,0.8394465,0.6910792,0.5466163,0.39824903,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10541886,0.15617609,0.21083772,0.26159495,0.23816854,0.21864653,0.19522011,0.1717937,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.20693332,0.30844778,0.40996224,0.5114767,0.5309987,0.5466163,0.5661383,0.58175594,0.60127795,0.93315214,1.2689307,1.6047094,1.9404879,2.2762666,2.1513257,2.0302892,1.9092526,1.7843118,1.6632754,1.4641509,1.261122,1.0619974,0.8628729,0.6637484,0.6481308,0.63641757,0.62470436,0.61299115,0.60127795,0.57394713,0.5505207,0.5231899,0.4997635,0.47633708,0.6481308,0.8238289,0.999527,1.175225,1.3509232,1.2494087,1.1517987,1.0502841,0.94876975,0.8511597,0.7418364,0.62860876,0.5192855,0.40996224,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.13665408,0.7418364,1.3470187,1.9522011,2.5573835,3.1625657,3.6428072,4.123049,4.60329,5.083532,5.563773,6.3993154,7.238762,8.074304,8.913751,9.749292,11.693685,13.634172,15.578565,17.519053,19.463446,19.404879,19.346313,19.29165,19.233086,19.174519,17.866545,16.554665,15.246691,13.934812,12.626837,12.615124,12.603411,12.595602,12.583888,12.576079,11.045554,9.518932,7.9923115,6.46569,4.939069,4.5017757,4.068387,3.631094,3.1977055,2.7643168,3.1313305,3.4983444,3.8653584,4.2323723,4.5993857,4.5681505,4.5369153,4.5017757,4.4705405,4.4393053,4.3612175,4.2870336,4.21285,4.138666,4.0605783,3.6467118,3.2289407,2.8111696,2.3933985,1.9756275,2.1200905,2.2645533,2.4090161,2.5534792,2.7018464,2.8072653,2.9165885,3.0220075,3.1313305,3.2367494,4.1308575,5.02887,5.9229784,6.817086,7.7111945,7.47693,7.238762,7.000593,6.7624245,6.524256,6.914696,7.3051367,7.6955767,8.086017,8.476458,8.730244,8.98403,9.24172,9.495506,9.749292,9.335425,8.921559,8.503788,8.089922,7.676055,7.2934237,6.910792,6.5281606,6.1455293,5.7628975,5.8644123,5.9659266,6.0713453,6.17286,6.2743745,6.27047,6.266566,6.2587566,6.2548523,6.250948,5.958118,5.6691923,5.380266,5.0913405,4.7985106,4.5993857,4.4002614,4.2011366,3.998108,3.7989833,3.5686235,3.3343596,3.1039999,2.8697357,2.639376,2.5261483,2.4129205,2.2996929,2.1864653,2.0732377,1.9443923,1.815547,1.6867018,1.5539521,1.4251068,1.678893,1.9287747,2.182561,2.436347,2.6862288,3.057147,3.4280653,3.7989833,4.165997,4.5369153,4.6345253,4.732136,4.829746,4.927356,5.024966,4.6150036,4.2050414,3.795079,3.3851168,2.9751544,2.5651922,2.15523,1.7452679,1.3353056,0.92534333,1.3274968,1.7296503,2.1318035,2.533957,2.9361105,3.0259118,3.1157131,3.2094188,3.2992198,3.3890212,4.7126136,6.036206,7.363703,8.687295,10.010887,9.491602,8.968412,8.445222,7.9220324,7.3988423,6.984976,6.571109,6.153338,5.7394714,5.3256044,5.3334136,5.3451266,5.35684,5.364649,5.376362,5.8566036,6.336845,6.813182,7.2934237,7.773665,7.3168497,6.8561306,6.395411,5.9346914,5.473972,4.9820175,4.4900627,3.998108,3.506153,3.0141985,3.0376248,3.0610514,3.0883822,3.1118085,3.1391394,3.154757,3.174279,3.1898966,3.2094188,3.2250361,4.337791,5.4505453,6.5633,7.676055,8.78881,8.710721,8.632633,8.554545,8.476458,8.398369,9.702439,11.00651,12.306676,13.610746,14.9109125,13.559989,12.209065,10.8542385,9.503315,8.148487,8.039165,7.9259367,7.812709,7.699481,7.5862536,7.0318284,6.477403,5.9229784,5.368553,4.814128,4.4002614,3.9863946,3.5764325,3.1625657,2.7486992,2.4988174,2.2489357,1.999054,1.7491722,1.4992905,1.3118792,1.1244678,0.93705654,0.74964523,0.5622339,0.63641757,0.7106012,0.78868926,0.8628729,0.93705654,1.4172981,1.8975395,2.377781,2.8580225,3.338264,4.3143644,5.2865605,6.262661,7.238762,8.210958,9.198771,10.182681,11.166591,12.154405,13.138313,12.70102,12.267632,11.834243,11.39695,10.963562,10.455989,9.948417,9.440845,8.933272,8.4257,8.246098,8.066495,7.8868923,7.703386,7.523783,6.657006,5.7902284,4.9234514,4.056674,3.1859922,3.7989833,4.4119744,5.024966,5.6379566,6.250948,7.2192397,8.183627,9.151918,10.120211,11.088503,10.307622,9.526741,8.745861,7.968885,7.1880045,7.7658563,8.347612,8.929368,9.507219,10.088976,11.916236,13.7474,15.578565,17.405825,19.23699,17.003672,14.766449,12.533132,10.295909,8.062591,7.8088045,7.558923,7.3051367,7.0513506,6.801469,6.0635366,5.3295093,4.5954814,3.8614538,3.1235218,3.2367494,3.3460727,3.455396,3.5647192,3.6740425,3.3187418,2.959537,2.6042364,2.2450314,1.8858263,2.358259,2.8306916,3.3031244,3.7794614,4.251894,3.78727,3.3265507,2.8619268,2.4012074,1.9365835,1.8663043,1.7921207,1.7218413,1.6476578,1.5734742,1.5617609,1.5500476,1.5383345,1.5266213,1.5110037,1.6242313,1.7335546,1.8428779,1.9522011,2.0615244,1.8311646,1.5969005,1.3665408,1.1322767,0.9019169,0.7340276,0.5700427,0.40605783,0.23816854,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.15617609,0.30844778,0.46462387,0.62079996,0.77307165,0.62079996,0.46462387,0.30844778,0.15617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.078088045,0.07418364,0.06637484,0.058566034,0.05075723,0.05466163,0.058566034,0.06637484,0.07027924,0.07418364,0.63641757,0.60908675,0.58175594,0.5544251,0.5270943,0.4997635,0.5583295,0.62079996,0.679366,0.7418364,0.80040246,0.76135844,0.71841,0.679366,0.64032197,0.60127795,0.5231899,0.44510186,0.3670138,0.28892577,0.21083772,0.3709182,0.5309987,0.6910792,0.8511597,1.0112402,0.8862993,0.75745404,0.62860876,0.5036679,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.16008049,0.14446288,0.12884527,0.113227665,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.08589685,0.1717937,0.25378615,0.339683,0.42557985,0.44510186,0.46462387,0.48414588,0.5036679,0.5231899,0.77697605,1.0307622,1.2806439,1.53443,1.7882162,1.7725986,1.756981,1.7413634,1.7257458,1.7140326,1.5617609,1.4133936,1.261122,1.1127546,0.96438736,0.94876975,0.93705654,0.92534333,0.9136301,0.9019169,0.8628729,0.8238289,0.78868926,0.74964523,0.7106012,0.97610056,1.2376955,1.4992905,1.7608855,2.0263848,1.8741131,1.7257458,1.5734742,1.4251068,1.2767396,1.1088502,0.94486535,0.78088045,0.61689556,0.44900626,0.359205,0.26940376,0.1796025,0.08980125,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.63251317,1.0893283,1.5461433,2.0068626,2.463678,2.7682211,3.076669,3.3851168,3.6935644,3.998108,4.786797,5.575486,6.364176,7.1489606,7.9376497,9.671205,11.400854,13.134409,14.867964,16.601519,16.632753,16.663988,16.69913,16.730364,16.761599,15.246691,13.731783,12.216875,10.701966,9.187058,9.335425,9.483793,9.628256,9.776623,9.924991,8.75367,7.578445,6.407124,5.2358036,4.0605783,3.7716527,3.4827268,3.193801,2.900971,2.612045,2.97125,3.3265507,3.6857557,4.041056,4.4002614,4.5447245,4.689187,4.83365,4.9781127,5.12648,4.775084,4.423688,4.0761957,3.7247996,3.3734035,2.9673457,2.5612879,2.1513257,1.7452679,1.33921,1.5812829,1.8233559,2.0654287,2.3075018,2.5495746,2.6940374,2.8345962,2.979059,3.1196175,3.2640803,3.9434462,4.6228123,5.3021784,5.9815445,6.66091,6.4110284,6.1611466,5.911265,5.661383,5.4115014,5.872221,6.3329406,6.79366,7.2543793,7.7111945,8.421796,9.128492,9.835189,10.541886,11.248583,10.764437,10.280292,9.796145,9.308095,8.823949,8.570163,8.316377,8.058686,7.8049,7.551114,7.785378,8.019642,8.253906,8.488171,8.726339,8.769287,8.8083315,8.85128,8.894228,8.937177,8.566258,8.191436,7.8205175,7.445695,7.0747766,6.7389984,6.3993154,6.0635366,5.7238536,5.388075,5.009348,4.6267166,4.2479897,3.8692627,3.4866312,3.310933,3.1391394,2.9634414,2.787743,2.612045,2.4441557,2.2723622,2.1005683,1.9326792,1.7608855,2.0615244,2.358259,2.6549935,2.951728,3.2484627,3.8067923,4.3612175,4.9156423,5.4700675,6.0244927,6.239235,6.453977,6.6687193,6.883461,7.098203,6.547683,5.9932575,5.4427366,4.8883114,4.337791,3.7091823,3.0805733,2.455869,1.8272603,1.1986516,1.5734742,1.9443923,2.3192148,2.690133,3.0610514,3.2094188,3.357786,3.506153,3.6506162,3.7989833,4.575959,5.349031,6.126007,6.899079,7.676055,7.621393,7.570636,7.5159745,7.465217,7.4105554,7.1294384,6.844417,6.559396,6.2743745,5.989353,5.801942,5.618435,5.4310236,5.2475166,5.0640097,5.5091114,5.9542136,6.3993154,6.844417,7.2856145,6.910792,6.532065,6.153338,5.7785153,5.3997884,5.0054436,4.6110992,4.2167544,3.8185053,3.4241607,3.5256753,3.6232853,3.7247996,3.8263142,3.9239242,4.0215344,4.11524,4.2089458,4.3065557,4.4002614,5.1499066,5.899552,6.649197,7.3988423,8.148487,7.941554,7.7307167,7.519879,7.309041,7.098203,8.472553,9.846903,11.217348,12.591698,13.962143,13.028991,12.091934,11.158782,10.221725,9.288573,9.050405,8.812236,8.574067,8.335898,8.101635,7.4417906,6.785851,6.126007,5.4700675,4.814128,4.474445,4.138666,3.7989833,3.4632049,3.1235218,2.8619268,2.6003318,2.338737,2.0732377,1.8116426,1.5500476,1.2884527,1.0268579,0.76135844,0.4997635,0.5505207,0.60127795,0.6481308,0.698888,0.74964523,1.2181735,1.6906061,2.1591344,2.631567,3.1000953,3.7013733,4.298747,4.900025,5.5013027,6.098676,6.813182,7.531592,8.246098,8.960603,9.675109,9.796145,9.921086,10.042123,10.163159,10.2881,10.081166,9.878138,9.671205,9.468176,9.261242,9.042596,8.823949,8.601398,8.382751,8.164105,7.328563,6.4969254,5.6652875,4.83365,3.998108,4.513489,5.024966,5.5364423,6.0518236,6.5633,7.1216297,7.676055,8.234385,8.792714,9.351044,9.105066,8.859089,8.6131115,8.371038,8.125061,8.058686,7.988407,7.9220324,7.8556576,7.7892823,10.631687,13.477997,16.324306,19.16671,22.01302,19.010534,16.008049,13.005564,10.003078,7.000593,7.363703,7.7307167,8.093826,8.460839,8.823949,7.773665,6.719476,5.6691923,4.6150036,3.5608149,3.9161155,4.267512,4.618908,4.9742084,5.3256044,4.618908,3.9161155,3.2094188,2.5066261,1.7999294,2.7135596,3.631094,4.5447245,5.4583545,6.375889,5.3997884,4.423688,3.4514916,2.475391,1.4992905,1.4094892,1.319688,1.2298868,1.1400855,1.0502841,1.0619974,1.0737107,1.0893283,1.1010414,1.1127546,1.4524376,1.7921207,2.1318035,2.4714866,2.8111696,2.5183394,2.2294137,1.9365835,1.6437533,1.3509232,1.1010414,0.8550641,0.60908675,0.359205,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.23426414,0.46462387,0.698888,0.92924774,1.1635119,0.92924774,0.698888,0.46462387,0.23426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.093705654,0.08980125,0.08589685,0.078088045,0.07418364,0.07027924,0.06637484,0.058566034,0.05466163,0.05075723,0.6637484,0.58175594,0.4958591,0.41386664,0.3318742,0.24988174,0.39434463,0.5349031,0.679366,0.8199245,0.96438736,0.92924774,0.8980125,0.8667773,0.8316377,0.80040246,0.6676528,0.5349031,0.40215343,0.26940376,0.13665408,0.31625658,0.4958591,0.679366,0.8589685,1.038571,0.92924774,0.8238289,0.7145056,0.60908675,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.078088045,0.07418364,0.06637484,0.058566034,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.06637484,0.13665408,0.20302892,0.26940376,0.3357786,0.359205,0.38263142,0.40605783,0.42557985,0.44900626,0.62079996,0.78868926,0.96048295,1.1283722,1.3001659,1.3938715,1.4836729,1.5773785,1.6710842,1.7608855,1.6632754,1.5617609,1.4641509,1.3626363,1.261122,1.2494087,1.2376955,1.2259823,1.2142692,1.1986516,1.1517987,1.1010414,1.0502841,0.999527,0.94876975,1.3001659,1.6515622,1.999054,2.35045,2.7018464,2.4988174,2.2996929,2.1005683,1.901444,1.698415,1.4797685,1.261122,1.038571,0.8199245,0.60127795,0.48024148,0.359205,0.23816854,0.12103647,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.1639849,0.1756981,0.18741131,0.19912452,0.21083772,0.5231899,0.8316377,1.1439898,1.4524376,1.7608855,1.8975395,2.0341935,2.1669433,2.3035975,2.436347,3.174279,3.912211,4.650143,5.388075,6.126007,7.648724,9.171441,10.694158,12.216875,13.735687,13.860628,13.981665,14.106606,14.227642,14.348679,12.630741,10.9089,9.190963,7.4691215,5.7511845,6.055728,6.3602715,6.6648145,6.969358,7.2739015,6.4578815,5.6418614,4.8219366,4.0059166,3.1859922,3.0415294,2.8970666,2.7526035,2.6081407,2.463678,2.8111696,3.1586614,3.506153,3.853645,4.2011366,4.521298,4.845363,5.169429,5.4895897,5.813655,5.1889505,4.564246,3.9356375,3.310933,2.6862288,2.2918842,1.893635,1.4953861,1.097137,0.698888,1.038571,1.3782539,1.7218413,2.0615244,2.4012074,2.5769055,2.7565079,2.9322062,3.1118085,3.2875066,3.7521305,4.2167544,4.6813784,5.1460023,5.610626,5.349031,5.087436,4.825841,4.564246,4.298747,4.829746,5.3607445,5.891743,6.4188375,6.949836,8.109444,9.269051,10.4286585,11.588266,12.751778,12.193448,11.639023,11.084598,10.530173,9.975748,9.846903,9.721962,9.593117,9.464272,9.339331,9.706344,10.073358,10.4403715,10.807385,11.174399,11.2642,11.354002,11.443803,11.533605,11.623405,11.170495,10.71368,10.260769,9.803954,9.351044,8.874706,8.398369,7.9259367,7.4495993,6.9732623,6.446168,5.919074,5.3919797,4.8648853,4.337791,4.0996222,3.8614538,3.6232853,3.3890212,3.1508527,2.9400148,2.7291772,2.5183394,2.3114061,2.1005683,2.4441557,2.7838387,3.1274261,3.4710135,3.8106966,4.552533,5.2943697,6.0323014,6.774138,7.5120697,7.843944,8.175818,8.511597,8.843472,9.175345,8.480362,7.785378,7.0903945,6.395411,5.700427,4.853172,4.009821,3.1664703,2.3192148,1.475864,1.815547,2.1591344,2.5027218,2.8463092,3.1859922,3.3929255,3.5959544,3.802888,4.0059166,4.21285,4.4393053,4.661856,4.8883114,5.1108627,5.337318,5.755089,6.17286,6.590631,7.008402,7.426173,7.269997,7.113821,6.9615493,6.805373,6.649197,6.27047,5.891743,5.5091114,5.1303844,4.7516575,5.1616197,5.571582,5.9815445,6.3915067,6.801469,6.504734,6.211904,5.9151692,5.618435,5.3256044,5.02887,4.728231,4.4314966,4.134762,3.8380275,4.0137253,4.1894236,4.3612175,4.5369153,4.7126136,4.884407,5.056201,5.2318993,5.4036927,5.575486,5.9620223,6.348558,6.7389984,7.125534,7.5120697,7.168483,6.8287997,6.4852123,6.141625,5.7980375,7.2426662,8.683391,10.128019,11.568744,13.013372,12.494087,11.978706,11.45942,10.944039,10.424754,10.061645,9.698535,9.339331,8.976221,8.6131115,7.8517528,7.094299,6.3329406,5.571582,4.814128,4.548629,4.2870336,4.025439,3.7638438,3.4983444,3.2250361,2.951728,2.6745155,2.4012074,2.1239948,1.7882162,1.4485333,1.1127546,0.77307165,0.43729305,0.46071947,0.48805028,0.5114767,0.5388075,0.5622339,1.0229534,1.4836729,1.9443923,2.4012074,2.8619268,3.0883822,3.310933,3.5373883,3.7638438,3.9863946,4.4314966,4.8765984,5.3217,5.7668023,6.211904,6.89127,7.570636,8.253906,8.933272,9.612638,9.710248,9.807858,9.905469,10.003078,10.100689,9.839094,9.581403,9.319808,9.058213,8.800523,8.0040245,7.2036223,6.407124,5.610626,4.814128,5.22409,5.6379566,6.0518236,6.461786,6.8756523,7.0240197,7.168483,7.3168497,7.465217,7.6135845,7.90251,8.191436,8.484266,8.773191,9.062118,8.347612,7.633106,6.918601,6.2040954,5.4856853,9.347139,13.208592,17.066143,20.927597,24.78905,21.017397,17.245745,13.477997,9.706344,5.938596,6.918601,7.90251,8.886419,9.866425,10.850334,9.479889,8.109444,6.7389984,5.368553,3.998108,4.5954814,5.1889505,5.786324,6.379793,6.9732623,5.9229784,4.8687897,3.8185053,2.7643168,1.7140326,3.06886,4.4275923,5.786324,7.141152,8.499884,7.012306,5.5247293,4.037152,2.5495746,1.0619974,0.95657855,0.8472553,0.7418364,0.63251317,0.5231899,0.5622339,0.60127795,0.63641757,0.6754616,0.7106012,1.2806439,1.8506867,2.4207294,2.9907722,3.5608149,3.2094188,2.8580225,2.5066261,2.1513257,1.7999294,1.4680552,1.1400855,0.80821127,0.48024148,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.30844778,0.62079996,0.92924774,1.2415999,1.5500476,1.2415999,0.92924774,0.62079996,0.30844778,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.10932326,0.10932326,0.10541886,0.10151446,0.10151446,0.08589685,0.07027924,0.05466163,0.039044023,0.023426414,0.6871748,0.5505207,0.41386664,0.27330816,0.13665408,0.0,0.22645533,0.44900626,0.6754616,0.9019169,1.1244678,1.1010414,1.0737107,1.0502841,1.0268579,0.999527,0.81211567,0.62470436,0.43729305,0.24988174,0.062470436,0.26159495,0.46071947,0.6637484,0.8628729,1.0619974,0.97610056,0.8862993,0.80040246,0.7106012,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.27330816,0.30063897,0.3240654,0.3513962,0.37482262,0.46071947,0.5505207,0.63641757,0.7262188,0.81211567,1.0112402,1.2142692,1.4133936,1.6125181,1.8116426,1.7608855,1.7140326,1.6632754,1.6125181,1.5617609,1.5500476,1.5383345,1.5266213,1.5110037,1.4992905,1.43682,1.3743496,1.3118792,1.2494087,1.1869383,1.6242313,2.0615244,2.4988174,2.9361105,3.3734035,3.1235218,2.87364,2.6237583,2.3738766,2.1239948,1.8506867,1.5734742,1.3001659,1.0268579,0.74964523,0.60127795,0.44900626,0.30063897,0.14836729,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,0.41386664,0.57394713,0.737932,0.9019169,1.0619974,1.0268579,0.9878138,0.94876975,0.9136301,0.8745861,1.5617609,2.2489357,2.9361105,3.6232853,4.3143644,5.6262436,6.9381227,8.250002,9.561881,10.87376,11.088503,11.29934,11.514082,11.72492,11.935758,10.010887,8.086017,6.1611466,4.2362766,2.3114061,2.77603,3.2367494,3.7013733,4.1620927,4.6267166,4.1620927,3.7013733,3.2367494,2.77603,2.3114061,2.3114061,2.3114061,2.3114061,2.3114061,2.3114061,2.6510892,2.9868677,3.3265507,3.6623292,3.998108,4.5017757,5.001539,5.5013027,6.001066,6.5008297,5.5989127,4.7009,3.7989833,2.900971,1.999054,1.6125181,1.2259823,0.8355421,0.44900626,0.062470436,0.4997635,0.93705654,1.3743496,1.8116426,2.2489357,2.463678,2.6745155,2.8892577,3.1000953,3.310933,3.5608149,3.8106966,4.0605783,4.3143644,4.564246,4.2870336,4.0137253,3.736513,3.4632049,3.1859922,3.78727,4.388548,4.985922,5.5871997,6.1884775,7.800996,9.413514,11.0260315,12.63855,14.251068,13.626364,13.001659,12.373051,11.748346,11.123642,11.123642,11.123642,11.123642,11.123642,11.123642,11.623405,12.123169,12.626837,13.1266,13.626364,13.763018,13.899672,14.036326,14.176885,14.313539,13.774731,13.235924,12.70102,12.162213,11.623405,11.014318,10.401327,9.788337,9.175345,8.562354,7.8868923,7.211431,6.5359693,5.8644123,5.1889505,4.8883114,4.5876727,4.2870336,3.9863946,3.6857557,3.435874,3.1859922,2.9361105,2.6862288,2.436347,2.8267872,3.213323,3.5998588,3.9863946,4.376835,5.298274,6.223617,7.1489606,8.074304,8.999647,9.448653,9.901564,10.350571,10.799577,11.248583,10.413041,9.573594,8.738052,7.898606,7.0630636,6.001066,4.939069,3.873167,2.8111696,1.7491722,2.0615244,2.3738766,2.6862288,2.998581,3.310933,3.5764325,3.8380275,4.0996222,4.3612175,4.6267166,4.298747,3.9746814,3.6506162,3.3265507,2.998581,3.8887846,4.775084,5.661383,6.551587,7.437886,7.4105554,7.387129,7.363703,7.336372,7.3129454,6.7389984,6.1611466,5.5871997,5.0132523,4.4393053,4.814128,5.1889505,5.563773,5.938596,6.3134184,6.098676,5.8878384,5.6730967,5.462259,5.251421,5.0483923,4.8492675,4.650143,4.4510183,4.251894,4.5017757,4.7516575,5.001539,5.251421,5.5013027,5.7511845,6.001066,6.250948,6.5008297,6.7507114,6.774138,6.801469,6.824895,6.8483214,6.8756523,6.3993154,5.9268827,5.4505453,4.9742084,4.5017757,6.012779,7.523783,9.0386915,10.549695,12.0606985,11.963089,11.861574,11.763964,11.66245,11.560935,11.076789,10.588739,10.100689,9.612638,9.124588,8.261715,7.3988423,6.5359693,5.6730967,4.814128,4.6267166,4.4393053,4.251894,4.0605783,3.873167,3.5881457,3.2992198,3.0141985,2.7252727,2.436347,2.0263848,1.6125181,1.1986516,0.78868926,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.37482262,0.8238289,1.2767396,1.7257458,2.174752,2.6237583,2.475391,2.3231194,2.174752,2.0263848,1.8741131,2.0498111,2.2255092,2.4012074,2.5769055,2.7486992,3.9863946,5.22409,6.461786,7.699481,8.937177,9.339331,9.737579,10.135828,10.537982,10.936231,10.6355915,10.338858,10.0382185,9.737579,9.43694,8.675582,7.914223,7.1489606,6.387602,5.6262436,5.938596,6.250948,6.5633,6.8756523,7.1880045,6.9264097,6.66091,6.3993154,6.13772,5.8761253,6.699954,7.523783,8.351517,9.175345,9.999174,8.636538,7.2739015,5.911265,4.548629,3.1859922,8.062591,12.939189,17.811884,22.688482,27.561176,23.02426,18.487345,13.950429,9.413514,4.8765984,6.473499,8.074304,9.675109,11.275913,12.8767185,11.186112,9.499411,7.812709,6.126007,4.4393053,5.2748475,6.114294,6.949836,7.7892823,8.624825,7.223144,5.825368,4.423688,3.0259118,1.6242313,3.4241607,5.22409,7.0240197,8.823949,10.6238785,8.624825,6.6257706,4.6267166,2.6237583,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,1.1127546,1.9131571,2.7135596,3.513962,4.3143644,3.900498,3.4866312,3.076669,2.6628022,2.2489357,1.8389735,1.4251068,1.0112402,0.60127795,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.38653582,0.77307165,1.1635119,1.5500476,1.9365835,1.5500476,1.1635119,0.77307165,0.38653582,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.5505207,0.44119745,0.3318742,0.21864653,0.10932326,0.0,0.1796025,0.359205,0.5388075,0.71841,0.9019169,0.8784905,0.8589685,0.8394465,0.8199245,0.80040246,0.6481308,0.4997635,0.3513962,0.19912452,0.05075723,0.21083772,0.3709182,0.5309987,0.6910792,0.8511597,0.79649806,0.7418364,0.6832704,0.62860876,0.57394713,0.5309987,0.48414588,0.44119745,0.39434463,0.3513962,0.3435874,0.3357786,0.3279698,0.32016098,0.31235218,0.29283017,0.27330816,0.25378615,0.23426414,0.21083772,0.19131571,0.1717937,0.15227169,0.13274968,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.19912452,0.25769055,0.31625658,0.37872702,0.43729305,0.43729305,0.43729305,0.43729305,0.43729305,0.43729305,0.5505207,0.6637484,0.77307165,0.8862993,0.999527,1.2142692,1.4251068,1.6359446,1.8506867,2.0615244,1.999054,1.9365835,1.8741131,1.8116426,1.7491722,1.7335546,1.7218413,1.7062237,1.6906061,1.6749885,1.6125181,1.5500476,1.4875772,1.4251068,1.3626363,1.8194515,2.2762666,2.7330816,3.193801,3.6506162,3.521771,3.3890212,3.260176,3.1313305,2.998581,2.7330816,2.4714866,2.2059872,1.9404879,1.6749885,1.6437533,1.6086137,1.5773785,1.5461433,1.5110037,1.4602464,1.4055848,1.3548276,1.3040704,1.2494087,1.3157835,1.3782539,1.4446288,1.5110037,1.5734742,1.7647898,1.9561055,2.1435168,2.3348327,2.5261483,2.3035975,2.084951,1.8663043,1.6437533,1.4251068,1.8897307,2.3543546,2.8189783,3.2836022,3.7482262,4.786797,5.8214636,6.8561306,7.890797,8.925464,9.128492,9.331521,9.530646,9.733675,9.936704,8.503788,7.066968,5.6340523,4.1972322,2.7643168,3.0102942,3.2562714,3.506153,3.7521305,3.998108,3.611572,3.2211318,2.8306916,2.4402514,2.0498111,2.1513257,2.2567444,2.358259,2.4597735,2.5612879,2.8892577,3.2172275,3.5451972,3.873167,4.2011366,4.5291066,4.853172,5.181142,5.5091114,5.8370814,5.138193,4.4432096,3.7443218,3.049338,2.35045,2.0068626,1.6593709,1.3157835,0.96829176,0.62470436,1.2142692,1.7999294,2.3855898,2.9751544,3.5608149,3.959064,4.3534083,4.747753,5.142098,5.5364423,5.6340523,5.7316628,5.8292727,5.9268827,6.0244927,5.364649,4.704805,4.044961,3.3851168,2.7252727,3.240654,3.7599394,4.279225,4.794606,5.3138914,6.6726236,8.031356,9.393991,10.752724,12.111456,11.775677,11.443803,11.108025,10.772245,10.436467,10.479416,10.522364,10.565312,10.608261,10.651209,11.0260315,11.404759,11.783486,12.158309,12.537036,12.67369,12.806439,12.943093,13.075843,13.212498,12.708829,12.209065,11.705398,11.20173,10.698062,10.22563,9.753197,9.280765,8.8083315,8.335898,7.800996,7.262188,6.7233806,6.1884775,5.64967,5.2475166,4.845363,4.4432096,4.041056,3.638903,3.5451972,3.4514916,3.3616903,3.2679846,3.174279,3.49444,3.814601,4.134762,4.454923,4.775084,5.6965227,6.6140575,7.535496,8.456935,9.37447,9.589212,9.803954,10.018696,10.2334385,10.44818,9.655587,8.866898,8.074304,7.28171,6.4891167,5.6652875,4.841459,4.0215344,3.1977055,2.3738766,2.5808098,2.7916477,2.998581,3.2055142,3.4124475,3.513962,3.619381,3.7208953,3.8224099,3.9239242,3.7013733,3.474918,3.2484627,3.0259118,2.7994564,3.5959544,4.388548,5.185046,5.9815445,6.774138,6.9615493,7.1450562,7.328563,7.5159745,7.699481,7.2270484,6.754616,6.282183,5.8097506,5.337318,5.5247293,5.7121406,5.899552,6.086963,6.2743745,6.133816,5.989353,5.8487945,5.704332,5.563773,5.3841705,5.2006636,5.0210614,4.841459,4.661856,4.8219366,4.9820175,5.142098,5.3021784,5.462259,5.8487945,6.239235,6.6257706,7.012306,7.3988423,7.4183645,7.4417906,7.461313,7.480835,7.5003567,6.9342184,6.36808,5.805846,5.239708,4.6735697,6.0713453,7.465217,8.859089,10.256865,11.650736,11.4516115,11.248583,11.0494585,10.850334,10.651209,10.22563,9.803954,9.382278,8.960603,8.538928,8.289046,8.039165,7.7892823,7.5394006,7.2856145,6.453977,5.6223392,4.7907014,3.959064,3.1235218,3.0063896,2.8853533,2.7643168,2.6432803,2.5261483,2.416825,2.3114061,2.2020829,2.096664,1.9873407,1.9170616,1.8467822,1.7765031,1.7062237,1.6359446,1.756981,1.8780174,1.999054,2.1161861,2.2372224,2.2567444,2.2723622,2.2918842,2.3075018,2.3231194,2.4285383,2.5300527,2.631567,2.7330816,2.8385005,3.8809757,4.927356,5.9737353,7.016211,8.062591,9.0152645,9.967939,10.920613,11.873287,12.825961,12.111456,11.400854,10.686349,9.975748,9.261242,8.839567,8.4178915,7.996216,7.570636,7.1489606,7.2543793,7.3597984,7.465217,7.570636,7.676055,7.519879,7.363703,7.211431,7.055255,6.899079,7.211431,7.519879,7.8283267,8.140678,8.449126,7.570636,6.688241,5.8097506,4.93126,4.0488653,7.734621,11.416472,15.098324,18.780174,22.462027,19.174519,15.8870125,12.599506,9.311999,6.0244927,7.1177254,8.210958,9.304191,10.393518,11.486752,10.350571,9.21439,8.074304,6.9381227,5.801942,6.329036,6.8561306,7.3832245,7.910319,8.437413,7.4574084,6.477403,5.4973984,4.5173936,3.5373883,4.661856,5.786324,6.910792,8.039165,9.163632,7.4417906,5.7238536,4.0020123,2.2840753,0.5622339,0.4997635,0.43729305,0.37482262,0.31235218,0.24988174,0.3240654,0.39824903,0.47633708,0.5505207,0.62470436,1.2259823,1.8233559,2.4246337,3.0259118,3.6232853,3.416352,3.2094188,3.0024853,2.795552,2.5886188,2.2684577,1.9522011,1.6359446,1.3157835,0.999527,0.8862993,0.76916724,0.6559396,0.5388075,0.42557985,0.6715572,0.9136301,1.1596074,1.4055848,1.6515622,1.33921,1.0268579,0.7106012,0.39824903,0.08589685,0.14836729,0.20693332,0.26940376,0.3279698,0.38653582,0.45681506,0.5231899,0.58956474,0.6559396,0.7262188,0.58175594,0.43338865,0.28892577,0.14446288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.113227665,0.113227665,0.113227665,0.113227665,0.113227665,0.093705654,0.078088045,0.058566034,0.042948425,0.023426414,0.41386664,0.3318742,0.24597734,0.1639849,0.08199245,0.0,0.13665408,0.26940376,0.40605783,0.5388075,0.6754616,0.659844,0.6442264,0.62860876,0.61689556,0.60127795,0.48805028,0.37482262,0.26159495,0.14836729,0.039044023,0.15617609,0.27721256,0.39824903,0.5192855,0.63641757,0.61689556,0.59346914,0.5700427,0.5466163,0.5231899,0.5583295,0.59346914,0.62860876,0.6637484,0.698888,0.6832704,0.6715572,0.6559396,0.64032197,0.62470436,0.58566034,0.5466163,0.5036679,0.46462387,0.42557985,0.38653582,0.3435874,0.30454338,0.26549935,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.05466163,0.10932326,0.1639849,0.21864653,0.27330816,0.3435874,0.41386664,0.48414588,0.5544251,0.62470436,0.60127795,0.57394713,0.5505207,0.5231899,0.4997635,0.63641757,0.77307165,0.9136301,1.0502841,1.1869383,1.4133936,1.6359446,1.8623998,2.0888553,2.3114061,2.2372224,2.1630387,2.0888553,2.0107672,1.9365835,1.9209659,1.901444,1.8858263,1.8663043,1.8506867,1.7882162,1.7257458,1.6632754,1.6008049,1.5383345,2.0146716,2.4910088,2.97125,3.4475873,3.9239242,3.9161155,3.9044023,3.8965936,3.8848803,3.873167,3.619381,3.3655949,3.1118085,2.854118,2.6003318,2.6862288,2.7682211,2.854118,2.9400148,3.0259118,2.8814487,2.7408905,2.5964274,2.455869,2.3114061,2.4285383,2.5456703,2.6667068,2.7838387,2.900971,3.1157131,3.3343596,3.5530062,3.7716527,3.9863946,3.5842414,3.182088,2.7799344,2.377781,1.9756275,2.2177005,2.4597735,2.7018464,2.9439192,3.1859922,3.9434462,4.7009,5.4583545,6.2158084,6.9732623,7.168483,7.3597984,7.551114,7.746334,7.9376497,6.9927845,6.0479193,5.1030536,4.1581883,3.213323,3.2445583,3.2757936,3.310933,3.3421683,3.3734035,3.057147,2.7408905,2.4207294,2.1044729,1.7882162,1.9912452,2.1981785,2.4012074,2.6081407,2.8111696,3.1313305,3.4475873,3.7638438,4.084005,4.4002614,4.5564375,4.7087092,4.8648853,5.0210614,5.173333,4.6813784,4.185519,3.68966,3.193801,2.7018464,2.397303,2.096664,1.7921207,1.4914817,1.1869383,1.9248703,2.6628022,3.4007344,4.138666,4.8765984,5.45445,6.028397,6.606249,7.1841,7.7619514,7.70729,7.6526284,7.5979667,7.5433054,7.4886436,6.4422636,5.395884,4.3534083,3.3070288,2.260649,2.697942,3.1313305,3.5686235,4.0020123,4.4393053,5.5442514,6.6531014,7.7619514,8.866898,9.975748,9.928895,9.885946,9.839094,9.796145,9.749292,9.835189,9.921086,10.003078,10.088976,10.174872,10.4286585,10.686349,10.940135,11.193921,11.4516115,11.584361,11.713207,11.845957,11.978706,12.111456,11.6468315,11.178304,10.709775,10.241247,9.776623,9.440845,9.108971,8.777096,8.445222,8.113348,7.7111945,7.3129454,6.910792,6.5125427,6.114294,5.606722,5.1030536,4.5993857,4.0918136,3.5881457,3.6506162,3.716991,3.7833657,3.8458362,3.912211,4.165997,4.415879,4.6696653,4.9234514,5.173333,6.0908675,7.0044975,7.918128,8.835662,9.749292,9.729771,9.710248,9.690726,9.671205,9.651682,8.902037,8.156297,7.406651,6.66091,5.911265,5.3295093,4.747753,4.165997,3.5842414,2.998581,3.1039999,3.2055142,3.3070288,3.408543,3.513962,3.455396,3.39683,3.338264,3.2836022,3.2250361,3.1000953,2.9751544,2.8502135,2.7252727,2.6003318,3.3031244,4.0059166,4.7087092,5.4115014,6.114294,6.5086384,6.902983,7.297328,7.6916723,8.086017,7.719003,7.348085,6.9771667,6.606249,6.239235,6.239235,6.239235,6.239235,6.239235,6.239235,6.165051,6.0908675,6.0205884,5.9464045,5.8761253,5.716045,5.5559645,5.395884,5.2358036,5.0757227,5.1460023,5.2162814,5.2865605,5.35684,5.423215,5.950309,6.473499,7.000593,7.523783,8.050878,8.066495,8.078208,8.093826,8.109444,8.125061,7.4691215,6.813182,6.1611466,5.505207,4.8492675,6.126007,7.406651,8.683391,9.96013,11.23687,10.936231,10.6355915,10.338858,10.0382185,9.737579,9.378374,9.023073,8.663869,8.308568,7.9493628,8.312472,8.675582,9.0386915,9.4018,9.761005,8.285142,6.8092775,5.3295093,3.853645,2.3738766,2.4207294,2.4714866,2.5183394,2.5651922,2.612045,2.8111696,3.0063896,3.2055142,3.4007344,3.5998588,3.4593005,3.3187418,3.1781836,3.0415294,2.900971,2.690133,2.4792955,2.2684577,2.0615244,1.8506867,2.0341935,2.2216048,2.4051118,2.5886188,2.77603,2.803361,2.8345962,2.8658314,2.893162,2.9243972,3.7794614,4.630621,5.481781,6.336845,7.1880045,8.691199,10.198298,11.701493,13.208592,14.711788,13.58732,12.4628525,11.338385,10.213917,9.089449,9.0035515,8.921559,8.839567,8.757574,8.675582,8.574067,8.468649,8.367134,8.265619,8.164105,8.113348,8.066495,8.019642,7.9727893,7.9259367,7.719003,7.5159745,7.309041,7.1060123,6.899079,6.5008297,6.1064854,5.708236,5.309987,4.911738,7.4027467,9.893755,12.380859,14.871868,17.362877,15.324779,13.286681,11.248583,9.21439,7.1762915,7.7619514,8.343708,8.929368,9.515028,10.100689,9.511124,8.925464,8.335898,7.7502384,7.1606736,7.37932,7.5979667,7.816613,8.031356,8.250002,7.6916723,7.1294384,6.571109,6.008875,5.4505453,5.899552,6.348558,6.801469,7.250475,7.699481,6.2587566,4.8219366,3.3812122,1.9404879,0.4997635,0.4997635,0.4997635,0.4997635,0.4997635,0.4997635,0.58566034,0.6754616,0.76135844,0.8511597,0.93705654,1.33921,1.737459,2.135708,2.5378613,2.9361105,2.9361105,2.9322062,2.9283018,2.9283018,2.9243972,2.7018464,2.4792955,2.2567444,2.0341935,1.8116426,1.620327,1.4290112,1.2337911,1.0424755,0.8511597,0.95267415,1.0541886,1.1557031,1.261122,1.3626363,1.1244678,0.8862993,0.6481308,0.41386664,0.1756981,0.29673457,0.41386664,0.5349031,0.6559396,0.77307165,0.9097257,1.0463798,1.1791295,1.3157835,1.4485333,1.1596074,0.8706817,0.58175594,0.28892577,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.27330816,0.21864653,0.1639849,0.10932326,0.05466163,0.0,0.08980125,0.1796025,0.26940376,0.359205,0.44900626,0.44119745,0.42948425,0.42167544,0.40996224,0.39824903,0.3240654,0.24988174,0.1756981,0.10151446,0.023426414,0.10541886,0.1835069,0.26549935,0.3435874,0.42557985,0.43338865,0.44510186,0.45681506,0.46462387,0.47633708,0.58956474,0.7066968,0.8199245,0.93315214,1.0502841,1.0268579,1.0034313,0.98390937,0.96048295,0.93705654,0.8784905,0.8160201,0.75745404,0.698888,0.63641757,0.57785153,0.5192855,0.45681506,0.39824903,0.3357786,0.26940376,0.20302892,0.13665408,0.06637484,0.0,0.0,0.0,0.0,0.0,0.0,0.08199245,0.1639849,0.24597734,0.3318742,0.41386664,0.49195468,0.57394713,0.6520352,0.7340276,0.81211567,0.76135844,0.7106012,0.6637484,0.61299115,0.5622339,0.7262188,0.8862993,1.0502841,1.2142692,1.3743496,1.6125181,1.8506867,2.0888553,2.3231194,2.5612879,2.475391,2.3855898,2.2996929,2.2137961,2.1239948,2.1044729,2.084951,2.0654287,2.0459068,2.0263848,1.9639144,1.901444,1.8389735,1.7765031,1.7140326,2.2098918,2.7057507,3.2055142,3.7013733,4.2011366,4.31046,4.4197836,4.5291066,4.6384296,4.7516575,4.50568,4.2597027,4.0137253,3.7716527,3.5256753,3.7287042,3.9317331,4.1308575,4.3338866,4.5369153,4.3065557,4.0722914,3.8419318,3.6076677,3.3734035,3.5451972,3.7130866,3.8848803,4.056674,4.224563,4.4705405,4.716518,4.958591,5.2045684,5.4505453,4.8648853,4.279225,3.6935644,3.1118085,2.5261483,2.5456703,2.5651922,2.5847144,2.6042364,2.6237583,3.1039999,3.5842414,4.0644827,4.5447245,5.024966,5.2084727,5.388075,5.571582,5.755089,5.938596,5.481781,5.02887,4.572055,4.1191444,3.6623292,3.4788225,3.2992198,3.1157131,2.9322062,2.7486992,2.5066261,2.260649,2.0146716,1.7686942,1.5266213,1.8311646,2.1396124,2.4480603,2.7565079,3.0610514,3.3694992,3.677947,3.9863946,4.290938,4.5993857,4.5837684,4.564246,4.548629,4.5291066,4.513489,4.220659,3.9278288,3.6349986,3.3421683,3.049338,2.7916477,2.5300527,2.2684577,2.0107672,1.7491722,2.639376,3.5256753,4.4119744,5.298274,6.1884775,6.9459314,7.70729,8.468649,9.226103,9.987461,9.780528,9.573594,9.366661,9.155824,8.94889,7.519879,6.0908675,4.661856,3.2289407,1.7999294,2.1513257,2.5066261,2.8580225,3.2094188,3.5608149,4.415879,5.270943,6.126007,6.9810715,7.8361354,8.082112,8.32809,8.574067,8.81614,9.062118,9.190963,9.315904,9.444749,9.573594,9.698535,9.8312845,9.964035,10.096785,10.229534,10.362284,10.491129,10.6238785,10.752724,10.881569,11.014318,10.58093,10.147541,9.714153,9.280765,8.85128,8.65606,8.464745,8.273428,8.078208,7.8868923,7.6252975,7.363703,7.098203,6.8366084,6.575013,5.9659266,5.3607445,4.7516575,4.1464753,3.5373883,3.7599394,3.9824903,4.2050414,4.4275923,4.650143,4.83365,5.0210614,5.2045684,5.388075,5.575486,6.4852123,7.394938,8.304664,9.21439,10.124115,9.870329,9.616543,9.358852,9.105066,8.85128,8.148487,7.445695,6.7429028,6.04011,5.337318,4.9937305,4.6540475,4.31046,3.9668727,3.6232853,3.6232853,3.619381,3.619381,3.6154766,3.611572,3.39683,3.1781836,2.959537,2.7408905,2.5261483,2.4988174,2.475391,2.4480603,2.4246337,2.4012074,3.0102942,3.619381,4.2284675,4.841459,5.4505453,6.055728,6.66091,7.266093,7.871275,8.476458,8.207053,7.941554,7.6721506,7.406651,7.137247,6.949836,6.7624245,6.575013,6.387602,6.2001905,6.196286,6.196286,6.192382,6.1884775,6.1884775,6.0479193,5.9073606,5.7668023,5.6262436,5.4856853,5.466163,5.446641,5.4271193,5.407597,5.388075,6.0518236,6.7116675,7.375416,8.039165,8.699008,8.710721,8.718531,8.730244,8.738052,8.749765,8.0040245,7.2582836,6.5164475,5.7707067,5.024966,6.184573,7.3441806,8.503788,9.663396,10.826907,10.424754,10.0265045,9.6243515,9.226103,8.823949,8.531119,8.238289,7.9493628,7.656533,7.363703,8.335898,9.311999,10.2881,11.2642,12.236397,10.116306,7.9923115,5.8683167,3.7482262,1.6242313,1.8389735,2.0537157,2.2684577,2.4831998,2.7018464,3.2016098,3.7052777,4.2089458,4.7087092,5.212377,5.001539,4.7907014,4.5837684,4.3729305,4.1620927,3.6232853,3.0805733,2.541766,2.0029583,1.4641509,1.815547,2.1669433,2.5183394,2.87364,3.2250361,3.182088,3.1391394,3.096191,3.0532427,3.0141985,3.6740425,4.3338866,4.9937305,5.6535745,6.3134184,8.371038,10.4286585,12.486279,14.543899,16.601519,15.063184,13.524849,11.986515,10.44818,8.913751,9.171441,9.4291315,9.686822,9.940608,10.198298,9.889851,9.581403,9.269051,8.960603,8.648251,8.710721,8.769287,8.831758,8.890324,8.94889,8.23048,7.5081654,6.7897553,6.0713453,5.349031,5.434928,5.520825,5.606722,5.688714,5.774611,7.0708723,8.371038,9.6673,10.963562,12.263727,11.475039,10.686349,9.901564,9.112875,8.324185,8.402273,8.480362,8.55845,8.636538,8.710721,8.675582,8.636538,8.601398,8.562354,8.52331,8.433509,8.339804,8.246098,8.156297,8.062591,7.9220324,7.7814736,7.6409154,7.504261,7.363703,7.137247,6.910792,6.688241,6.461786,6.239235,5.0757227,3.9161155,2.7565079,1.5969005,0.43729305,0.4997635,0.5622339,0.62470436,0.6871748,0.74964523,0.8511597,0.94876975,1.0502841,1.1517987,1.2494087,1.4485333,1.6515622,1.8506867,2.0498111,2.2489357,2.4519646,2.6549935,2.8580225,3.0610514,3.2640803,3.135235,3.0063896,2.8814487,2.7526035,2.6237583,2.3543546,2.084951,1.815547,1.5461433,1.2767396,1.2337911,1.1947471,1.1557031,1.116659,1.0737107,0.9136301,0.74964523,0.58566034,0.42557985,0.26159495,0.44119745,0.62079996,0.80430686,0.98390937,1.1635119,1.3665408,1.5656652,1.7686942,1.9717231,2.174752,1.7413634,1.3040704,0.8706817,0.43338865,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.08589685,0.08589685,0.08589685,0.08589685,0.08589685,0.08589685,0.08199245,0.078088045,0.078088045,0.07418364,0.13665408,0.10932326,0.08199245,0.05466163,0.027330816,0.0,0.046852827,0.08980125,0.13665408,0.1796025,0.22645533,0.21864653,0.21474212,0.21083772,0.20693332,0.19912452,0.1639849,0.12494087,0.08589685,0.05075723,0.011713207,0.05075723,0.093705654,0.13274968,0.1717937,0.21083772,0.25378615,0.29673457,0.339683,0.38263142,0.42557985,0.62079996,0.8160201,1.0112402,1.2064602,1.4016805,1.3704453,1.33921,1.3118792,1.2806439,1.2494087,1.1713207,1.0893283,1.0112402,0.92924774,0.8511597,0.76916724,0.6910792,0.60908675,0.5309987,0.44900626,0.359205,0.26940376,0.1796025,0.08980125,0.0,0.0,0.0,0.0,0.0,0.0,0.10932326,0.21864653,0.3318742,0.44119745,0.5505207,0.64032197,0.7301232,0.8199245,0.9097257,0.999527,0.92534333,0.8511597,0.77307165,0.698888,0.62470436,0.81211567,0.999527,1.1869383,1.3743496,1.5617609,1.8116426,2.0615244,2.3114061,2.5612879,2.8111696,2.7135596,2.612045,2.514435,2.4129205,2.3114061,2.2918842,2.2684577,2.2450314,2.2216048,2.1981785,2.135708,2.0732377,2.0107672,1.9482968,1.8858263,2.4051118,2.9243972,3.4397783,3.959064,4.474445,4.704805,4.9351645,5.165524,5.395884,5.6262436,5.388075,5.153811,4.919547,4.6852827,4.4510183,4.7711797,5.0913405,5.4115014,5.7316628,6.0518236,5.727758,5.4036927,5.083532,4.759466,4.4393053,4.661856,4.884407,5.1069584,5.3256044,5.548156,5.8214636,6.094772,6.36808,6.6413884,6.910792,6.1455293,5.376362,4.6110992,3.8419318,3.076669,2.87364,2.6706111,2.4675822,2.2645533,2.0615244,2.2645533,2.4675822,2.6706111,2.87364,3.076669,3.2484627,3.4202564,3.59205,3.7638438,3.9356375,3.970777,4.0059166,4.041056,4.0761957,4.1113358,3.7130866,3.3187418,2.920493,2.522244,2.1239948,1.9522011,1.7804074,1.6086137,1.43682,1.261122,1.6710842,2.0810463,2.4910088,2.900971,3.310933,3.611572,3.9083066,4.2050414,4.5017757,4.7985106,4.6110992,4.4197836,4.2284675,4.041056,3.8497405,3.7599394,3.6701381,3.5803368,3.4905357,3.4007344,3.182088,2.9634414,2.7486992,2.5300527,2.3114061,3.349977,4.388548,5.423215,6.461786,7.5003567,8.441318,9.386183,10.327144,11.268105,12.212971,11.8537655,11.490656,11.131451,10.772245,10.413041,8.597494,6.7819467,4.9663997,3.1508527,1.33921,1.6086137,1.8780174,2.1474214,2.416825,2.6862288,3.2914112,3.892689,4.493967,5.099149,5.700427,6.2353306,6.7702336,7.3051367,7.8400397,8.374943,8.546737,8.714626,8.886419,9.054309,9.226103,9.2339115,9.245625,9.253433,9.265146,9.276859,9.4018,9.530646,9.655587,9.784432,9.913278,9.515028,9.116779,8.718531,8.324185,7.9259367,7.871275,7.8205175,7.7658563,7.715099,7.6643414,7.5394006,7.4105554,7.2856145,7.1606736,7.0357327,6.329036,5.618435,4.9078336,4.1972322,3.4866312,3.8692627,4.2479897,4.6267166,5.009348,5.388075,5.505207,5.6223392,5.7394714,5.8566036,5.9737353,6.8795567,7.785378,8.691199,9.593117,10.498938,10.010887,9.518932,9.030883,8.538928,8.050878,7.3910336,6.735094,6.0791545,5.4193106,4.7633705,4.661856,4.5564375,4.454923,4.3534083,4.251894,4.142571,4.0332475,3.9278288,3.8185053,3.7130866,3.3343596,2.9556324,2.5808098,2.2020829,1.8233559,1.901444,1.9756275,2.0498111,2.1239948,2.1981785,2.717464,3.2367494,3.7521305,4.271416,4.786797,5.602817,6.4188375,7.230953,8.046973,8.862993,8.699008,8.531119,8.367134,8.203149,8.039165,7.6643414,7.2856145,6.910792,6.5359693,6.1611466,6.2314262,6.297801,6.364176,6.434455,6.5008297,6.379793,6.2587566,6.141625,6.0205884,5.899552,5.7902284,5.6809053,5.571582,5.4583545,5.349031,6.1494336,6.949836,7.7502384,8.550641,9.351044,9.354948,9.358852,9.366661,9.370565,9.37447,8.538928,7.703386,6.871748,6.036206,5.2006636,6.2431393,7.2856145,8.32809,9.370565,10.413041,9.913278,9.413514,8.913751,8.413987,7.914223,7.6838636,7.4574084,7.230953,7.000593,6.774138,8.36323,9.948417,11.537509,13.1266,14.711788,11.943566,9.17925,6.4110284,3.6428072,0.8745861,1.2572175,1.639849,2.0224805,2.4051118,2.787743,3.5959544,4.4041657,5.2084727,6.016684,6.824895,6.5437784,6.266566,5.985449,5.704332,5.423215,4.5564375,3.6857557,2.815074,1.9443923,1.0737107,1.5969005,2.1161861,2.6354716,3.154757,3.6740425,3.5608149,3.4436827,3.330455,3.213323,3.1000953,3.5686235,4.0332475,4.5017757,4.970304,5.4388323,8.046973,10.6590185,13.2671585,15.879204,18.487345,16.539047,14.586847,12.63855,10.686349,8.738052,9.335425,9.932799,10.530173,11.127546,11.72492,11.205634,10.690253,10.170968,9.655587,9.136301,9.304191,9.47208,9.639969,9.807858,9.975748,8.738052,7.504261,6.27047,5.036679,3.7989833,4.369026,4.9351645,5.5013027,6.0713453,6.6374836,6.7429028,6.8483214,6.9537406,7.0591593,7.1606736,7.6252975,8.086017,8.550641,9.01136,9.475985,9.0465,8.6131115,8.183627,7.7541428,7.3246584,7.8361354,8.351517,8.862993,9.37447,9.885946,9.483793,9.081639,8.679486,8.277332,7.8751793,8.156297,8.433509,8.714626,8.995743,9.276859,8.374943,7.47693,6.575013,5.6730967,4.775084,3.8965936,3.0141985,2.135708,1.2533131,0.37482262,0.4997635,0.62470436,0.74964523,0.8745861,0.999527,1.1127546,1.2259823,1.33921,1.4485333,1.5617609,1.5617609,1.5617609,1.5617609,1.5617609,1.5617609,1.9717231,2.377781,2.7838387,3.193801,3.5998588,3.5686235,3.533484,3.5022488,3.4710135,3.435874,3.0883822,2.7408905,2.3933985,2.0459068,1.698415,1.5188124,1.3353056,1.1517987,0.96829176,0.78868926,0.698888,0.61299115,0.5231899,0.43729305,0.3513962,0.58956474,0.8316377,1.0698062,1.3118792,1.5500476,1.8194515,2.0888553,2.358259,2.631567,2.900971,2.3192148,1.7413634,1.1596074,0.58175594,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.078088045,0.08589685,0.08980125,0.093705654,0.10151446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.6481308,0.92534333,1.1986516,1.475864,1.7491722,1.7140326,1.6749885,1.6359446,1.6008049,1.5617609,1.4641509,1.3626363,1.261122,1.1635119,1.0619974,0.96438736,0.8628729,0.76135844,0.6637484,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.0,0.0,0.0,0.0,0.0,0.13665408,0.27330816,0.41386664,0.5505207,0.6871748,0.78868926,0.8862993,0.9878138,1.0893283,1.1869383,1.0893283,0.9878138,0.8862993,0.78868926,0.6871748,0.9019169,1.1127546,1.3235924,1.5383345,1.7491722,2.0107672,2.2762666,2.5378613,2.7994564,3.0610514,2.951728,2.8385005,2.7252727,2.612045,2.4988174,2.475391,2.4480603,2.4246337,2.4012074,2.3738766,2.3114061,2.2489357,2.1864653,2.1239948,2.0615244,2.6003318,3.1391394,3.6740425,4.21285,4.7516575,5.099149,5.4505453,5.801942,6.1494336,6.5008297,6.2743745,6.0518236,5.825368,5.5989127,5.376362,5.813655,6.250948,6.688241,7.125534,7.562827,7.1489606,6.7389984,6.3251314,5.911265,5.5013027,5.774611,6.0518236,6.3251314,6.5984397,6.8756523,7.1762915,7.47693,7.773665,8.074304,8.374943,7.426173,6.473499,5.5247293,4.575959,3.6232853,3.2016098,2.77603,2.35045,1.9248703,1.4992905,1.4251068,1.3509232,1.2767396,1.1986516,1.1244678,1.2884527,1.4485333,1.6125181,1.7765031,1.9365835,2.463678,2.9868677,3.513962,4.037152,4.564246,3.951255,3.338264,2.7252727,2.1122816,1.4992905,1.4016805,1.3001659,1.1986516,1.1010414,0.999527,1.5110037,2.0263848,2.5378613,3.049338,3.5608149,3.8497405,4.138666,4.423688,4.7126136,5.001539,4.6384296,4.2753205,3.912211,3.5491016,3.1859922,3.2992198,3.4124475,3.5256753,3.638903,3.7482262,3.5764325,3.4007344,3.2250361,3.049338,2.87364,4.0605783,5.251421,6.4383593,7.6252975,8.812236,9.936704,11.061172,12.185639,13.314012,14.438479,13.923099,13.411622,12.900145,12.388668,11.873287,9.675109,7.47693,5.2748475,3.076669,0.8745861,1.0619974,1.2494087,1.43682,1.6242313,1.8116426,2.1630387,2.514435,2.8619268,3.213323,3.5608149,4.388548,5.212377,6.036206,6.8639393,7.687768,7.898606,8.113348,8.324185,8.538928,8.749765,8.636538,8.52331,8.413987,8.300759,8.187531,8.312472,8.437413,8.562354,8.687295,8.812236,8.449126,8.086017,7.726812,7.363703,7.000593,7.08649,7.1762915,7.262188,7.348085,7.437886,7.4495993,7.461313,7.47693,7.4886436,7.5003567,6.688241,5.8761253,5.0640097,4.251894,3.435874,3.9746814,4.513489,5.0483923,5.5871997,6.126007,6.1767645,6.223617,6.2743745,6.3251314,6.375889,7.2739015,8.175818,9.073831,9.975748,10.87376,10.151445,9.425227,8.699008,7.9766936,7.250475,6.6374836,6.0244927,5.4115014,4.7985106,4.1894236,4.3260775,4.462732,4.5993857,4.73604,4.8765984,4.661856,4.4510183,4.2362766,4.025439,3.8106966,3.2757936,2.736986,2.1981785,1.6632754,1.1244678,1.3001659,1.475864,1.6515622,1.8233559,1.999054,2.4246337,2.8502135,3.2757936,3.7013733,4.123049,5.1499066,6.1767645,7.1997175,8.226576,9.249529,9.187058,9.124588,9.062118,8.999647,8.937177,8.374943,7.812709,7.250475,6.688241,6.126007,6.262661,6.3993154,6.5359693,6.676528,6.813182,6.7116675,6.6140575,6.5125427,6.4110284,6.3134184,6.114294,5.911265,5.7121406,5.5130157,5.3138914,6.250948,7.1880045,8.125061,9.062118,9.999174,9.999174,9.999174,9.999174,9.999174,9.999174,9.073831,8.148487,7.223144,6.3017054,5.376362,6.3017054,7.223144,8.148487,9.073831,9.999174,9.4018,8.800523,8.1992445,7.601871,7.000593,6.8366084,6.676528,6.5125427,6.348558,6.1884775,8.386656,10.588739,12.786918,14.989,17.18718,13.774731,10.362284,6.949836,3.5373883,0.12494087,0.6754616,1.2259823,1.7765031,2.3231194,2.87364,3.9863946,5.099149,6.211904,7.3246584,8.437413,8.086017,7.7385254,7.387129,7.0357327,6.688241,5.4856853,4.2870336,3.0883822,1.8858263,0.6871748,1.3743496,2.0615244,2.7486992,3.435874,4.123049,3.9356375,3.7482262,3.5608149,3.3734035,3.1859922,3.4632049,3.736513,4.0137253,4.2870336,4.564246,7.726812,10.885473,14.051944,17.210606,20.37317,18.011007,15.648844,13.286681,10.924518,8.562354,9.499411,10.436467,11.373524,12.31058,13.251541,12.525322,11.799104,11.076789,10.350571,9.6243515,9.901564,10.174872,10.44818,10.725393,10.998701,9.249529,7.5003567,5.7511845,3.998108,2.2489357,3.2992198,4.349504,5.3997884,6.4500723,7.5003567,6.4110284,5.3256044,4.2362766,3.1508527,2.0615244,3.775557,5.4856853,7.1997175,8.913751,10.6238785,9.686822,8.749765,7.812709,6.8756523,5.938596,7.000593,8.062591,9.124588,10.186585,11.248583,10.537982,9.823476,9.112875,8.398369,7.687768,8.386656,9.085544,9.788337,10.487225,11.186112,9.612638,8.039165,6.461786,4.8883114,3.310933,2.7135596,2.1122816,1.5110037,0.9136301,0.31235218,0.4997635,0.6871748,0.8745861,1.0619974,1.2494087,1.3743496,1.4992905,1.6242313,1.7491722,1.8741131,1.6749885,1.475864,1.2767396,1.0737107,0.8745861,1.4875772,2.1005683,2.7135596,3.3265507,3.9356375,3.998108,4.0605783,4.126953,4.1894236,4.251894,3.8263142,3.4007344,2.9751544,2.5495746,2.1239948,1.7999294,1.475864,1.1517987,0.8238289,0.4997635,0.48805028,0.47633708,0.46071947,0.44900626,0.43729305,0.737932,1.038571,1.33921,1.6359446,1.9365835,2.2762666,2.612045,2.951728,3.2875066,3.6232853,2.900971,2.174752,1.4485333,0.7262188,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.1756981,0.1639849,0.14836729,0.13665408,0.12494087,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.19131571,0.3318742,0.46852827,0.60908675,0.74964523,0.9917182,1.2337911,1.475864,1.7218413,1.9639144,1.901444,1.8389735,1.7765031,1.7140326,1.6515622,1.7804074,1.9092526,2.0420024,2.1708477,2.2996929,2.1669433,2.0302892,1.893635,1.7608855,1.6242313,1.3118792,0.999527,0.6871748,0.37482262,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.20302892,0.40605783,0.60908675,0.80821127,1.0112402,1.2415999,1.4719596,1.7023194,1.9326792,2.1630387,1.901444,1.6359446,1.3743496,1.1127546,0.8511597,1.0229534,1.1947471,1.3665408,1.5383345,1.7140326,2.0888553,2.4675822,2.8463092,3.2211318,3.5998588,3.4475873,3.2953155,3.1430438,2.9907722,2.8385005,2.8189783,2.7994564,2.77603,2.7565079,2.736986,2.6940374,2.6471848,2.6042364,2.5573835,2.514435,2.9243972,3.338264,3.7482262,4.1620927,4.575959,4.939069,5.298274,5.661383,6.0244927,6.387602,6.2470436,6.1064854,5.9659266,5.8292727,5.688714,6.055728,6.422742,6.7897553,7.1567693,7.523783,7.1450562,6.7663293,6.3836975,6.0049706,5.6262436,5.903456,6.184573,6.46569,6.746807,7.0240197,7.113821,7.2036223,7.2934237,7.3832245,7.473026,6.6140575,5.7511845,4.8883114,4.025439,3.1625657,2.8111696,2.455869,2.1044729,1.7530766,1.4016805,1.4446288,1.4914817,1.53443,1.5812829,1.6242313,1.7413634,1.8584955,1.9756275,2.096664,2.2137961,2.5300527,2.8463092,3.1664703,3.4827268,3.7989833,3.2836022,2.7643168,2.2489357,1.7296503,1.2142692,1.1713207,1.1322767,1.0932326,1.0541886,1.0112402,1.542239,2.0732377,2.6042364,3.1313305,3.6623292,3.853645,4.0488653,4.240181,4.4314966,4.6267166,4.376835,4.123049,3.873167,3.6232853,3.3734035,3.4905357,3.6037633,3.7208953,3.8341231,3.951255,3.9746814,3.998108,4.025439,4.0488653,4.0761957,5.040583,6.0049706,6.969358,7.9337454,8.898132,9.597021,10.295909,10.990892,11.68978,12.388668,11.900618,11.412568,10.924518,10.436467,9.948417,8.257811,6.5633,4.872694,3.1781836,1.4875772,1.6281357,1.7725986,1.9131571,2.05762,2.1981785,2.4714866,2.7408905,3.0102942,3.279698,3.5491016,4.380739,5.2162814,6.0479193,6.8795567,7.7111945,8.078208,8.449126,8.81614,9.183154,9.550168,9.468176,9.386183,9.304191,9.218294,9.136301,9.190963,9.245625,9.304191,9.358852,9.413514,8.991838,8.566258,8.144583,7.7229075,7.3012323,7.2582836,7.2192397,7.180196,7.141152,7.098203,7.008402,6.918601,6.8287997,6.7389984,6.649197,5.9268827,5.2006636,4.474445,3.7482262,3.0259118,3.4788225,3.9317331,4.380739,4.83365,5.2865605,5.3256044,5.3607445,5.3997884,5.4388323,5.473972,6.2314262,6.984976,7.7385254,8.495979,9.249529,8.636538,8.023546,7.4105554,6.801469,6.1884775,5.6652875,5.142098,4.618908,4.095718,3.5764325,3.736513,3.900498,4.0605783,4.224563,4.388548,4.290938,4.1972322,4.1035266,4.0059166,3.912211,3.3538816,2.7916477,2.233318,1.6710842,1.1127546,1.2376955,1.3626363,1.4875772,1.6125181,1.737459,2.096664,2.455869,2.8189783,3.1781836,3.5373883,4.435401,5.3334136,6.2314262,7.125534,8.023546,8.13287,8.238289,8.347612,8.453031,8.562354,8.13287,7.703386,7.2739015,6.844417,6.4110284,6.578918,6.746807,6.914696,7.082586,7.250475,7.266093,7.2856145,7.3012323,7.320754,7.336372,7.082586,6.8287997,6.571109,6.3173227,6.0635366,6.9927845,7.9220324,8.85128,9.784432,10.71368,10.670732,10.631687,10.592644,10.553599,10.510651,10.135828,9.761005,9.386183,9.01136,8.636538,9.331521,10.0265045,10.721489,11.416472,12.111456,11.303245,10.498938,9.690726,8.882515,8.074304,7.968885,7.859562,7.7541428,7.6448197,7.5394006,9.026978,10.518459,12.006037,13.497519,14.989,12.763491,10.541886,8.320281,6.098676,3.8770714,3.6154766,3.3538816,3.096191,2.8345962,2.5769055,3.4436827,4.3143644,5.185046,6.055728,6.9264097,7.0630636,7.1997175,7.336372,7.47693,7.6135845,6.3407493,5.067914,3.795079,2.522244,1.2494087,1.6867018,2.1200905,2.5534792,2.9907722,3.4241607,3.3616903,3.2992198,3.2367494,3.174279,3.1118085,3.3031244,3.4905357,3.6818514,3.873167,4.0605783,6.9615493,9.86252,12.763491,15.660558,18.56153,16.605423,14.653222,12.697116,10.741011,8.78881,9.475985,10.163159,10.850334,11.537509,12.224684,11.537509,10.850334,10.163159,9.475985,8.78881,9.245625,9.702439,10.159255,10.61607,11.076789,9.315904,7.558923,5.801942,4.044961,2.2879796,3.310933,4.3338866,5.35684,6.375889,7.3988423,6.4305506,5.4583545,4.4900627,3.521771,2.5495746,3.8067923,5.0640097,6.321227,7.578445,8.835662,8.160201,7.480835,6.805373,6.126007,5.4505453,6.2431393,7.039637,7.8361354,8.628729,9.425227,9.288573,9.148014,9.01136,8.874706,8.738052,8.902037,9.066022,9.2339115,9.397896,9.561881,8.207053,6.852226,5.4973984,4.142571,2.787743,2.6432803,2.4988174,2.3543546,2.2059872,2.0615244,1.8780174,1.6945106,1.5070993,1.3235924,1.1361811,1.2533131,1.3743496,1.4914817,1.6086137,1.7257458,1.6125181,1.4992905,1.3860629,1.2767396,1.1635119,1.8506867,2.5378613,3.2250361,3.912211,4.5993857,4.950782,5.298274,5.64967,6.001066,6.348558,5.8800297,5.4115014,4.939069,4.4705405,4.0020123,3.3226464,2.6432803,1.9678187,1.2884527,0.61299115,0.57394713,0.5309987,0.49195468,0.45291066,0.41386664,0.659844,0.9058213,1.1557031,1.4016805,1.6515622,1.9209659,2.1903696,2.4597735,2.7291772,2.998581,2.5456703,2.096664,1.6437533,1.1908426,0.737932,0.74574083,0.75354964,0.76135844,0.76916724,0.77697605,0.62470436,0.47633708,0.3240654,0.1756981,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.058566034,0.07027924,0.078088045,0.08980125,0.10151446,0.10151446,0.14836729,0.19912452,0.24988174,0.30063897,0.3513962,0.3240654,0.30063897,0.27330816,0.24988174,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.30454338,0.5114767,0.7145056,0.92143893,1.1244678,1.3353056,1.5461433,1.7530766,1.9639144,2.174752,2.0888553,1.999054,1.9131571,1.8233559,1.737459,2.096664,2.455869,2.8189783,3.1781836,3.5373883,3.3655949,3.1977055,3.0259118,2.8580225,2.6862288,2.174752,1.6632754,1.1517987,0.63641757,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.26940376,0.5349031,0.80430686,1.0698062,1.33921,1.698415,2.05762,2.416825,2.77603,3.1391394,2.7135596,2.2879796,1.8623998,1.43682,1.0112402,1.1439898,1.2767396,1.4094892,1.542239,1.6749885,2.1669433,2.6588979,3.1508527,3.6467118,4.138666,3.9434462,3.7521305,3.5608149,3.3655949,3.174279,3.1586614,3.1430438,3.1313305,3.1157131,3.1000953,3.0727646,3.0454338,3.018103,2.9907722,2.9634414,3.2484627,3.5373883,3.8263142,4.1113358,4.4002614,4.775084,5.1499066,5.5247293,5.899552,6.2743745,6.2197127,6.165051,6.1103897,6.055728,6.001066,6.297801,6.5945354,6.89127,7.191909,7.4886436,7.141152,6.79366,6.446168,6.098676,5.7511845,6.036206,6.321227,6.606249,6.89127,7.1762915,7.055255,6.9342184,6.813182,6.6960497,6.575013,5.801942,5.024966,4.251894,3.474918,2.7018464,2.4207294,2.1396124,1.8584955,1.5812829,1.3001659,1.4641509,1.6281357,1.796025,1.9600099,2.1239948,2.1981785,2.2684577,2.3426414,2.416825,2.4871042,2.5964274,2.7057507,2.8189783,2.9283018,3.0376248,2.6159496,2.194274,1.7686942,1.3470187,0.92534333,0.94486535,0.96438736,0.98390937,1.0034313,1.0268579,1.5734742,2.1200905,2.6667068,3.213323,3.7638438,3.8614538,3.959064,4.056674,4.154284,4.251894,4.1113358,3.9746814,3.8380275,3.7013733,3.5608149,3.6818514,3.7989833,3.9161155,4.0332475,4.1503797,4.376835,4.5993857,4.825841,5.0483923,5.2748475,6.016684,6.75852,7.504261,8.246098,8.987934,9.257338,9.526741,9.796145,10.069453,10.338858,9.874233,9.413514,8.94889,8.488171,8.023546,6.8405128,5.6535745,4.4705405,3.2836022,2.1005683,2.1981785,2.2957885,2.3933985,2.4910088,2.5886188,2.77603,2.9673457,3.1586614,3.3460727,3.5373883,4.376835,5.2162814,6.055728,6.899079,7.7385254,8.261715,8.781001,9.304191,9.82738,10.350571,10.295909,10.2451515,10.194394,10.139732,10.088976,10.073358,10.05774,10.042123,10.0265045,10.010887,9.530646,9.0465,8.566258,8.082112,7.601871,7.433982,7.266093,7.098203,6.930314,6.7624245,6.571109,6.375889,6.184573,5.9932575,5.801942,5.1616197,4.5252023,3.8887846,3.2484627,2.612045,2.979059,3.3460727,3.7130866,4.084005,4.4510183,4.474445,4.5017757,4.5252023,4.548629,4.575959,5.185046,5.794133,6.4032197,7.016211,7.6252975,7.125534,6.6257706,6.126007,5.6262436,5.12648,4.6930914,4.2597027,3.8263142,3.39683,2.9634414,3.1508527,3.338264,3.5256753,3.7130866,3.900498,3.9239242,3.9434462,3.9668727,3.9902992,4.0137253,3.4280653,2.8463092,2.2645533,1.6827974,1.1010414,1.175225,1.2494087,1.3235924,1.4016805,1.475864,1.7686942,2.0654287,2.358259,2.6549935,2.951728,3.7208953,4.4900627,5.2592297,6.028397,6.801469,7.0786815,7.355894,7.633106,7.910319,8.187531,7.890797,7.5940623,7.2934237,6.996689,6.699954,6.899079,7.094299,7.2934237,7.4886436,7.687768,7.824422,7.957172,8.093826,8.226576,8.36323,8.050878,7.7424297,7.433982,7.1216297,6.813182,7.734621,8.65606,9.581403,10.502842,11.424281,11.346193,11.2642,11.186112,11.10412,11.0260315,11.20173,11.373524,11.549222,11.72492,11.900618,12.365242,12.829865,13.29449,13.759113,14.223738,13.208592,12.193448,11.178304,10.163159,9.151918,9.097258,9.0465,8.991838,8.941081,8.886419,9.6673,10.44818,11.229061,12.006037,12.786918,11.756155,10.721489,9.690726,8.65606,7.6252975,6.5554914,5.4856853,4.415879,3.3460727,2.2762666,2.900971,3.5295796,4.1581883,4.786797,5.4115014,6.036206,6.66091,7.2856145,7.914223,8.538928,7.191909,5.8487945,4.5017757,3.1586614,1.8116426,1.9951496,2.1786566,2.358259,2.541766,2.7252727,2.787743,2.8502135,2.912684,2.9751544,3.0376248,3.1430438,3.2484627,3.3538816,3.4593005,3.5608149,6.2001905,8.835662,11.475039,14.114414,16.749886,15.203742,13.653695,12.107552,10.561408,9.01136,9.448653,9.885946,10.323239,10.764437,11.20173,10.549695,9.901564,9.249529,8.601398,7.9493628,8.589685,9.230007,9.870329,10.510651,11.150972,9.386183,7.621393,5.8566036,4.0918136,2.3231194,3.3187418,4.3143644,5.309987,6.3056097,7.3012323,6.446168,5.5950084,4.743849,3.8887846,3.0376248,3.8419318,4.6423345,5.446641,6.2470436,7.0513506,6.6335793,6.2158084,5.7980375,5.380266,4.9624953,5.4895897,6.016684,6.5437784,7.0708723,7.601871,8.039165,8.476458,8.913751,9.351044,9.788337,9.4174185,9.0465,8.675582,8.308568,7.9376497,6.801469,5.6691923,4.533011,3.39683,2.260649,2.5730011,2.8814487,3.193801,3.5022488,3.8106966,3.2562714,2.697942,2.1396124,1.5812829,1.0268579,1.1361811,1.2455044,1.3548276,1.4641509,1.5734742,1.5500476,1.5266213,1.4992905,1.475864,1.4485333,2.2137961,2.9751544,3.736513,4.5017757,5.263134,5.899552,6.5359693,7.1762915,7.812709,8.449126,7.9337454,7.4183645,6.902983,6.3915067,5.8761253,4.845363,3.814601,2.7838387,1.7530766,0.7262188,0.6559396,0.58956474,0.5231899,0.45681506,0.38653582,0.58175594,0.77697605,0.97219616,1.1674163,1.3626363,1.5656652,1.7686942,1.9717231,2.1708477,2.3738766,2.194274,2.0146716,1.8350691,1.6554666,1.475864,1.4914817,1.5031948,1.5188124,1.53443,1.5500476,1.2494087,0.94876975,0.6481308,0.3513962,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.039044023,0.046852827,0.05075723,0.058566034,0.06637484,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.44900626,0.5231899,0.48805028,0.44900626,0.41386664,0.37482262,0.3357786,0.26940376,0.20302892,0.13665408,0.06637484,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.42167544,0.6910792,0.96048295,1.2298868,1.4992905,1.678893,1.8545911,2.0341935,2.2098918,2.3855898,2.2762666,2.1630387,2.0498111,1.9365835,1.8233559,2.416825,3.0063896,3.5959544,4.185519,4.775084,4.5681505,4.365122,4.1581883,3.9551594,3.7482262,3.0376248,2.3231194,1.6125181,0.9019169,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.3318742,0.6637484,0.9956226,1.3314011,1.6632754,2.1513257,2.6432803,3.1313305,3.6232853,4.1113358,3.5256753,2.9361105,2.35045,1.7608855,1.175225,1.2689307,1.358732,1.4524376,1.5461433,1.6359446,2.2450314,2.854118,3.4593005,4.068387,4.6735697,4.4432096,4.2089458,3.978586,3.7443218,3.513962,3.5022488,3.49444,3.4827268,3.4710135,3.4632049,3.4514916,3.4436827,3.4319696,3.4241607,3.4124475,3.5764325,3.736513,3.900498,4.0605783,4.224563,4.6110992,5.001539,5.388075,5.774611,6.1611466,6.192382,6.223617,6.250948,6.282183,6.3134184,6.5398736,6.7663293,6.996689,7.223144,7.4495993,7.1333427,6.8209906,6.504734,6.1884775,5.8761253,6.165051,6.453977,6.746807,7.0357327,7.3246584,6.996689,6.6648145,6.336845,6.0049706,5.6730967,4.985922,4.298747,3.611572,2.9243972,2.2372224,2.0302892,1.8233559,1.6164225,1.4055848,1.1986516,1.4836729,1.7686942,2.0537157,2.338737,2.6237583,2.6510892,2.67842,2.7057507,2.7330816,2.7643168,2.6667068,2.5690966,2.4714866,2.3738766,2.2762666,1.9482968,1.620327,1.2923572,0.96438736,0.63641757,0.71841,0.79649806,0.8784905,0.95657855,1.038571,1.6008049,2.1669433,2.7330816,3.2992198,3.8614538,3.8653584,3.8692627,3.8692627,3.873167,3.873167,3.8497405,3.8263142,3.7989833,3.775557,3.7482262,3.8692627,3.9902992,4.1113358,4.2284675,4.349504,4.775084,5.2006636,5.6262436,6.0518236,6.473499,6.996689,7.5159745,8.03526,8.554545,9.073831,8.917655,8.761478,8.601398,8.445222,8.289046,7.8517528,7.4105554,6.9732623,6.5359693,6.098676,5.423215,4.743849,4.068387,3.3890212,2.7135596,2.7643168,2.8189783,2.8697357,2.9243972,2.9751544,3.084478,3.193801,3.3031244,3.416352,3.5256753,4.3729305,5.2201858,6.067441,6.914696,7.7619514,8.441318,9.116779,9.796145,10.471607,11.150972,11.127546,11.10412,11.080693,11.061172,11.037745,10.951848,10.865952,10.783959,10.698062,10.612165,10.069453,9.526741,8.98403,8.441318,7.898606,7.605776,7.309041,7.016211,6.719476,6.426646,6.1299114,5.833177,5.5403466,5.2436123,4.950782,4.4002614,3.8497405,3.2992198,2.7486992,2.1981785,2.4831998,2.7643168,3.049338,3.330455,3.611572,3.6232853,3.638903,3.6506162,3.6623292,3.6740425,4.138666,4.60329,5.0718184,5.5364423,6.001066,5.610626,5.22409,4.8375545,4.4510183,4.0605783,3.7208953,3.377308,3.0337205,2.6940374,2.35045,2.5612879,2.77603,2.9868677,3.2016098,3.4124475,3.5530062,3.6935644,3.8341231,3.970777,4.1113358,3.506153,2.900971,2.2957885,1.6906061,1.0893283,1.1127546,1.1361811,1.1635119,1.1869383,1.2142692,1.4407244,1.6710842,1.901444,2.1318035,2.3621633,3.0063896,3.6467118,4.290938,4.93126,5.575486,6.0205884,6.4695945,6.918601,7.363703,7.812709,7.648724,7.480835,7.3168497,7.152865,6.98888,7.2153354,7.4417906,7.6682463,7.898606,8.125061,8.378847,8.628729,8.882515,9.136301,9.386183,9.023073,8.65606,8.292951,7.9259367,7.562827,8.476458,9.393991,10.307622,11.221252,12.138786,12.01775,11.896713,11.775677,11.6585455,11.537509,12.263727,12.986042,13.712261,14.438479,15.160794,15.398962,15.633226,15.867491,16.101755,16.33602,15.113941,13.891863,12.6697855,11.447707,10.22563,10.22563,10.229534,10.2334385,10.2334385,10.237343,10.307622,10.377901,10.44818,10.518459,10.588739,10.744915,10.901091,11.061172,11.217348,11.373524,9.495506,7.6135845,5.735567,3.853645,1.9756275,2.358259,2.7447948,3.1313305,3.513962,3.900498,5.0132523,6.126007,7.238762,8.351517,9.464272,8.043069,6.6257706,5.2084727,3.7911747,2.3738766,2.3035975,2.233318,2.1669433,2.096664,2.0263848,2.2137961,2.4012074,2.5886188,2.77603,2.9634414,2.9829633,3.0024853,3.0220075,3.0415294,3.0610514,5.4388323,7.812709,10.186585,12.564366,14.938243,13.798158,12.658072,11.517986,10.377901,9.237816,9.425227,9.612638,9.80005,9.987461,10.174872,9.561881,8.94889,8.335898,7.726812,7.113821,7.9337454,8.757574,9.581403,10.401327,11.225157,9.452558,7.6799593,5.9073606,4.134762,2.3621633,3.330455,4.298747,5.263134,6.2314262,7.1997175,6.46569,5.7316628,4.9937305,4.2597027,3.5256753,3.873167,4.220659,4.5681505,4.9156423,5.263134,5.1030536,4.9468775,4.7907014,4.630621,4.474445,4.73604,4.9937305,5.2553253,5.5130157,5.774611,6.785851,7.800996,8.812236,9.823476,10.838621,9.932799,9.026978,8.121157,7.2192397,6.3134184,5.395884,4.482254,3.5686235,2.6510892,1.737459,2.5027218,3.2679846,4.0332475,4.7985106,5.563773,4.630621,3.7013733,2.7721257,1.8428779,0.9136301,1.0151446,1.116659,1.2181735,1.3235924,1.4251068,1.4875772,1.5500476,1.6125181,1.6749885,1.737459,2.5769055,3.4124475,4.251894,5.087436,5.9268827,6.8483214,7.773665,8.699008,9.6243515,10.549695,9.991365,9.4291315,8.870802,8.308568,7.7502384,6.36808,4.985922,3.6037633,2.2216048,0.8394465,0.7418364,0.6481308,0.5544251,0.45681506,0.3631094,0.5036679,0.6481308,0.78868926,0.93315214,1.0737107,1.2103647,1.3431144,1.4797685,1.6164225,1.7491722,1.8428779,1.9365835,2.0263848,2.1200905,2.2137961,2.233318,2.2567444,2.280171,2.3035975,2.3231194,1.8741131,1.4251068,0.97610056,0.5231899,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.031235218,0.03513962,0.039044023,0.046852827,0.05075723,0.19912452,0.30063897,0.39824903,0.4997635,0.60127795,0.698888,0.6481308,0.60127795,0.5505207,0.4997635,0.44900626,0.359205,0.26940376,0.1796025,0.08980125,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.5349031,0.8706817,1.2064602,1.5383345,1.8741131,2.018576,2.1669433,2.3114061,2.455869,2.6003318,2.463678,2.3231194,2.1864653,2.0498111,1.9131571,2.7330816,3.5530062,4.3729305,5.192855,6.012779,5.7707067,5.532538,5.2943697,5.0522966,4.814128,3.900498,2.9868677,2.0732377,1.1635119,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.39824903,0.79649806,1.1908426,1.5890918,1.9873407,2.6081407,3.2289407,3.8458362,4.466636,5.087436,4.337791,3.5881457,2.8385005,2.0888553,1.33921,1.3899672,1.4407244,1.4953861,1.5461433,1.6008049,2.3231194,3.0454338,3.767748,4.4900627,5.212377,4.939069,4.6657605,4.396357,4.123049,3.8497405,3.8458362,3.8419318,3.8341231,3.8302186,3.8263142,3.8341231,3.8419318,3.8458362,3.853645,3.8614538,3.900498,3.9356375,3.9746814,4.0137253,4.0488653,4.4510183,4.8492675,5.251421,5.64967,6.0518236,6.165051,6.278279,6.395411,6.5086384,6.6257706,6.7819467,6.9381227,7.098203,7.2543793,7.4105554,7.1294384,6.8483214,6.5633,6.282183,6.001066,6.2938967,6.590631,6.883461,7.180196,7.47693,6.9342184,6.395411,5.8566036,5.3138914,4.775084,4.173806,3.5764325,2.9751544,2.3738766,1.7765031,1.639849,1.5031948,1.3704453,1.2337911,1.1010414,1.5031948,1.9092526,2.3153105,2.7213683,3.1235218,3.1079042,3.0883822,3.0727646,3.0532427,3.0376248,2.7330816,2.4285383,2.1239948,1.815547,1.5110037,1.2806439,1.0463798,0.8160201,0.58175594,0.3513962,0.48805028,0.62860876,0.76916724,0.9097257,1.0502841,1.6320401,2.2137961,2.7994564,3.3812122,3.9629683,3.8692627,3.775557,3.6857557,3.59205,3.4983444,3.5881457,3.6740425,3.7638438,3.8497405,3.9356375,4.0605783,4.181615,4.3065557,4.4275923,4.548629,5.173333,5.801942,6.426646,7.0513506,7.676055,7.9727893,8.269524,8.566258,8.866898,9.163632,8.577971,7.9923115,7.406651,6.8209906,6.239235,5.825368,5.4115014,5.001539,4.5876727,4.173806,4.0059166,3.8341231,3.6662338,3.49444,3.3265507,3.3343596,3.338264,3.3460727,3.3538816,3.3616903,3.3929255,3.4241607,3.4514916,3.4827268,3.513962,4.369026,5.22409,6.0791545,6.9342184,7.7892823,8.62092,9.452558,10.284196,11.115833,11.951375,11.959184,11.963089,11.970898,11.978706,11.986515,11.834243,11.678067,11.521891,11.365715,11.213444,10.608261,10.006983,9.405705,8.804427,8.1992445,7.7775693,7.355894,6.9342184,6.5086384,6.086963,5.688714,5.2943697,4.8961205,4.4978714,4.0996222,3.638903,3.174279,2.7135596,2.2489357,1.7882162,1.9834363,2.182561,2.3816853,2.5769055,2.77603,2.77603,2.77603,2.77603,2.77603,2.77603,3.096191,3.416352,3.736513,4.056674,4.376835,4.0996222,3.8263142,3.5491016,3.2757936,2.998581,2.7486992,2.494913,2.241127,1.9912452,1.737459,1.9756275,2.2137961,2.4480603,2.6862288,2.9243972,3.182088,3.4397783,3.697469,3.9551594,4.21285,3.5842414,2.9556324,2.330928,1.7023194,1.0737107,1.0502841,1.0268579,0.999527,0.97610056,0.94876975,1.116659,1.2806439,1.4446288,1.6086137,1.7765031,2.2918842,2.803361,3.3187418,3.8341231,4.349504,4.9663997,5.5832953,6.2040954,6.8209906,7.437886,7.406651,7.3715115,7.3402762,7.309041,7.2739015,7.531592,7.7892823,8.046973,8.304664,8.562354,8.933272,9.304191,9.671205,10.042123,10.413041,9.991365,9.573594,9.151918,8.734148,8.312472,9.218294,10.128019,11.033841,11.943566,12.849388,12.689307,12.529227,12.369146,12.209065,12.0489855,13.325725,14.59856,15.875299,17.148134,18.424873,18.42878,18.436588,18.440493,18.444397,18.448301,17.019289,15.590279,14.161267,12.728352,11.29934,11.357906,11.416472,11.471134,11.5297,11.588266,10.947944,10.307622,9.6673,9.026978,8.386656,9.733675,11.080693,12.431617,13.778636,15.125654,12.435521,9.745388,7.055255,4.365122,1.6749885,1.8194515,1.9600099,2.1005683,2.2450314,2.3855898,3.9863946,5.5871997,7.1880045,8.78881,10.38571,8.898132,7.406651,5.919074,4.4275923,2.9361105,2.6159496,2.2918842,1.9717231,1.6476578,1.3235924,1.6359446,1.9482968,2.260649,2.5769055,2.8892577,2.822883,2.7565079,2.6940374,2.6276627,2.5612879,4.6735697,6.785851,8.898132,11.014318,13.1266,12.392572,11.6585455,10.928422,10.194394,9.464272,9.4018,9.339331,9.276859,9.21439,9.151918,8.574067,8.00012,7.426173,6.8483214,6.2743745,7.28171,8.285142,9.288573,10.295909,11.29934,9.518932,7.7385254,5.958118,4.181615,2.4012074,3.338264,4.279225,5.2201858,6.1611466,7.098203,6.481308,5.8644123,5.2475166,4.630621,4.0137253,3.9044023,3.7989833,3.68966,3.5842414,3.474918,3.5764325,3.6818514,3.7833657,3.8848803,3.9863946,3.978586,3.970777,3.9668727,3.959064,3.951255,5.5364423,7.125534,8.710721,10.299813,11.888905,10.44818,9.007456,7.5667315,6.126007,4.689187,3.9942036,3.2992198,2.6042364,1.9092526,1.2142692,2.4324427,3.6506162,4.872694,6.0908675,7.3129454,6.008875,4.7087092,3.4046388,2.1005683,0.80040246,0.8941081,0.9917182,1.0854238,1.1791295,1.2767396,1.4251068,1.5734742,1.7257458,1.8741131,2.0263848,2.9361105,3.8497405,4.7633705,5.6730967,6.5867267,7.800996,9.01136,10.22563,11.435994,12.650263,12.045081,11.4398985,10.834716,10.229534,9.6243515,7.890797,6.153338,4.4197836,2.6862288,0.94876975,0.8277333,0.7066968,0.58175594,0.46071947,0.3357786,0.42557985,0.5192855,0.60908675,0.698888,0.78868926,0.8550641,0.92143893,0.9917182,1.0580931,1.1244678,1.4914817,1.8545911,2.2216048,2.5847144,2.951728,2.979059,3.0102942,3.0415294,3.06886,3.1000953,2.4988174,1.901444,1.3001659,0.698888,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.011713207,0.015617609,0.015617609,0.019522011,0.023426414,0.023426414,0.24988174,0.37482262,0.4997635,0.62470436,0.74964523,0.8745861,0.81211567,0.74964523,0.6871748,0.62470436,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.6481308,1.0502841,1.4485333,1.8506867,2.2489357,2.3621633,2.475391,2.5886188,2.7018464,2.8111696,2.6510892,2.4871042,2.3231194,2.1630387,1.999054,3.049338,4.0996222,5.1499066,6.2001905,7.250475,6.9732623,6.699954,6.426646,6.1494336,5.8761253,4.7633705,3.6506162,2.5378613,1.4251068,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.46071947,0.92534333,1.3860629,1.8506867,2.3114061,3.0610514,3.8106966,4.564246,5.3138914,6.0635366,5.1499066,4.2362766,3.3265507,2.4129205,1.4992905,1.5110037,1.5266213,1.5383345,1.5500476,1.5617609,2.4012074,3.2367494,4.0761957,4.911738,5.7511845,5.4388323,5.12648,4.814128,4.5017757,4.1894236,4.1894236,4.1894236,4.1894236,4.1894236,4.1894236,4.21285,4.2362766,4.263607,4.2870336,4.3143644,4.224563,4.138666,4.0488653,3.9629683,3.873167,4.2870336,4.7009,5.1108627,5.5247293,5.938596,6.13772,6.336845,6.5359693,6.7389984,6.9381227,7.0240197,7.113821,7.1997175,7.2856145,7.375416,7.125534,6.8756523,6.6257706,6.375889,6.126007,6.426646,6.7233806,7.0240197,7.3246584,7.6252975,6.8756523,6.126007,5.376362,4.6267166,3.873167,3.3616903,2.8502135,2.338737,1.8233559,1.3118792,1.2494087,1.1869383,1.1244678,1.0619974,0.999527,1.5266213,2.0498111,2.5769055,3.1000953,3.6232853,3.5608149,3.4983444,3.435874,3.3734035,3.310933,2.7994564,2.2879796,1.7765031,1.261122,0.74964523,0.61299115,0.47633708,0.3357786,0.19912452,0.062470436,0.26159495,0.46071947,0.6637484,0.8628729,1.0619974,1.6632754,2.260649,2.8619268,3.4632049,4.0605783,3.873167,3.6857557,3.4983444,3.310933,3.1235218,3.3265507,3.5256753,3.7247996,3.9239242,4.123049,4.251894,4.376835,4.5017757,4.6267166,4.7516575,5.575486,6.3993154,7.223144,8.050878,8.874706,8.94889,9.023073,9.101162,9.175345,9.249529,8.238289,7.223144,6.211904,5.2006636,4.1894236,3.7989833,3.4124475,3.0259118,2.639376,2.2489357,2.5886188,2.9243972,3.2640803,3.5998588,3.9356375,3.900498,3.8614538,3.8263142,3.78727,3.7482262,3.7013733,3.6506162,3.5998588,3.5491016,3.4983444,4.3612175,5.22409,6.086963,6.949836,7.812709,8.800523,9.788337,10.77615,11.763964,12.751778,12.786918,12.825961,12.861101,12.900145,12.939189,12.712734,12.486279,12.263727,12.037272,11.810817,11.150972,10.487225,9.823476,9.163632,8.499884,7.9493628,7.3988423,6.8483214,6.3017054,5.7511845,5.251421,4.7516575,4.251894,3.7482262,3.2484627,2.87364,2.4988174,2.1239948,1.7491722,1.3743496,1.4875772,1.6008049,1.7140326,1.8233559,1.9365835,1.9248703,1.9131571,1.901444,1.8858263,1.8741131,2.0498111,2.2255092,2.4012074,2.5769055,2.7486992,2.5886188,2.4246337,2.260649,2.1005683,1.9365835,1.7765031,1.6125181,1.4485333,1.2884527,1.1244678,1.3860629,1.6515622,1.9131571,2.174752,2.436347,2.8111696,3.1859922,3.5608149,3.9356375,4.3143644,3.6623292,3.0141985,2.3621633,1.7140326,1.0619974,0.9878138,0.9136301,0.8394465,0.76135844,0.6871748,0.78868926,0.8862993,0.9878138,1.0893283,1.1869383,1.5734742,1.9639144,2.35045,2.736986,3.1235218,3.912211,4.7009,5.4856853,6.2743745,7.0630636,7.1606736,7.262188,7.363703,7.461313,7.562827,7.8517528,8.136774,8.4257,8.710721,8.999647,9.487698,9.975748,10.4637985,10.951848,11.435994,10.963562,10.487225,10.010887,9.538455,9.062118,9.964035,10.862047,11.763964,12.661977,13.563893,13.360865,13.16174,12.962616,12.763491,12.564366,14.387722,16.211079,18.038338,19.861694,21.688955,21.4625,21.236044,21.013493,20.787037,20.560583,18.924637,17.288692,15.648844,14.012899,12.373051,12.486279,12.599506,12.712734,12.825961,12.939189,11.588266,10.237343,8.886419,7.5394006,6.1884775,8.726339,11.2642,13.798158,16.33602,18.87388,15.375536,11.873287,8.374943,4.8765984,1.3743496,1.2767396,1.175225,1.0737107,0.97610056,0.8745861,2.9634414,5.0483923,7.137247,9.226103,11.311053,9.749292,8.187531,6.6257706,5.0640097,3.4983444,2.9243972,2.35045,1.7765031,1.1986516,0.62470436,1.0619974,1.4992905,1.9365835,2.3738766,2.8111696,2.6628022,2.514435,2.3621633,2.2137961,2.0615244,3.912211,5.7628975,7.6135845,9.464272,11.311053,10.986988,10.662923,10.338858,10.010887,9.686822,9.37447,9.062118,8.749765,8.437413,8.125061,7.5862536,7.0513506,6.5125427,5.9737353,5.4388323,6.6257706,7.812709,8.999647,10.186585,11.373524,9.589212,7.800996,6.012779,4.224563,2.436347,3.349977,4.263607,5.173333,6.086963,7.000593,6.5008297,6.001066,5.5013027,5.001539,4.5017757,3.9356375,3.3734035,2.8111696,2.2489357,1.6867018,2.0498111,2.4129205,2.77603,3.1391394,3.4983444,3.2250361,2.951728,2.6745155,2.4012074,2.1239948,4.2870336,6.4500723,8.6131115,10.77615,12.939189,10.963562,8.987934,7.012306,5.036679,3.0610514,2.5886188,2.1122816,1.6359446,1.1635119,0.6871748,2.3621633,4.037152,5.7121406,7.387129,9.062118,7.387129,5.7121406,4.037152,2.3621633,0.6871748,0.77307165,0.8628729,0.94876975,1.038571,1.1244678,1.3626363,1.6008049,1.8389735,2.0732377,2.3114061,3.2992198,4.2870336,5.2748475,6.262661,7.250475,8.749765,10.249056,11.748346,13.251541,14.750832,14.098797,13.450665,12.798631,12.150499,11.498465,9.413514,7.3246584,5.2358036,3.1508527,1.0619974,0.9136301,0.76135844,0.61299115,0.46071947,0.31235218,0.3513962,0.38653582,0.42557985,0.46071947,0.4997635,0.4997635,0.4997635,0.4997635,0.4997635,0.4997635,1.1361811,1.7765031,2.4129205,3.049338,3.6857557,3.7247996,3.7638438,3.7989833,3.8380275,3.873167,3.1235218,2.3738766,1.6242313,0.8745861,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.737932,0.8238289,0.9136301,0.999527,1.0893283,1.175225,1.1322767,1.0893283,1.0463798,1.0034313,0.96438736,0.9058213,0.8511597,0.79649806,0.7418364,0.6871748,0.6832704,0.679366,0.6715572,0.6676528,0.6637484,0.679366,0.6910792,0.7066968,0.7223144,0.737932,1.0112402,1.2806439,1.5539521,1.8272603,2.1005683,2.15523,2.2098918,2.2645533,2.3192148,2.3738766,2.2489357,2.1200905,1.9912452,1.8663043,1.737459,2.6667068,3.5959544,4.5291066,5.4583545,6.387602,6.2938967,6.2040954,6.1103897,6.016684,5.9268827,4.970304,4.0137253,3.0610514,2.1044729,1.1517987,1.0112402,0.8745861,0.737932,0.60127795,0.46071947,0.8667773,1.2728351,1.678893,2.0810463,2.4871042,3.1391394,3.7911747,4.4432096,5.099149,5.7511845,4.892216,4.0332475,3.1781836,2.3192148,1.4641509,1.5266213,1.5890918,1.6515622,1.7140326,1.7765031,2.5769055,3.3734035,4.173806,4.9742084,5.774611,5.466163,5.1616197,4.853172,4.5447245,4.2362766,4.3338866,4.4275923,4.521298,4.618908,4.7126136,4.728231,4.747753,4.7633705,4.7828927,4.7985106,4.732136,4.6657605,4.5993857,4.5291066,4.462732,4.950782,5.4388323,5.9268827,6.4110284,6.899079,7.238762,7.57454,7.914223,8.250002,8.58578,8.566258,8.542832,8.519405,8.495979,8.476458,8.218767,7.9649806,7.7111945,7.453504,7.1997175,7.3910336,7.578445,7.7697606,7.9610763,8.148487,7.2465706,6.3407493,5.434928,4.5291066,3.6232853,3.1586614,2.6940374,2.2294137,1.7647898,1.3001659,1.2689307,1.2415999,1.2103647,1.1791295,1.1517987,1.6320401,2.1161861,2.5964274,3.0805733,3.5608149,3.408543,3.2562714,3.1039999,2.951728,2.7994564,2.358259,1.9209659,1.4797685,1.038571,0.60127795,0.5036679,0.40996224,0.31625658,0.21864653,0.12494087,0.3631094,0.60127795,0.8394465,1.0737107,1.3118792,1.9170616,2.522244,3.1274261,3.7326086,4.337791,4.2011366,4.068387,3.9317331,3.7989833,3.6623292,3.7794614,3.892689,4.0059166,4.123049,4.2362766,4.2948427,4.3534083,4.40807,4.466636,4.5252023,5.1460023,5.7707067,6.3915067,7.016211,7.6370106,8.066495,8.495979,8.929368,9.358852,9.788337,8.804427,7.824422,6.8405128,5.8566036,4.8765984,4.447114,4.0215344,3.59205,3.1664703,2.736986,2.959537,3.182088,3.4046388,3.6271896,3.8497405,3.9668727,4.084005,4.2011366,4.318269,4.4393053,4.376835,4.318269,4.2557983,4.1972322,4.138666,4.884407,5.6340523,6.379793,7.1294384,7.8751793,8.663869,9.456462,10.2451515,11.033841,11.826434,11.763964,11.705398,11.6468315,11.584361,11.525795,11.564839,11.603884,11.6468315,11.685876,11.72492,10.955752,10.19049,9.421323,8.65606,7.8868923,7.6135845,7.336372,7.0630636,6.785851,6.5125427,6.196286,5.883934,5.5676775,5.251421,4.939069,4.650143,4.3612175,4.0761957,3.78727,3.4983444,3.4124475,3.3265507,3.2367494,3.1508527,3.0610514,3.0610514,3.0610514,3.0610514,3.0610514,3.0610514,3.084478,3.1079042,3.1313305,3.1508527,3.174279,3.0883822,3.0063896,2.920493,2.8345962,2.7486992,2.5573835,2.366068,2.1708477,1.979532,1.7882162,2.1044729,2.4207294,2.7408905,3.057147,3.3734035,3.619381,3.8614538,4.1035266,4.3455997,4.5876727,3.998108,3.4124475,2.8267872,2.2372224,1.6515622,1.5812829,1.5149081,1.4485333,1.3782539,1.3118792,1.3353056,1.358732,1.3782539,1.4016805,1.4251068,1.6906061,1.9600099,2.2294137,2.494913,2.7643168,3.506153,4.251894,4.997635,5.743376,6.4891167,6.7389984,6.9927845,7.2465706,7.4964523,7.7502384,8.093826,8.441318,8.784905,9.128492,9.475985,10.003078,10.530173,11.057267,11.584361,12.111456,11.966993,11.82253,11.678067,11.533605,11.389141,11.943566,12.501896,13.0602255,13.618555,14.176885,14.059752,13.946525,13.829392,13.716166,13.599033,14.770353,15.941674,17.10909,18.28041,19.451733,18.959778,18.471727,17.979773,17.491722,16.999767,15.992432,14.985096,13.97776,12.970425,11.963089,12.568271,13.173453,13.778636,14.383818,14.989,13.528754,12.072412,10.61607,9.155824,7.699481,9.487698,11.275913,13.06413,14.848442,16.636658,13.973856,11.311053,8.648251,5.989353,3.3265507,2.9322062,2.541766,2.1474214,1.756981,1.3626363,3.1118085,4.8570766,6.606249,8.351517,10.100689,9.589212,9.073831,8.562354,8.050878,7.5394006,6.348558,5.1616197,3.9746814,2.787743,1.6008049,1.7413634,1.8819219,2.018576,2.1591344,2.2996929,2.3270237,2.3543546,2.3816853,2.4090161,2.436347,3.8224099,5.2084727,6.590631,7.9766936,9.362757,9.358852,9.351044,9.347139,9.343235,9.339331,8.823949,8.308568,7.793187,7.277806,6.7624245,6.5281606,6.2938967,6.055728,5.8214636,5.5871997,6.493021,7.3988423,8.300759,9.20658,10.112402,8.538928,6.969358,5.395884,3.8224099,2.2489357,2.9556324,3.6662338,4.3729305,5.0796275,5.786324,5.520825,5.251421,4.985922,4.716518,4.4510183,4.193328,3.9356375,3.677947,3.4202564,3.1625657,3.3226464,3.4827268,3.6428072,3.802888,3.9629683,3.8185053,3.677947,3.533484,3.3929255,3.2484627,4.7985106,6.3446536,7.890797,9.440845,10.986988,9.4018,7.816613,6.2314262,4.646239,3.0610514,2.7213683,2.3816853,2.0420024,1.7023194,1.3626363,2.5651922,3.767748,4.970304,6.17286,7.375416,6.1181984,4.860981,3.6037633,2.3465457,1.0893283,1.0893283,1.0932326,1.0932326,1.097137,1.1010414,1.2728351,1.4446288,1.6164225,1.7882162,1.9639144,2.7643168,3.5686235,4.369026,5.173333,5.9737353,7.238762,8.499884,9.761005,11.0260315,12.287154,11.795199,11.303245,10.81129,10.315431,9.823476,8.32809,6.8287997,5.3334136,3.8341231,2.338737,2.1239948,1.9092526,1.6945106,1.475864,1.261122,1.0932326,0.92143893,0.75354964,0.58175594,0.41386664,0.40996224,0.40605783,0.40605783,0.40215343,0.39824903,0.9136301,1.4251068,1.9365835,2.4480603,2.9634414,3.0063896,3.0532427,3.096191,3.1430438,3.1859922,2.6237583,2.05762,1.4914817,0.92924774,0.3631094,0.29673457,0.22645533,0.16008049,0.093705654,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.2259823,1.2767396,1.3235924,1.3743496,1.4251068,1.475864,1.4524376,1.4290112,1.4055848,1.3860629,1.3626363,1.3665408,1.3665408,1.3704453,1.3743496,1.3743496,1.3665408,1.3548276,1.3431144,1.3353056,1.3235924,1.3040704,1.2845483,1.2650263,1.2455044,1.2259823,1.3704453,1.5149081,1.6593709,1.8038338,1.9482968,1.9482968,1.9443923,1.9443923,1.9404879,1.9365835,1.8467822,1.7530766,1.6593709,1.5656652,1.475864,2.2840753,3.096191,3.9044023,4.716518,5.5247293,5.6145306,5.704332,5.794133,5.883934,5.9737353,5.1772375,4.380739,3.5842414,2.7838387,1.9873407,1.7765031,1.5617609,1.3509232,1.1361811,0.92534333,1.2728351,1.620327,1.9678187,2.3153105,2.6628022,3.2172275,3.7716527,4.3260775,4.884407,5.4388323,4.6345253,3.8341231,3.0298162,2.2294137,1.4251068,1.5383345,1.6515622,1.7608855,1.8741131,1.9873407,2.7486992,3.513962,4.2753205,5.036679,5.801942,5.4973984,5.196759,4.892216,4.591577,4.2870336,4.478349,4.6657605,4.8570766,5.0483923,5.2358036,5.2475166,5.2592297,5.267039,5.278752,5.2865605,5.239708,5.192855,5.1460023,5.099149,5.0483923,5.610626,6.1767645,6.7389984,7.3012323,7.8634663,8.335898,8.812236,9.288573,9.761005,10.237343,10.104593,9.971844,9.839094,9.706344,9.573594,9.315904,9.054309,8.796618,8.535024,8.273428,8.355421,8.433509,8.515501,8.59359,8.675582,7.6135845,6.5554914,5.493494,4.435401,3.3734035,2.9556324,2.541766,2.1239948,1.7062237,1.2884527,1.2884527,1.2923572,1.2962615,1.2962615,1.3001659,1.7413634,2.1786566,2.619854,3.0610514,3.4983444,3.2562714,3.0141985,2.7721257,2.5300527,2.2879796,1.9209659,1.5539521,1.1869383,0.8160201,0.44900626,0.39824903,0.3435874,0.29283017,0.23816854,0.18741131,0.46071947,0.737932,1.0112402,1.2884527,1.5617609,2.1708477,2.7838387,3.3929255,4.0020123,4.6110992,4.5291066,4.447114,4.365122,4.283129,4.2011366,4.2284675,4.2597027,4.290938,4.318269,4.349504,4.3416953,4.3299823,4.318269,4.31046,4.298747,4.7204223,5.138193,5.559869,5.9815445,6.3993154,7.1841,7.968885,8.75367,9.538455,10.323239,9.370565,8.421796,7.4691215,6.5164475,5.563773,5.095245,4.6267166,4.1581883,3.6935644,3.2250361,3.3343596,3.4397783,3.5491016,3.6545205,3.7638438,4.0332475,4.3065557,4.579864,4.853172,5.12648,5.056201,4.985922,4.9156423,4.845363,4.775084,5.407597,6.04011,6.6726236,7.3051367,7.9376497,8.531119,9.120684,9.714153,10.307622,10.901091,10.741011,10.584834,10.4286585,10.268578,10.112402,10.416945,10.721489,11.0260315,11.330575,11.639023,10.764437,9.893755,9.019169,8.148487,7.2739015,7.2739015,7.2739015,7.2739015,7.2739015,7.2739015,7.1450562,7.016211,6.883461,6.754616,6.6257706,6.426646,6.223617,6.0244927,5.825368,5.6262436,5.337318,5.0483923,4.7633705,4.474445,4.185519,4.2011366,4.21285,4.224563,4.2362766,4.251894,4.1191444,3.9902992,3.8614538,3.7287042,3.5998588,3.59205,3.5842414,3.5764325,3.5686235,3.5608149,3.338264,3.1157131,2.893162,2.6706111,2.4480603,2.822883,3.193801,3.5686235,3.9395418,4.3143644,4.423688,4.533011,4.6423345,4.7516575,4.860981,4.337791,3.8106966,3.2875066,2.7643168,2.2372224,2.1786566,2.1161861,2.05762,1.999054,1.9365835,1.8819219,1.8272603,1.7725986,1.717937,1.6632754,1.8116426,1.9561055,2.1044729,2.25284,2.4012074,3.1039999,3.8067923,4.50568,5.2084727,5.911265,6.3173227,6.7233806,7.1294384,7.531592,7.9376497,8.339804,8.741957,9.14411,9.546264,9.948417,10.518459,11.084598,11.650736,12.220779,12.786918,12.974329,13.157836,13.341343,13.528754,13.712261,13.927003,14.141745,14.356487,14.571229,14.785972,14.75864,14.727406,14.69617,14.668839,14.637604,15.152986,15.668366,16.183748,16.69913,17.21451,16.457056,15.7035055,14.946052,14.192502,13.438952,13.0602255,12.681499,12.306676,11.927949,11.549222,12.6463585,13.743496,14.840633,15.941674,17.03881,15.473146,13.907481,12.341816,10.77615,9.21439,10.249056,11.287627,12.326198,13.360865,14.399435,12.576079,10.748819,8.925464,7.098203,5.2748475,4.591577,3.9044023,3.2211318,2.533957,1.8506867,3.2562714,4.6657605,6.0713453,7.480835,8.886419,9.425227,9.964035,10.498938,11.037745,11.576552,9.776623,7.9766936,6.1767645,4.376835,2.5769055,2.416825,2.260649,2.1005683,1.9443923,1.7882162,1.9912452,2.1981785,2.4012074,2.6081407,2.8111696,3.7326086,4.6540475,5.571582,6.493021,7.4144597,7.726812,8.043069,8.359325,8.671678,8.987934,8.269524,7.551114,6.8366084,6.1181984,5.3997884,5.466163,5.5364423,5.602817,5.6691923,5.735567,6.3602715,6.9810715,7.605776,8.226576,8.85128,7.492548,6.133816,4.7789884,3.4202564,2.0615244,2.5651922,3.06886,3.5686235,4.0722914,4.575959,4.5408196,4.50568,4.4705405,4.435401,4.4002614,4.447114,4.493967,4.5408196,4.591577,4.6384296,4.5954814,4.552533,4.5095844,4.466636,4.423688,4.415879,4.4041657,4.396357,4.3846436,4.376835,5.3060827,6.239235,7.172387,8.105539,9.0386915,7.843944,6.649197,5.4505453,4.2557983,3.0610514,2.8580225,2.6510892,2.4480603,2.241127,2.0380979,2.7682211,3.4983444,4.2284675,4.958591,5.688714,4.8492675,4.0059166,3.1664703,2.3270237,1.4875772,1.4055848,1.3235924,1.2415999,1.1557031,1.0737107,1.183034,1.2884527,1.397776,1.5031948,1.6125181,2.2294137,2.8463092,3.4632049,4.084005,4.7009,5.7238536,6.7507114,7.773665,8.800523,9.823476,9.491602,9.155824,8.8200445,8.484266,8.148487,7.2426662,6.336845,5.4271193,4.521298,3.611572,3.3343596,3.0532427,2.7721257,2.4910088,2.2137961,1.8350691,1.456342,1.0815194,0.7027924,0.3240654,0.32016098,0.31625658,0.30844778,0.30454338,0.30063897,0.6871748,1.0737107,1.4641509,1.8506867,2.2372224,2.2918842,2.3426414,2.3933985,2.4480603,2.4988174,2.1200905,1.7413634,1.358732,0.98000497,0.60127795,0.48805028,0.37872702,0.26940376,0.16008049,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.7140326,1.7257458,1.737459,1.7491722,1.7608855,1.7765031,1.7725986,1.7686942,1.7686942,1.7647898,1.7608855,1.8233559,1.8819219,1.9443923,2.0029583,2.0615244,2.0459068,2.0341935,2.018576,2.0029583,1.9873407,1.9326792,1.8780174,1.8233559,1.7686942,1.7140326,1.7296503,1.7491722,1.7647898,1.7843118,1.7999294,1.7413634,1.678893,1.620327,1.5617609,1.4992905,1.4407244,1.3860629,1.3274968,1.2689307,1.2142692,1.901444,2.592523,3.2836022,3.970777,4.661856,4.9351645,5.2084727,5.481781,5.7511845,6.0244927,5.3841705,4.743849,4.1035266,3.4632049,2.8267872,2.5378613,2.2489357,1.9639144,1.6749885,1.3860629,1.678893,1.9678187,2.2567444,2.5456703,2.8385005,3.2953155,3.7521305,4.2089458,4.6657605,5.12648,4.376835,3.631094,2.8814487,2.135708,1.3860629,1.5500476,1.7140326,1.8741131,2.0380979,2.1981785,2.9243972,3.6506162,4.376835,5.099149,5.825368,5.5286336,5.2318993,4.93126,4.6345253,4.337791,4.6228123,4.9078336,5.192855,5.477876,5.7628975,5.7668023,5.7668023,5.7707067,5.7707067,5.774611,5.74728,5.7199492,5.6926184,5.6652875,5.6379566,6.2743745,6.910792,7.551114,8.187531,8.823949,9.43694,10.049932,10.662923,11.275913,11.888905,11.6468315,11.400854,11.158782,10.916709,10.674636,10.409137,10.143637,9.878138,9.616543,9.351044,9.319808,9.288573,9.261242,9.230007,9.198771,7.984503,6.7702336,5.5559645,4.3416953,3.1235218,2.7565079,2.3855898,2.0146716,1.6437533,1.2767396,1.3118792,1.3431144,1.3782539,1.4133936,1.4485333,1.8467822,2.2450314,2.6432803,3.0415294,3.435874,3.1039999,2.7721257,2.4402514,2.1083772,1.7765031,1.4797685,1.1869383,0.8902037,0.59346914,0.30063897,0.28892577,0.28111696,0.26940376,0.26159495,0.24988174,0.5622339,0.8745861,1.1869383,1.4992905,1.8116426,2.4285383,3.0415294,3.6584249,4.271416,4.8883114,4.8570766,4.825841,4.7985106,4.7672753,4.73604,4.6813784,4.6267166,4.572055,4.5173936,4.462732,4.3846436,4.3065557,4.2284675,4.154284,4.0761957,4.290938,4.5095844,4.728231,4.9468775,5.1616197,6.3017054,7.4417906,8.581876,9.721962,10.862047,9.940608,9.019169,8.093826,7.172387,6.250948,5.743376,5.2358036,4.728231,4.220659,3.7130866,3.7052777,3.697469,3.68966,3.6818514,3.6740425,4.1035266,4.5291066,4.958591,5.3841705,5.813655,5.7316628,5.6535745,5.571582,5.493494,5.4115014,5.930787,6.446168,6.9654536,7.480835,8.00012,8.3944645,8.78881,9.183154,9.581403,9.975748,9.718058,9.464272,9.2104845,8.956698,8.699008,9.269051,9.839094,10.409137,10.979179,11.549222,10.573121,9.593117,8.617016,7.6409154,6.66091,6.9381227,7.211431,7.4886436,7.7619514,8.039165,8.093826,8.148487,8.203149,8.257811,8.312472,8.1992445,8.086017,7.9766936,7.8634663,7.7502384,7.262188,6.774138,6.2860875,5.801942,5.3138914,5.337318,5.3607445,5.388075,5.4115014,5.4388323,5.153811,4.872694,4.591577,4.3065557,4.025439,4.095718,4.165997,4.2362766,4.3065557,4.376835,4.123049,3.8692627,3.619381,3.3655949,3.1118085,3.541293,3.9668727,4.396357,4.8219366,5.251421,5.2279944,5.2045684,5.181142,5.1616197,5.138193,4.6735697,4.21285,3.7482262,3.2875066,2.8267872,2.7721257,2.7213683,2.6667068,2.6159496,2.5612879,2.4285383,2.2957885,2.1669433,2.0341935,1.901444,1.9287747,1.9561055,1.9834363,2.0107672,2.0380979,2.697942,3.357786,4.01763,4.677474,5.337318,5.8956475,6.453977,7.008402,7.5667315,8.125061,8.58578,9.0465,9.503315,9.964035,10.424754,11.033841,11.639023,12.24811,12.853292,13.462379,13.97776,14.493141,15.008522,15.523903,16.039284,15.9104395,15.781594,15.656653,15.527808,15.398962,15.453624,15.5082855,15.566852,15.621513,15.676175,15.535617,15.395058,15.254499,15.113941,14.973383,13.954333,12.935285,11.916236,10.893282,9.874233,10.128019,10.381805,10.631687,10.885473,11.139259,12.728352,14.317443,15.906535,17.495626,19.088623,17.413633,15.74255,14.0714655,12.396477,10.725393,11.014318,11.29934,11.588266,11.873287,12.162213,11.174399,10.186585,9.198771,8.210958,7.223144,6.2470436,5.270943,4.290938,3.3148375,2.338737,3.4046388,4.4705405,5.5403466,6.606249,7.676055,9.261242,10.850334,12.439425,14.024612,15.613705,13.200784,10.787864,8.374943,5.9620223,3.5491016,3.096191,2.639376,2.1864653,1.7296503,1.2767396,1.6593709,2.0380979,2.4207294,2.803361,3.1859922,3.6428072,4.095718,4.552533,5.009348,5.462259,6.098676,6.7311897,7.367607,8.0040245,8.636538,7.719003,6.7975645,5.8761253,4.958591,4.037152,4.40807,4.7789884,5.1460023,5.5169206,5.8878384,6.2275214,6.5672045,6.9068875,7.2465706,7.5862536,6.446168,5.3021784,4.1581883,3.018103,1.8741131,2.1708477,2.4714866,2.7682211,3.0649557,3.3616903,3.5608149,3.7560349,3.9551594,4.154284,4.349504,4.7009,5.056201,5.407597,5.758993,6.114294,5.8683167,5.6223392,5.376362,5.134289,4.8883114,5.009348,5.134289,5.2553253,5.376362,5.5013027,5.8175592,6.133816,6.453977,6.7702336,7.08649,6.282183,5.477876,4.6735697,3.8692627,3.0610514,2.9907722,2.9243972,2.854118,2.7838387,2.7135596,2.97125,3.2289407,3.4866312,3.7443218,3.998108,3.5764325,3.154757,2.7330816,2.3114061,1.8858263,1.7218413,1.5539521,1.3860629,1.2181735,1.0502841,1.0932326,1.1361811,1.1791295,1.2181735,1.261122,1.6945106,2.1278992,2.5612879,2.9907722,3.4241607,4.21285,5.001539,5.786324,6.575013,7.363703,7.1841,7.008402,6.8287997,6.6531014,6.473499,6.1572423,5.840986,5.520825,5.2045684,4.8883114,4.5408196,4.1972322,3.853645,3.506153,3.1625657,2.5769055,1.9912452,1.4055848,0.8238289,0.23816854,0.23035973,0.22255093,0.21474212,0.20693332,0.19912452,0.46071947,0.7262188,0.9878138,1.2494087,1.5110037,1.5734742,1.6320401,1.6906061,1.7530766,1.8116426,1.6164225,1.4212024,1.2259823,1.0307622,0.8394465,0.6832704,0.5309987,0.37872702,0.22645533,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.1981785,2.174752,2.1513257,2.1239948,2.1005683,2.0732377,2.0927596,2.1083772,2.1278992,2.1435168,2.1630387,2.280171,2.397303,2.514435,2.631567,2.7486992,2.7291772,2.7096553,2.690133,2.6706111,2.6510892,2.5612879,2.4714866,2.3816853,2.2918842,2.1981785,2.0888553,1.979532,1.8702087,1.7608855,1.6515622,1.53443,1.4133936,1.2962615,1.1791295,1.0619974,1.038571,1.0190489,0.9956226,0.97219616,0.94876975,1.5188124,2.0888553,2.6588979,3.2289407,3.7989833,4.2557983,4.7087092,5.165524,5.618435,6.0752497,5.591104,5.1108627,4.6267166,4.1464753,3.6623292,3.2992198,2.9361105,2.5769055,2.2137961,1.8506867,2.0810463,2.3153105,2.5456703,2.7799344,3.0141985,3.3734035,3.7326086,4.0918136,4.4510183,4.814128,4.1191444,3.4280653,2.7330816,2.0420024,1.3509232,1.5617609,1.7765031,1.9873407,2.1981785,2.4129205,3.1000953,3.78727,4.474445,5.1616197,5.8487945,5.5559645,5.263134,4.9742084,4.6813784,4.388548,4.7672753,5.1460023,5.5286336,5.9073606,6.2860875,6.282183,6.278279,6.2743745,6.266566,6.262661,6.2548523,6.2470436,6.239235,6.2314262,6.223617,6.9381227,7.648724,8.36323,9.073831,9.788337,10.537982,11.287627,12.037272,12.786918,13.536563,13.185166,12.83377,12.47847,12.127073,11.775677,11.506273,11.23687,10.963562,10.694158,10.424754,10.284196,10.143637,10.003078,9.866425,9.725866,8.355421,6.984976,5.6145306,4.2440853,2.87364,2.5534792,2.2294137,1.9092526,1.5851873,1.261122,1.3314011,1.397776,1.4641509,1.53443,1.6008049,1.9561055,2.3114061,2.6667068,3.018103,3.3734035,2.951728,2.5300527,2.1083772,1.6867018,1.261122,1.038571,0.8160201,0.59346914,0.3709182,0.14836729,0.1835069,0.21474212,0.24597734,0.28111696,0.31235218,0.6637484,1.0112402,1.3626363,1.7140326,2.0615244,2.6823244,3.3031244,3.9239242,4.5408196,5.1616197,5.185046,5.2084727,5.2318993,5.251421,5.2748475,5.134289,4.9937305,4.853172,4.716518,4.575959,4.4314966,4.283129,4.138666,3.9942036,3.8497405,3.8653584,3.8809757,3.8965936,3.9083066,3.9239242,5.4193106,6.914696,8.410083,9.905469,11.400854,10.506746,9.616543,8.722435,7.8283267,6.9381227,6.3915067,5.840986,5.2943697,4.747753,4.2011366,4.0761957,3.9551594,3.8341231,3.7091823,3.5881457,4.169902,4.7516575,5.3334136,5.919074,6.5008297,6.4110284,6.321227,6.2314262,6.141625,6.0518236,6.453977,6.8561306,7.2582836,7.660437,8.062591,8.261715,8.456935,8.65606,8.85128,9.050405,8.699008,8.343708,7.9923115,7.6409154,7.2856145,8.121157,8.956698,9.792241,10.627783,11.4633255,10.381805,9.296382,8.214863,7.1333427,6.0518236,6.5984397,7.1489606,7.699481,8.250002,8.800523,9.0386915,9.280765,9.518932,9.761005,9.999174,9.975748,9.948417,9.924991,9.901564,9.874233,9.187058,8.499884,7.812709,7.125534,6.4383593,6.473499,6.5125427,6.551587,6.5867267,6.6257706,6.1884775,5.755089,5.3217,4.884407,4.4510183,4.5993857,4.743849,4.892216,5.040583,5.1889505,4.903929,4.6228123,4.3416953,4.056674,3.775557,4.2557983,4.7399445,5.22409,5.704332,6.1884775,6.0323014,5.8761253,5.7238536,5.5676775,5.4115014,5.0132523,4.6110992,4.21285,3.8106966,3.4124475,3.3655949,3.3226464,3.2757936,3.232845,3.1859922,2.979059,2.7682211,2.5573835,2.3465457,2.135708,2.0459068,1.9522011,1.8584955,1.7686942,1.6749885,2.2918842,2.9087796,3.5256753,4.1464753,4.7633705,5.473972,6.180669,6.89127,7.601871,8.312472,8.831758,9.347139,9.866425,10.381805,10.901091,11.549222,12.193448,12.841579,13.48971,14.13784,14.981192,15.828446,16.671797,17.519053,18.362404,17.893875,17.421442,16.952915,16.484386,16.011953,16.152512,16.29307,16.43363,16.574188,16.710842,15.918248,15.12175,14.329156,13.532659,12.73616,11.4516115,10.167064,8.882515,7.5979667,6.3134184,7.195813,8.078208,8.960603,9.8429985,10.725393,12.806439,14.89139,16.972437,19.053482,21.138433,19.358027,17.57762,15.797212,14.016804,12.236397,11.775677,11.311053,10.850334,10.38571,9.924991,9.776623,9.6243515,9.475985,9.323712,9.175345,7.9064145,6.6335793,5.364649,4.095718,2.8267872,3.5530062,4.279225,5.009348,5.735567,6.461786,9.101162,11.736633,14.376009,17.01148,19.650856,16.624945,13.599033,10.573121,7.551114,4.5252023,3.7716527,3.018103,2.2684577,1.5149081,0.76135844,1.3235924,1.8819219,2.4441557,3.0024853,3.5608149,3.5530062,3.541293,3.533484,3.521771,3.513962,4.466636,5.423215,6.375889,7.3324676,8.289046,7.164578,6.044015,4.919547,3.7989833,2.6745155,3.3460727,4.0215344,4.6930914,5.364649,6.036206,6.094772,6.153338,6.211904,6.266566,6.3251314,5.395884,4.4705405,3.541293,2.6159496,1.6867018,1.7804074,1.8741131,1.9639144,2.05762,2.1513257,2.5808098,3.0102942,3.4397783,3.8692627,4.298747,4.958591,5.6145306,6.2743745,6.930314,7.5862536,7.141152,6.6921453,6.2431393,5.7980375,5.349031,5.606722,5.860508,6.114294,6.36808,6.6257706,6.329036,6.028397,5.7316628,5.434928,5.138193,4.7243266,4.3065557,3.892689,3.4788225,3.0610514,3.1274261,3.193801,3.2562714,3.3226464,3.3890212,3.174279,2.9556324,2.7408905,2.5261483,2.3114061,2.3075018,2.3035975,2.2957885,2.2918842,2.2879796,2.0341935,1.7843118,1.5305257,1.2767396,1.0268579,1.0034313,0.98000497,0.95657855,0.93315214,0.9136301,1.1596074,1.4055848,1.6554666,1.901444,2.1513257,2.7018464,3.2484627,3.7989833,4.349504,4.900025,4.8805027,4.860981,4.841459,4.8180323,4.7985106,5.0718184,5.3451266,5.618435,5.891743,6.1611466,5.7511845,5.3412223,4.93126,4.521298,4.1113358,3.3187418,2.5261483,1.7335546,0.94096094,0.14836729,0.14055848,0.12884527,0.12103647,0.10932326,0.10151446,0.23816854,0.37482262,0.5114767,0.6481308,0.78868926,0.8550641,0.92143893,0.9917182,1.0580931,1.1244678,1.116659,1.1049459,1.0932326,1.0854238,1.0737107,0.8784905,0.6832704,0.48805028,0.29673457,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.6862288,2.6237583,2.5612879,2.4988174,2.436347,2.3738766,2.4129205,2.4480603,2.4871042,2.5261483,2.5612879,2.736986,2.912684,3.0883822,3.2640803,3.435874,3.4124475,3.3890212,3.3616903,3.338264,3.310933,3.1859922,3.0610514,2.9361105,2.8111696,2.6862288,2.4480603,2.2137961,1.9756275,1.737459,1.4992905,1.3235924,1.1517987,0.97610056,0.80040246,0.62470436,0.63641757,0.6481308,0.6637484,0.6754616,0.6871748,1.1361811,1.5890918,2.0380979,2.4871042,2.9361105,3.5764325,4.21285,4.8492675,5.4856853,6.126007,5.801942,5.473972,5.1499066,4.825841,4.5017757,4.0605783,3.6232853,3.1859922,2.7486992,2.3114061,2.4871042,2.6628022,2.8385005,3.0141985,3.1859922,3.4514916,3.7130866,3.9746814,4.2362766,4.5017757,3.8614538,3.2250361,2.5886188,1.9482968,1.3118792,1.5734742,1.8389735,2.1005683,2.3621633,2.6237583,3.2757936,3.9239242,4.575959,5.22409,5.8761253,5.5871997,5.298274,5.0132523,4.7243266,4.4393053,4.911738,5.388075,5.8644123,6.336845,6.813182,6.801469,6.785851,6.774138,6.7624245,6.7507114,6.7624245,6.774138,6.785851,6.801469,6.813182,7.601871,8.386656,9.175345,9.964035,10.748819,11.639023,12.525322,13.411622,14.301826,15.188125,14.723501,14.262781,13.798158,13.337439,12.8767185,12.599506,12.326198,12.0489855,11.775677,11.498465,11.248583,10.998701,10.748819,10.498938,10.249056,8.726339,7.1997175,5.6730967,4.1503797,2.6237583,2.35045,2.0732377,1.7999294,1.5266213,1.2494087,1.3509232,1.4485333,1.5500476,1.6515622,1.7491722,2.0615244,2.3738766,2.6862288,2.998581,3.310933,2.7994564,2.2879796,1.7765031,1.261122,0.74964523,0.60127795,0.44900626,0.30063897,0.14836729,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.76135844,1.1517987,1.5383345,1.9248703,2.3114061,2.9361105,3.5608149,4.1894236,4.814128,5.4388323,5.5130157,5.5871997,5.661383,5.735567,5.813655,5.5871997,5.3607445,5.138193,4.911738,4.689187,4.474445,4.263607,4.0488653,3.8380275,3.6232853,3.435874,3.2484627,3.0610514,2.87364,2.6862288,4.5369153,6.387602,8.238289,10.088976,11.935758,11.076789,10.213917,9.351044,8.488171,7.6252975,7.0357327,6.4500723,5.8644123,5.2748475,4.689187,4.4510183,4.21285,3.9746814,3.736513,3.4983444,4.2362766,4.9742084,5.7121406,6.4500723,7.1880045,7.08649,6.98888,6.8873653,6.785851,6.688241,6.9732623,7.262188,7.551114,7.8361354,8.125061,8.125061,8.125061,8.125061,8.125061,8.125061,7.676055,7.223144,6.774138,6.3251314,5.8761253,6.9732623,8.074304,9.175345,10.276386,11.373524,10.186585,8.999647,7.812709,6.6257706,5.4388323,6.262661,7.08649,7.914223,8.738052,9.561881,9.987461,10.413041,10.838621,11.2642,11.685876,11.748346,11.810817,11.873287,11.935758,11.998228,11.111929,10.22563,9.339331,8.449126,7.562827,7.6135845,7.6643414,7.7111945,7.7619514,7.812709,7.223144,6.6374836,6.0518236,5.462259,4.8765984,5.099149,5.3256044,5.548156,5.774611,6.001066,5.688714,5.376362,5.0640097,4.7516575,4.4393053,4.9742084,5.5130157,6.0518236,6.5867267,7.125534,6.8366084,6.551587,6.262661,5.9737353,5.688714,5.349031,5.0132523,4.6735697,4.337791,3.998108,3.9629683,3.9239242,3.8887846,3.8497405,3.8106966,3.5256753,3.2367494,2.951728,2.6628022,2.3738766,2.1630387,1.9482968,1.737459,1.5266213,1.3118792,1.8858263,2.463678,3.0376248,3.611572,4.1894236,5.0483923,5.911265,6.774138,7.6370106,8.499884,9.073831,9.651682,10.22563,10.799577,11.373524,12.0606985,12.751778,13.438952,14.126127,14.813302,15.988527,17.163752,18.338978,19.514202,20.689428,19.873407,19.061293,18.249176,17.437061,16.624945,16.8514,17.073952,17.300406,17.526861,17.749413,16.300879,14.848442,13.399908,11.951375,10.498938,8.94889,7.3988423,5.8487945,4.298747,2.7486992,4.263607,5.774611,7.2856145,8.800523,10.311526,12.888432,15.461433,18.038338,20.61134,23.188246,21.298513,19.412687,17.526861,15.637131,13.751305,12.537036,11.326671,10.112402,8.898132,7.687768,8.374943,9.062118,9.749292,10.436467,11.123642,9.561881,8.00012,6.4383593,4.8765984,3.310933,3.7013733,4.087909,4.474445,4.860981,5.251421,8.937177,12.626837,16.312593,19.998348,23.68801,20.049105,16.414106,12.775204,9.136301,5.5013027,4.4510183,3.4007344,2.35045,1.3001659,0.24988174,0.9878138,1.7257458,2.463678,3.2016098,3.9356375,3.4632049,2.9868677,2.514435,2.0380979,1.5617609,2.8385005,4.1113358,5.388075,6.66091,7.9376497,6.6140575,5.2865605,3.9629683,2.639376,1.3118792,2.2879796,3.2640803,4.2362766,5.212377,6.1884775,5.9620223,5.735567,5.5130157,5.2865605,5.0640097,4.349504,3.638903,2.9243972,2.2137961,1.4992905,1.3860629,1.2767396,1.1635119,1.0502841,0.93705654,1.6008049,2.260649,2.9243972,3.5881457,4.251894,5.212377,6.1767645,7.137247,8.101635,9.062118,8.413987,7.7619514,7.113821,6.461786,5.813655,6.2001905,6.5867267,6.9732623,7.363703,7.7502384,6.8366084,5.9268827,5.0132523,4.0996222,3.1859922,3.1625657,3.1391394,3.1118085,3.0883822,3.0610514,3.2640803,3.4632049,3.6623292,3.8614538,4.0605783,3.3734035,2.6862288,1.999054,1.3118792,0.62470436,1.038571,1.4485333,1.8623998,2.2762666,2.6862288,2.35045,2.0107672,1.6749885,1.33921,0.999527,0.9136301,0.8238289,0.737932,0.6481308,0.5622339,0.62470436,0.6871748,0.74964523,0.81211567,0.8745861,1.1869383,1.4992905,1.8116426,2.1239948,2.436347,2.5769055,2.7135596,2.8502135,2.9868677,3.1235218,3.9863946,4.8492675,5.7121406,6.575013,7.437886,6.9615493,6.4891167,6.012779,5.5364423,5.0640097,4.0605783,3.0610514,2.0615244,1.0619974,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.13665408,0.21083772,0.28892577,0.3631094,0.43729305,0.61299115,0.78868926,0.96438736,1.1361811,1.3118792,1.0737107,0.8394465,0.60127795,0.3631094,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.5612879,2.4910088,2.416825,2.3465457,2.2723622,2.1981785,2.338737,2.4792955,2.619854,2.7604125,2.900971,3.0727646,3.2445583,3.416352,3.5881457,3.7638438,3.7989833,3.8341231,3.8692627,3.9044023,3.9356375,3.8106966,3.6818514,3.5569105,3.4280653,3.2992198,3.0063896,2.7096553,2.416825,2.1200905,1.8233559,1.7062237,1.5890918,1.4719596,1.3548276,1.2376955,1.2337911,1.2337911,1.2298868,1.2259823,1.2259823,1.5539521,1.8858263,2.2137961,2.5456703,2.87364,3.5530062,4.2284675,4.9078336,5.5832953,6.262661,6.012779,5.7628975,5.5130157,5.263134,5.0132523,4.6110992,4.21285,3.8106966,3.4124475,3.0141985,3.1235218,3.2367494,3.349977,3.4632049,3.5764325,3.8106966,4.044961,4.279225,4.513489,4.7516575,4.263607,3.7794614,3.2953155,2.8111696,2.3231194,2.5730011,2.8189783,3.06886,3.3148375,3.5608149,4.084005,4.607195,5.1303844,5.6535745,6.1767645,5.891743,5.606722,5.3217,5.036679,4.7516575,5.1460023,5.5442514,5.9425,6.3407493,6.7389984,6.8209906,6.902983,6.984976,7.066968,7.1489606,7.08649,7.0240197,6.9615493,6.899079,6.8366084,7.473026,8.105539,8.741957,9.378374,10.010887,10.71368,11.412568,12.111456,12.814248,13.513136,13.192975,12.8767185,12.560462,12.244205,11.924045,11.818625,11.709302,11.603884,11.49456,11.389141,10.838621,10.2881,9.737579,9.187058,8.636538,7.355894,6.0791545,4.7985106,3.5178664,2.2372224,2.0537157,1.8741131,1.6906061,1.5070993,1.3235924,1.4407244,1.5617609,1.678893,1.796025,1.9131571,2.096664,2.2762666,2.4597735,2.6432803,2.8267872,2.3855898,1.9443923,1.5031948,1.0659018,0.62470436,0.5466163,0.46852827,0.39434463,0.31625658,0.23816854,0.39824903,0.5622339,0.7262188,0.8862993,1.0502841,1.3665408,1.678893,1.9951496,2.3114061,2.6237583,3.154757,3.6857557,4.2167544,4.743849,5.2748475,5.395884,5.520825,5.6418614,5.7668023,5.8878384,5.6730967,5.462259,5.251421,5.036679,4.825841,4.50568,4.1894236,3.873167,3.5569105,3.2367494,3.1391394,3.0415294,2.9439192,2.8463092,2.7486992,4.3455997,5.938596,7.535496,9.128492,10.725393,10.147541,9.56969,8.991838,8.413987,7.8361354,7.238762,6.6413884,6.044015,5.446641,4.8492675,4.661856,4.474445,4.2870336,4.0996222,3.912211,4.6696653,5.4271193,6.184573,6.942027,7.699481,7.6409154,7.578445,7.519879,7.461313,7.3988423,7.6135845,7.8283267,8.046973,8.261715,8.476458,8.570163,8.663869,8.761478,8.855185,8.94889,8.445222,7.941554,7.433982,6.930314,6.426646,7.3402762,8.253906,9.171441,10.085071,10.998701,10.147541,9.296382,8.441318,7.590158,6.7389984,7.676055,8.617016,9.557977,10.498938,11.435994,11.900618,12.361338,12.825961,13.286681,13.751305,13.833297,13.919194,14.005091,14.090988,14.176885,13.333533,12.494087,11.654641,10.815194,9.975748,9.745388,9.515028,9.284669,9.054309,8.823949,8.207053,7.590158,6.9732623,6.356367,5.7394714,5.903456,6.067441,6.2314262,6.3993154,6.5633,6.473499,6.3836975,6.2938967,6.2040954,6.114294,6.5633,7.012306,7.461313,7.914223,8.36323,8.296855,8.226576,8.160201,8.093826,8.023546,7.621393,7.2153354,6.8092775,6.4032197,6.001066,5.805846,5.6145306,5.423215,5.2318993,5.036679,4.8102236,4.5837684,4.3534083,4.126953,3.900498,3.5842414,3.2640803,2.9478238,2.631567,2.3114061,2.6862288,3.057147,3.4319696,3.802888,4.173806,4.8765984,5.575486,6.2743745,6.9732623,7.676055,8.378847,9.085544,9.788337,10.495033,11.20173,12.009941,12.818152,13.630268,14.438479,15.250595,16.378967,17.503435,18.631807,19.76018,20.888552,20.459068,20.025679,19.596195,19.16671,18.737226,18.374117,18.011007,17.651802,17.288692,16.925583,15.793307,14.664935,13.536563,12.404286,11.275913,10.0226,8.769287,7.5159745,6.266566,5.0132523,6.321227,7.629202,8.933272,10.241247,11.549222,14.461906,17.37459,20.287273,23.199959,26.112642,23.961317,21.813896,19.662569,17.511244,15.363823,14.118319,12.8767185,11.6351185,10.393518,9.151918,9.530646,9.913278,10.295909,10.67854,11.061172,9.80005,8.538928,7.2739015,6.012779,4.7516575,5.044488,5.3334136,5.6262436,5.919074,6.211904,9.237816,12.263727,15.285735,18.311647,21.337559,18.057861,14.782067,11.506273,8.226576,4.950782,4.0332475,3.1157131,2.1981785,1.2806439,0.3631094,0.96438736,1.5617609,2.1630387,2.7643168,3.3616903,3.4632049,3.5686235,3.6701381,3.7716527,3.8770714,5.4036927,6.930314,8.456935,9.983557,11.514082,9.729771,7.9493628,6.165051,4.380739,2.6003318,3.1235218,3.6467118,4.165997,4.689187,5.212377,5.0210614,4.825841,4.6345253,4.4432096,4.251894,3.8458362,3.4397783,3.0337205,2.631567,2.2255092,2.1669433,2.1083772,2.0537157,1.9951496,1.9365835,2.416825,2.8970666,3.377308,3.8575494,4.337791,5.1108627,5.8878384,6.66091,7.437886,8.210958,7.6643414,7.1177254,6.571109,6.0205884,5.473972,5.989353,6.5008297,7.012306,7.523783,8.039165,7.000593,5.9620223,4.9234514,3.8887846,2.8502135,2.795552,2.7447948,2.6940374,2.639376,2.5886188,2.736986,2.8892577,3.0376248,3.1859922,3.338264,2.7916477,2.2489357,1.7023194,1.1557031,0.61299115,0.94096094,1.2728351,1.6008049,1.9326792,2.260649,1.9717231,1.678893,1.3860629,1.0932326,0.80040246,0.7301232,0.659844,0.58956474,0.5192855,0.44900626,0.58175594,0.7145056,0.8472553,0.98000497,1.1127546,1.397776,1.6827974,1.9678187,2.25284,2.5378613,2.7057507,2.87364,3.0415294,3.2094188,3.3734035,4.0059166,4.6384296,5.270943,5.903456,6.5359693,6.0908675,5.6418614,5.196759,4.747753,4.298747,3.4671092,2.6354716,1.8038338,0.96829176,0.13665408,0.10932326,0.08199245,0.05466163,0.027330816,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.1717937,0.24597734,0.31625658,0.39044023,0.46071947,0.6832704,0.9058213,1.1283722,1.3509232,1.5734742,1.3118792,1.0502841,0.78868926,0.5231899,0.26159495,0.21083772,0.15617609,0.10541886,0.05075723,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.436347,2.3543546,2.2723622,2.1903696,2.1083772,2.0263848,2.2684577,2.5105307,2.7526035,2.9946766,3.2367494,3.408543,3.5764325,3.7482262,3.9161155,4.087909,4.181615,4.279225,4.3729305,4.466636,4.564246,4.4314966,4.3026514,4.173806,4.041056,3.912211,3.5608149,3.2094188,2.854118,2.5027218,2.1513257,2.0888553,2.0302892,1.9717231,1.9092526,1.8506867,1.8311646,1.815547,1.796025,1.7804074,1.7608855,1.9717231,2.182561,2.3933985,2.6042364,2.8111696,3.5295796,4.2479897,4.9663997,5.6809053,6.3993154,6.223617,6.0518236,5.8761253,5.700427,5.5247293,5.1616197,4.7985106,4.4393053,4.0761957,3.7130866,3.7638438,3.8106966,3.8614538,3.912211,3.9629683,4.169902,4.376835,4.5837684,4.7907014,5.001539,4.6657605,4.3338866,4.0020123,3.6701381,3.338264,3.5686235,3.802888,4.0332475,4.267512,4.5017757,4.8961205,5.290465,5.6848097,6.0791545,6.473499,6.192382,5.911265,5.6262436,5.3451266,5.0640097,5.3841705,5.704332,6.0205884,6.3407493,6.66091,6.8405128,7.016211,7.195813,7.3715115,7.551114,7.4105554,7.2739015,7.137247,7.000593,6.8639393,7.3441806,7.8283267,8.308568,8.792714,9.276859,9.788337,10.299813,10.81129,11.326671,11.838148,11.666354,11.490656,11.318862,11.147068,10.975275,11.033841,11.096312,11.154878,11.213444,11.275913,10.424754,9.573594,8.726339,7.8751793,7.0240197,5.989353,4.9546866,3.9200199,2.8853533,1.8506867,1.7608855,1.6710842,1.5812829,1.4914817,1.4016805,1.53443,1.6710842,1.8038338,1.9404879,2.0732377,2.1278992,2.1786566,2.233318,2.2840753,2.338737,1.9717231,1.6008049,1.2337911,0.8667773,0.4997635,0.4958591,0.48805028,0.48414588,0.48024148,0.47633708,0.7262188,0.97610056,1.2259823,1.475864,1.7257458,1.9678187,2.2098918,2.4519646,2.6940374,2.9361105,3.3734035,3.8067923,4.2440853,4.677474,5.1108627,5.282656,5.4505453,5.6223392,5.794133,5.9620223,5.7628975,5.563773,5.3607445,5.1616197,4.9624953,4.5408196,4.1191444,3.6935644,3.2718892,2.8502135,2.8424048,2.8345962,2.8267872,2.8189783,2.8111696,4.154284,5.493494,6.832704,8.171914,9.511124,9.218294,8.929368,8.636538,8.343708,8.050878,7.4417906,6.8366084,6.2275214,5.618435,5.0132523,4.8765984,4.73604,4.5993857,4.462732,4.3260775,5.1030536,5.8800297,6.657006,7.433982,8.210958,8.191436,8.171914,8.152391,8.13287,8.113348,8.253906,8.398369,8.538928,8.683391,8.823949,9.0152645,9.20658,9.393991,9.585307,9.776623,9.21439,8.65606,8.093826,7.535496,6.9732623,7.703386,8.433509,9.163632,9.893755,10.6238785,10.108498,9.589212,9.073831,8.554545,8.039165,9.093353,10.147541,11.20173,12.2559185,13.314012,13.813775,14.313539,14.813302,15.313066,15.812829,15.918248,16.02757,16.13299,16.242313,16.351637,15.559043,14.766449,13.973856,13.181262,12.388668,11.877192,11.365715,10.858143,10.346666,9.839094,9.190963,8.542832,7.8947015,7.2465706,6.5984397,6.703859,6.8092775,6.914696,7.0201154,7.125534,7.2582836,7.3910336,7.523783,7.656533,7.7892823,8.148487,8.511597,8.874706,9.237816,9.600925,9.753197,9.905469,10.05774,10.2100115,10.362284,9.889851,9.4174185,8.944985,8.472553,8.00012,7.6526284,7.3051367,6.957645,6.610153,6.262661,6.094772,5.9268827,5.758993,5.591104,5.423215,5.001539,4.579864,4.1581883,3.736513,3.310933,3.4827268,3.6506162,3.8224099,3.9942036,4.1620927,4.7009,5.2358036,5.774611,6.3134184,6.8483214,7.6838636,8.519405,9.354948,10.19049,11.0260315,11.959184,12.888432,13.821584,14.754736,15.687888,16.769407,17.847023,18.928543,20.006157,21.087677,21.040823,20.99397,20.943214,20.89636,20.849508,19.900738,18.948065,17.999294,17.050524,16.101755,15.289639,14.481428,13.6693125,12.861101,12.0489855,11.096312,10.139732,9.183154,8.23048,7.2739015,8.378847,9.479889,10.58093,11.685876,12.786918,16.039284,19.287746,22.53621,25.788576,29.037039,26.624119,24.211199,21.798277,19.389261,16.976341,15.7035055,14.430671,13.157836,11.885,10.612165,10.690253,10.768341,10.84643,10.920613,10.998701,10.0382185,9.073831,8.113348,7.1489606,6.1884775,6.3836975,6.5828223,6.7780423,6.9771667,7.1762915,9.538455,11.900618,14.262781,16.624945,18.987108,16.07052,13.153932,10.2334385,7.3168497,4.4002614,3.6154766,2.8306916,2.0459068,1.261122,0.47633708,0.93705654,1.4016805,1.8623998,2.3231194,2.787743,3.4671092,4.1464753,4.825841,5.5091114,6.1884775,7.968885,9.749292,11.525795,13.306203,15.086611,12.845484,10.608261,8.367134,6.126007,3.8887846,3.959064,4.029343,4.095718,4.165997,4.2362766,4.0761957,3.9161155,3.7560349,3.5959544,3.435874,3.338264,3.240654,3.1430438,3.049338,2.951728,2.9478238,2.9439192,2.9439192,2.9400148,2.9361105,3.2367494,3.533484,3.8302186,4.126953,4.423688,5.0132523,5.5989127,6.1884775,6.774138,7.363703,6.918601,6.473499,6.028397,5.5832953,5.138193,5.774611,6.4110284,7.0513506,7.687768,8.324185,7.1606736,6.001066,4.8375545,3.6740425,2.514435,2.4324427,2.3543546,2.2723622,2.194274,2.1122816,2.2137961,2.3114061,2.4129205,2.514435,2.612045,2.2098918,1.8077383,1.4055848,1.0034313,0.60127795,0.8472553,1.0932326,1.3431144,1.5890918,1.8389735,1.5890918,1.3431144,1.0932326,0.8472553,0.60127795,0.5466163,0.4958591,0.44119745,0.39044023,0.3357786,0.5388075,0.7418364,0.94486535,1.1478943,1.3509232,1.6086137,1.8663043,2.1239948,2.3816853,2.639376,2.8345962,3.0337205,3.2289407,3.4280653,3.6232853,4.029343,4.4314966,4.83365,5.2358036,5.6379566,5.2162814,4.7985106,4.376835,3.959064,3.5373883,2.87364,2.2059872,1.542239,0.8784905,0.21083772,0.1717937,0.12884527,0.08589685,0.042948425,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.20693332,0.27721256,0.3474918,0.41777104,0.48805028,0.75745404,1.0268579,1.2962615,1.5656652,1.8389735,1.5500476,1.261122,0.97610056,0.6871748,0.39824903,0.32016098,0.23816854,0.16008049,0.078088045,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.3114061,2.2216048,2.1278992,2.0341935,1.9443923,1.8506867,2.194274,2.541766,2.8853533,3.2289407,3.5764325,3.7443218,3.9083066,4.0761957,4.2440853,4.4119744,4.5681505,4.7243266,4.8765984,5.0327744,5.1889505,5.056201,4.9234514,4.7907014,4.657952,4.5252023,4.11524,3.7052777,3.2953155,2.8853533,2.475391,2.4714866,2.4714866,2.4675822,2.463678,2.463678,2.4285383,2.397303,2.366068,2.330928,2.2996929,2.3894942,2.4792955,2.5690966,2.6588979,2.7486992,3.506153,4.263607,5.0210614,5.7785153,6.5359693,6.4383593,6.336845,6.239235,6.13772,6.036206,5.7121406,5.388075,5.0640097,4.73604,4.4119744,4.4002614,4.388548,4.376835,4.3612175,4.349504,4.5291066,4.7087092,4.8883114,5.0718184,5.251421,5.0718184,4.8883114,4.7087092,4.5291066,4.349504,4.5681505,4.786797,5.001539,5.2201858,5.4388323,5.704332,5.9737353,6.239235,6.5086384,6.774138,6.4969254,6.2158084,5.9346914,5.6535745,5.376362,5.618435,5.860508,6.1025805,6.3446536,6.5867267,6.860035,7.1333427,7.406651,7.676055,7.9493628,7.7385254,7.523783,7.3129454,7.098203,6.8873653,7.2192397,7.5472097,7.8790836,8.207053,8.538928,8.862993,9.187058,9.511124,9.839094,10.163159,10.135828,10.108498,10.081166,10.053836,10.0265045,10.25296,10.479416,10.705871,10.936231,11.162686,10.010887,8.862993,7.7111945,6.5633,5.4115014,4.6228123,3.8341231,3.0415294,2.25284,1.4641509,1.4641509,1.4680552,1.4680552,1.4719596,1.475864,1.6281357,1.7804074,1.9326792,2.084951,2.2372224,2.1591344,2.0810463,2.0068626,1.9287747,1.8506867,1.5539521,1.261122,0.96438736,0.6715572,0.37482262,0.44119745,0.5114767,0.57785153,0.6442264,0.7106012,1.0502841,1.3860629,1.7257458,2.0615244,2.4012074,2.5690966,2.7408905,2.9087796,3.0805733,3.2484627,3.5881457,3.9317331,4.271416,4.6110992,4.950782,5.169429,5.3841705,5.602817,5.8214636,6.036206,5.8487945,5.661383,5.473972,5.2865605,5.099149,4.572055,4.044961,3.5178664,2.9907722,2.463678,2.5456703,2.6276627,2.7096553,2.7916477,2.87364,3.959064,5.044488,6.1299114,7.2153354,8.300759,8.292951,8.285142,8.277332,8.269524,8.261715,7.6448197,7.027924,6.4110284,5.794133,5.173333,5.087436,5.001539,4.911738,4.825841,4.73604,5.5364423,6.3329406,7.1294384,7.9259367,8.726339,8.745861,8.765383,8.784905,8.804427,8.823949,8.894228,8.964508,9.034787,9.105066,9.175345,9.460366,9.745388,10.03041,10.315431,10.600452,9.983557,9.370565,8.75367,8.140678,7.523783,8.070399,8.6131115,9.159728,9.706344,10.249056,10.069453,9.885946,9.702439,9.518932,9.339331,10.506746,11.678067,12.849388,14.016804,15.188125,15.726933,16.261835,16.800642,17.33945,17.874353,18.003199,18.135948,18.264793,18.393639,18.526388,17.780647,17.034906,16.289165,15.543426,14.801589,14.008995,13.220306,12.431617,11.639023,10.850334,10.170968,9.495506,8.81614,8.140678,7.461313,7.5081654,7.551114,7.5979667,7.6409154,7.687768,8.043069,8.398369,8.75367,9.108971,9.464272,9.737579,10.010887,10.2881,10.561408,10.838621,11.209538,11.584361,11.955279,12.326198,12.70102,12.158309,11.619501,11.080693,10.541886,9.999174,9.499411,8.995743,8.492075,7.988407,7.4886436,7.37932,7.2739015,7.164578,7.0591593,6.949836,6.422742,5.8956475,5.368553,4.841459,4.3143644,4.279225,4.2479897,4.2167544,4.181615,4.1503797,4.5252023,4.900025,5.2748475,5.64967,6.0244927,6.98888,7.9532676,8.921559,9.885946,10.850334,11.904523,12.958711,14.016804,15.070992,16.125181,17.155943,18.19061,19.221373,20.256039,21.2868,21.62258,21.958359,22.294136,22.62601,22.96179,21.423454,19.889025,18.35069,16.812357,15.274021,14.785972,14.294017,13.805966,13.314012,12.825961,12.166118,11.510178,10.8542385,10.194394,9.538455,10.436467,11.334479,12.228588,13.1266,14.024612,17.612759,21.200905,24.78905,28.373291,31.961437,29.28692,26.612406,23.937891,21.263374,18.58886,17.284788,15.980719,14.6805525,13.376482,12.076316,11.845957,11.619501,11.393045,11.166591,10.936231,10.276386,9.612638,8.94889,8.289046,7.6252975,7.726812,7.8283267,7.9337454,8.03526,8.136774,9.839094,11.537509,13.235924,14.938243,16.636658,14.079274,11.521891,8.964508,6.407124,3.8497405,3.1977055,2.5456703,1.893635,1.2415999,0.58566034,0.9136301,1.2376955,1.5617609,1.8858263,2.2137961,3.4710135,4.728231,5.985449,7.2426662,8.499884,10.534078,12.564366,14.59856,16.628849,18.663042,15.965101,13.2671585,10.569217,7.871275,5.173333,4.7907014,4.4119744,4.029343,3.6467118,3.2640803,3.135235,3.0063896,2.8814487,2.7526035,2.6237583,2.8345962,3.0454338,3.2562714,3.4632049,3.6740425,3.7287042,3.7794614,3.8341231,3.8848803,3.9356375,4.0527697,4.165997,4.283129,4.396357,4.513489,4.911738,5.3138914,5.7121406,6.114294,6.5125427,6.168956,5.8292727,5.4856853,5.142098,4.7985106,5.563773,6.3251314,7.08649,7.8517528,8.6131115,7.3246584,6.036206,4.7516575,3.4632049,2.174752,2.069333,1.9600099,1.8506867,1.7452679,1.6359446,1.6867018,1.737459,1.7882162,1.8389735,1.8858263,1.6281357,1.3665408,1.1088502,0.8472553,0.58566034,0.75354964,0.91753453,1.0815194,1.2494087,1.4133936,1.2103647,1.0073358,0.80430686,0.60127795,0.39824903,0.3631094,0.3318742,0.29673457,0.26159495,0.22645533,0.4958591,0.76916724,1.0424755,1.3157835,1.5890918,1.8194515,2.0459068,2.2762666,2.5066261,2.736986,2.9634414,3.193801,3.4202564,3.6467118,3.873167,4.0488653,4.220659,4.3924527,4.564246,4.73604,4.3455997,3.951255,3.5608149,3.1664703,2.77603,2.2762666,1.7804074,1.2806439,0.78478485,0.28892577,0.23035973,0.1717937,0.113227665,0.058566034,0.0,0.03513962,0.07027924,0.10541886,0.14055848,0.1756981,0.24207294,0.30844778,0.37872702,0.44510186,0.5114767,0.8316377,1.1478943,1.4641509,1.7843118,2.1005683,1.7882162,1.475864,1.1635119,0.8511597,0.5388075,0.42948425,0.3240654,0.21474212,0.10932326,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.1864653,2.084951,1.9834363,1.8819219,1.7765031,1.6749885,2.1239948,2.5690966,3.018103,3.4632049,3.912211,4.0761957,4.2440853,4.40807,4.572055,4.73604,4.950782,5.169429,5.3841705,5.5989127,5.813655,5.677001,5.5442514,5.407597,5.270943,5.138193,4.6696653,4.2011366,3.736513,3.2679846,2.7994564,2.854118,2.9087796,2.9634414,3.018103,3.076669,3.0259118,2.979059,2.9322062,2.8853533,2.8385005,2.8072653,2.77603,2.7486992,2.717464,2.6862288,3.4866312,4.283129,5.0796275,5.8761253,6.676528,6.649197,6.6257706,6.5984397,6.575013,6.551587,6.262661,5.9737353,5.688714,5.3997884,5.1108627,5.036679,4.9624953,4.8883114,4.814128,4.73604,4.8883114,5.040583,5.196759,5.349031,5.5013027,5.473972,5.446641,5.4193106,5.388075,5.3607445,5.563773,5.7668023,5.969831,6.17286,6.375889,6.5164475,6.6531014,6.79366,6.9342184,7.0747766,6.7975645,6.520352,6.2431393,5.9659266,5.688714,5.852699,6.016684,6.180669,6.348558,6.5125427,6.8795567,7.2465706,7.6135845,7.9805984,8.351517,8.062591,7.773665,7.4886436,7.1997175,6.910792,7.0903945,7.266093,7.445695,7.621393,7.800996,7.9376497,8.074304,8.210958,8.351517,8.488171,8.605303,8.722435,8.839567,8.956698,9.073831,9.468176,9.866425,10.260769,10.655114,11.0494585,9.600925,8.148487,6.699954,5.251421,3.7989833,3.2562714,2.7096553,2.1630387,1.620327,1.0737107,1.1713207,1.2650263,1.358732,1.456342,1.5500476,1.7218413,1.8897307,2.0615244,2.2294137,2.4012074,2.194274,1.9834363,1.7765031,1.5695697,1.3626363,1.1400855,0.91753453,0.6949836,0.47243267,0.24988174,0.39044023,0.5309987,0.6715572,0.80821127,0.94876975,1.3743496,1.7999294,2.2255092,2.6510892,3.076669,3.174279,3.2718892,3.3655949,3.4632049,3.5608149,3.8067923,4.0527697,4.298747,4.5408196,4.786797,5.0522966,5.3177958,5.5832953,5.8487945,6.114294,5.938596,5.7628975,5.5871997,5.4115014,5.2358036,4.60329,3.970777,3.338264,2.7057507,2.0732377,2.2489357,2.4207294,2.592523,2.7643168,2.9361105,3.767748,4.5993857,5.4271193,6.2587566,7.08649,7.363703,7.6409154,7.918128,8.1992445,8.476458,7.8478484,7.2192397,6.590631,5.9659266,5.337318,5.298274,5.263134,5.22409,5.1889505,5.1499066,5.9659266,6.785851,7.601871,8.421796,9.237816,9.296382,9.358852,9.4174185,9.475985,9.538455,9.534551,9.530646,9.530646,9.526741,9.526741,9.905469,10.284196,10.666827,11.045554,11.424281,10.756628,10.085071,9.413514,8.745861,8.074304,8.433509,8.796618,9.155824,9.515028,9.874233,10.0265045,10.178777,10.331048,10.48332,10.6355915,11.924045,13.208592,14.493141,15.77769,17.062239,17.636185,18.214037,18.787983,19.36193,19.935879,20.08815,20.244326,20.396597,20.548868,20.701141,20.002253,19.303364,18.608381,17.909492,17.210606,16.140799,15.070992,14.001186,12.93138,11.861574,11.154878,10.44818,9.741484,9.030883,8.324185,8.308568,8.296855,8.281238,8.265619,8.250002,8.827853,9.405705,9.983557,10.561408,11.139259,11.326671,11.514082,11.701493,11.888905,12.076316,12.665881,13.25935,13.852819,14.446288,15.035853,14.430671,13.821584,13.216402,12.607315,11.998228,11.342289,10.686349,10.0265045,9.370565,8.710721,8.663869,8.617016,8.570163,8.52331,8.476458,7.843944,7.211431,6.578918,5.9464045,5.3138914,5.0757227,4.841459,4.607195,4.3729305,4.138666,4.349504,4.564246,4.775084,4.985922,5.2006636,6.2938967,7.3910336,8.484266,9.581403,10.674636,11.8537655,13.028991,14.208119,15.383345,16.562475,17.546383,18.534197,19.518106,20.502016,21.485926,22.204336,22.922745,23.641155,24.355661,25.074072,22.950077,20.826082,18.698183,16.574188,14.450192,14.278399,14.11051,13.938716,13.770826,13.599033,13.239828,12.880623,12.521418,12.158309,11.799104,12.494087,13.185166,13.8762455,14.571229,15.262308,19.186234,23.114061,27.037985,30.96191,34.885834,31.949724,29.013613,26.073599,23.137487,20.201378,18.866072,17.53467,16.20327,14.871868,13.536563,13.005564,12.470661,11.939662,11.408664,10.87376,10.510651,10.151445,9.788337,9.425227,9.062118,9.069926,9.077735,9.085544,9.093353,9.101162,10.135828,11.174399,12.212971,13.251541,14.286208,12.08803,9.893755,7.6955767,5.4973984,3.2992198,2.7799344,2.260649,1.7413634,1.2181735,0.698888,0.8862993,1.0737107,1.261122,1.4485333,1.6359446,3.4710135,5.3060827,7.141152,8.976221,10.81129,13.09927,15.383345,17.66742,19.951496,22.239475,19.080814,15.926057,12.771299,9.616543,6.461786,5.6262436,4.7907014,3.959064,3.1235218,2.2879796,2.194274,2.096664,2.0029583,1.9092526,1.8116426,2.330928,2.8463092,3.3655949,3.8809757,4.4002614,4.50568,4.6150036,4.7243266,4.829746,4.939069,4.8687897,4.802415,4.73604,4.6657605,4.5993857,4.814128,5.024966,5.2358036,5.4505453,5.661383,5.423215,5.181142,4.942973,4.7009,4.462732,5.349031,6.239235,7.125534,8.011833,8.898132,7.4886436,6.0752497,4.661856,3.2484627,1.8389735,1.7023194,1.5656652,1.4329157,1.2962615,1.1635119,1.1635119,1.1635119,1.1635119,1.1635119,1.1635119,1.0463798,0.92924774,0.80821127,0.6910792,0.57394713,0.6559396,0.7418364,0.8238289,0.9058213,0.9878138,0.8316377,0.6715572,0.5153811,0.359205,0.19912452,0.1835069,0.1639849,0.14836729,0.12884527,0.113227665,0.45681506,0.79649806,1.1400855,1.4836729,1.8233559,2.0263848,2.2294137,2.4324427,2.6354716,2.8385005,3.096191,3.3538816,3.611572,3.8692627,4.126953,4.068387,4.009821,3.951255,3.8965936,3.8380275,3.4710135,3.1079042,2.7408905,2.377781,2.0107672,1.6827974,1.3509232,1.0229534,0.6910792,0.3631094,0.28892577,0.21864653,0.14446288,0.07418364,0.0,0.042948425,0.08589685,0.12884527,0.1717937,0.21083772,0.27721256,0.3435874,0.40605783,0.47243267,0.5388075,0.9019169,1.2689307,1.6320401,1.999054,2.3621633,2.0263848,1.6867018,1.3509232,1.0112402,0.6754616,0.5388075,0.40605783,0.26940376,0.13665408,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.0615244,1.9482968,1.8389735,1.7257458,1.6125181,1.4992905,2.0498111,2.6003318,3.1508527,3.7013733,4.251894,4.4119744,4.575959,4.73604,4.900025,5.0640097,5.337318,5.610626,5.8878384,6.1611466,6.4383593,6.3017054,6.1611466,6.0244927,5.8878384,5.7511845,5.22409,4.7009,4.173806,3.6506162,3.1235218,3.2367494,3.349977,3.4632049,3.5764325,3.6857557,3.6232853,3.5608149,3.4983444,3.435874,3.3734035,3.2250361,3.076669,2.9243972,2.77603,2.6237583,3.4632049,4.298747,5.138193,5.9737353,6.813182,6.8639393,6.910792,6.9615493,7.012306,7.0630636,6.813182,6.5633,6.3134184,6.0635366,5.813655,5.6730967,5.5364423,5.3997884,5.263134,5.12648,5.251421,5.376362,5.5013027,5.6262436,5.7511845,5.8761253,6.001066,6.126007,6.250948,6.375889,6.5633,6.7507114,6.9381227,7.125534,7.3129454,7.3246584,7.336372,7.348085,7.363703,7.375416,7.098203,6.824895,6.551587,6.2743745,6.001066,6.086963,6.1767645,6.262661,6.348558,6.4383593,6.899079,7.363703,7.824422,8.289046,8.749765,8.386656,8.023546,7.6643414,7.3012323,6.9381227,6.9615493,6.98888,7.012306,7.0357327,7.0630636,7.012306,6.9615493,6.910792,6.8639393,6.813182,7.0747766,7.336372,7.601871,7.8634663,8.125061,8.687295,9.249529,9.811763,10.373997,10.936231,9.187058,7.437886,5.688714,3.9356375,2.1864653,1.8858263,1.5890918,1.2884527,0.9878138,0.6871748,0.8745861,1.0619974,1.2494087,1.43682,1.6242313,1.8116426,1.999054,2.1864653,2.3738766,2.5612879,2.2255092,1.8858263,1.5500476,1.2142692,0.8745861,0.7262188,0.57394713,0.42557985,0.27330816,0.12494087,0.3357786,0.5505207,0.76135844,0.97610056,1.1869383,1.698415,2.2137961,2.7252727,3.2367494,3.7482262,3.775557,3.7989833,3.8263142,3.8497405,3.873167,4.025439,4.173806,4.3260775,4.474445,4.6267166,4.939069,5.251421,5.563773,5.8761253,6.1884775,6.0244927,5.8644123,5.700427,5.5364423,5.376362,4.6384296,3.900498,3.1625657,2.4246337,1.6867018,1.9482968,2.2137961,2.475391,2.736986,2.998581,3.5764325,4.1503797,4.7243266,5.298274,5.8761253,6.4383593,7.000593,7.562827,8.125061,8.687295,8.050878,7.4144597,6.774138,6.13772,5.5013027,5.5130157,5.5247293,5.5364423,5.548156,5.563773,6.3993154,7.238762,8.074304,8.913751,9.749292,9.850807,9.948417,10.049932,10.151445,10.249056,10.174872,10.100689,10.0265045,9.948417,9.874233,10.350571,10.826907,11.29934,11.775677,12.24811,11.525795,10.799577,10.073358,9.351044,8.624825,8.800523,8.976221,9.151918,9.323712,9.499411,9.987461,10.475512,10.963562,11.4516115,11.935758,13.337439,14.739119,16.136894,17.538574,18.936352,19.549341,20.162333,20.775324,21.388315,22.001307,22.1731,22.348799,22.524496,22.700195,22.875893,22.223858,21.575727,20.92369,20.27556,19.623526,18.276506,16.925583,15.57466,14.223738,12.8767185,12.138786,11.400854,10.662923,9.924991,9.187058,9.112875,9.0386915,8.960603,8.886419,8.812236,9.612638,10.413041,11.213444,12.013845,12.814248,12.911859,13.013372,13.110983,13.212498,13.314012,14.126127,14.938243,15.750359,16.562475,17.37459,16.69913,16.023666,15.348206,14.676648,14.001186,13.189071,12.376955,11.560935,10.748819,9.936704,9.948417,9.964035,9.975748,9.987461,9.999174,9.261242,8.52331,7.7892823,7.0513506,6.3134184,5.8761253,5.4388323,5.001539,4.564246,4.123049,4.173806,4.224563,4.2753205,4.3260775,4.376835,5.5989127,6.824895,8.050878,9.276859,10.498938,11.799104,13.09927,14.399435,15.699601,16.999767,17.936825,18.87388,19.810938,20.751898,21.688955,22.78609,23.887133,24.988174,26.089216,27.186354,24.476698,21.763138,19.049578,16.33602,13.626364,13.774731,13.923099,14.07537,14.223738,14.376009,14.313539,14.251068,14.188598,14.126127,14.063657,14.551707,15.035853,15.523903,16.011953,16.500004,20.76361,25.023314,29.28692,33.55053,37.814137,34.612526,31.410915,28.213211,25.0116,21.813896,20.45126,19.088623,17.725986,16.36335,15.000713,14.161267,13.325725,12.486279,11.650736,10.81129,10.748819,10.686349,10.6238785,10.561408,10.498938,10.413041,10.323239,10.237343,10.151445,10.061645,10.436467,10.81129,11.186112,11.560935,11.935758,10.100689,8.261715,6.426646,4.5876727,2.7486992,2.3621633,1.9756275,1.5890918,1.1986516,0.81211567,0.8628729,0.9136301,0.96438736,1.0112402,1.0619974,3.474918,5.8878384,8.300759,10.71368,13.1266,15.664462,18.19842,20.73628,23.274141,25.812004,22.200432,18.58886,14.973383,11.361811,7.7502384,6.461786,5.173333,3.8887846,2.6003318,1.3118792,1.2494087,1.1869383,1.1244678,1.0619974,0.999527,1.8233559,2.6510892,3.474918,4.298747,5.12648,5.2865605,5.4505453,5.610626,5.774611,5.938596,5.688714,5.4388323,5.1889505,4.939069,4.689187,4.7126136,4.73604,4.7633705,4.786797,4.814128,4.6735697,4.5369153,4.4002614,4.263607,4.123049,5.138193,6.1494336,7.1606736,8.175818,9.187058,7.648724,6.114294,4.575959,3.0376248,1.4992905,1.33921,1.175225,1.0112402,0.8511597,0.6871748,0.63641757,0.58566034,0.5388075,0.48805028,0.43729305,0.46071947,0.48805028,0.5114767,0.5388075,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.0,0.0,0.0,0.0,0.0,0.41386664,0.8238289,1.2376955,1.6515622,2.0615244,2.2372224,2.4129205,2.5886188,2.7643168,2.9361105,3.2250361,3.513962,3.7989833,4.087909,4.376835,4.087909,3.7989833,3.513962,3.2250361,2.9361105,2.6003318,2.260649,1.9248703,1.5890918,1.2494087,1.0893283,0.92534333,0.76135844,0.60127795,0.43729305,0.3513962,0.26159495,0.1756981,0.08589685,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.31235218,0.37482262,0.43729305,0.4997635,0.5622339,0.97610056,1.3860629,1.7999294,2.2137961,2.6237583,2.260649,1.901444,1.5383345,1.175225,0.81211567,0.6481308,0.48805028,0.3240654,0.1639849,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.7882162,1.6710842,1.5578566,1.4407244,1.3274968,1.2142692,1.6593709,2.1005683,2.5456703,2.9907722,3.435874,3.5764325,3.716991,3.8575494,3.998108,4.138666,4.4393053,4.73604,5.036679,5.337318,5.6379566,5.700427,5.7628975,5.825368,5.8878384,5.950309,5.5169206,5.083532,4.6540475,4.220659,3.78727,3.8965936,4.0020123,4.1113358,4.2167544,4.3260775,4.2167544,4.1035266,3.9942036,3.8848803,3.775557,3.513962,3.2484627,2.9868677,2.7252727,2.463678,3.2250361,3.9863946,4.7516575,5.5130157,6.2743745,6.3407493,6.4032197,6.4695945,6.5359693,6.5984397,6.4149327,6.2314262,6.044015,5.860508,5.6730967,5.5442514,5.4154058,5.2865605,5.153811,5.024966,5.1108627,5.196759,5.278752,5.364649,5.4505453,5.6340523,5.813655,5.997162,6.180669,6.364176,6.551587,6.7389984,6.9264097,7.113821,7.3012323,7.2934237,7.289519,7.2856145,7.28171,7.2739015,7.0357327,6.79366,6.5554914,6.3134184,6.0752497,6.165051,6.2548523,6.3446536,6.434455,6.524256,6.9342184,7.3402762,7.746334,8.156297,8.562354,8.312472,8.062591,7.812709,7.562827,7.3129454,7.348085,7.3832245,7.4183645,7.453504,7.4886436,7.3988423,7.309041,7.2192397,7.1294384,7.0357327,7.328563,7.621393,7.914223,8.207053,8.499884,8.683391,8.870802,9.054309,9.24172,9.425227,7.9337454,6.4383593,4.9468775,3.455396,1.9639144,1.717937,1.4719596,1.2259823,0.98390937,0.737932,0.9136301,1.0932326,1.2689307,1.4485333,1.6242313,1.7413634,1.8545911,1.9717231,2.084951,2.1981785,1.9053483,1.6086137,1.3157835,1.0190489,0.7262188,0.62860876,0.5309987,0.43338865,0.3357786,0.23816854,0.39824903,0.5622339,0.7262188,0.8862993,1.0502841,1.4407244,1.8311646,2.2216048,2.6081407,2.998581,3.018103,3.0415294,3.0610514,3.0805733,3.1000953,3.2914112,3.4866312,3.677947,3.8692627,4.0605783,4.298747,4.533011,4.7672753,5.001539,5.2358036,5.1616197,5.087436,5.0132523,4.939069,4.860981,4.2440853,3.6271896,3.0102942,2.3933985,1.7765031,2.0654287,2.3543546,2.6432803,2.9361105,3.2250361,3.8770714,4.5291066,5.181142,5.833177,6.4891167,6.9810715,7.473026,7.9649806,8.456935,8.94889,8.339804,7.7307167,7.1216297,6.5086384,5.899552,5.708236,5.520825,5.3295093,5.138193,4.950782,5.6418614,6.336845,7.027924,7.719003,8.413987,8.495979,8.581876,8.667773,8.75367,8.835662,8.741957,8.648251,8.550641,8.456935,8.36323,8.886419,9.405705,9.928895,10.452085,10.975275,10.409137,9.839094,9.272955,8.706817,8.136774,8.253906,8.367134,8.484266,8.597494,8.710721,9.339331,9.967939,10.596548,11.221252,11.849861,13.427239,15.004618,16.581997,18.159374,19.736753,20.494207,21.247757,22.001307,22.75876,23.51231,23.793427,24.07845,24.359566,24.640682,24.925705,24.156536,23.383465,22.614298,21.84513,21.075964,19.646952,18.221846,16.792833,15.363823,13.938716,13.232019,12.521418,11.814721,11.108025,10.401327,10.323239,10.2451515,10.167064,10.088976,10.010887,10.6355915,11.256392,11.881096,12.501896,13.1266,13.138313,13.153932,13.169549,13.185166,13.200784,13.954333,14.711788,15.465338,16.218887,16.976341,16.55857,16.140799,15.723028,15.305257,14.8874855,13.993378,13.09927,12.201257,11.307149,10.413041,10.241247,10.073358,9.901564,9.733675,9.561881,8.917655,8.273428,7.629202,6.9810715,6.336845,6.0205884,5.704332,5.3841705,5.067914,4.7516575,4.7243266,4.7009,4.6735697,4.650143,4.6267166,5.7394714,6.8561306,7.968885,9.085544,10.198298,11.478943,12.755682,14.032422,15.309161,16.585901,17.558098,18.534197,19.506393,20.47859,21.450787,22.40346,23.356134,24.30881,25.261482,26.214157,24.211199,22.20824,20.205282,18.202324,16.199366,15.828446,15.461433,15.090515,14.719597,14.348679,14.438479,14.528281,14.618082,14.711788,14.801589,15.035853,15.274021,15.51219,15.750359,15.988527,20.138906,24.29319,28.443571,32.597855,36.748234,34.573483,32.394825,30.21617,28.041416,25.86276,24.543072,23.223385,21.903696,20.58401,19.26432,18.42878,17.597141,16.765503,15.933866,15.098324,14.450192,13.802062,13.150026,12.501896,11.849861,11.361811,10.869856,10.381805,9.889851,9.4018,9.511124,9.620447,9.729771,9.839094,9.948417,8.398369,6.8483214,5.298274,3.7482262,2.1981785,1.893635,1.5890918,1.2845483,0.98000497,0.6754616,0.737932,0.80040246,0.8628729,0.92534333,0.9878138,4.041056,7.098203,10.151445,13.208592,16.261835,18.627903,20.99397,23.356134,25.722202,28.08827,24.340044,20.591818,16.843592,13.09927,9.351044,8.304664,7.2582836,6.2158084,5.169429,4.126953,4.0644827,4.0059166,3.9434462,3.8848803,3.8263142,4.3338866,4.841459,5.349031,5.8566036,6.364176,6.2587566,6.1572423,6.055728,5.9542136,5.8487945,5.563773,5.2748475,4.985922,4.7009,4.4119744,4.3534083,4.290938,4.2323723,4.173806,4.1113358,4.173806,4.2362766,4.298747,4.3612175,4.423688,5.036679,5.645766,6.2548523,6.8639393,7.473026,6.2431393,5.0132523,3.7833657,2.5534792,1.3235924,1.2337911,1.1439898,1.0541886,0.96438736,0.8745861,0.8628729,0.8511597,0.8394465,0.8238289,0.81211567,0.8784905,0.94096094,1.0073358,1.0737107,1.1361811,1.077615,1.0190489,0.95657855,0.8980125,0.8394465,0.6871748,0.5388075,0.38653582,0.23816854,0.08589685,0.10932326,0.12884527,0.14836729,0.1678893,0.18741131,0.48414588,0.78088045,1.0815194,1.3782539,1.6749885,1.9482968,2.2216048,2.4910088,2.7643168,3.0376248,3.154757,3.2718892,3.3890212,3.506153,3.6232853,3.435874,3.2484627,3.0610514,2.87364,2.6862288,2.358259,2.0263848,1.698415,1.3665408,1.038571,0.9019169,0.76135844,0.62470436,0.48805028,0.3513962,0.30063897,0.25378615,0.20693332,0.16008049,0.113227665,0.16008049,0.20693332,0.25378615,0.30063897,0.3513962,0.42557985,0.4997635,0.57394713,0.6481308,0.7262188,1.0502841,1.3743496,1.698415,2.0263848,2.35045,2.0459068,1.7452679,1.4407244,1.1400855,0.8394465,0.6910792,0.5427119,0.39434463,0.24597734,0.10151446,0.093705654,0.08980125,0.08589685,0.078088045,0.07418364,0.06637484,0.05466163,0.046852827,0.03513962,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.023426414,0.019522011,0.015617609,0.015617609,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.5110037,1.3938715,1.2767396,1.1596074,1.0424755,0.92534333,1.2650263,1.6047094,1.9443923,2.2840753,2.6237583,2.7408905,2.8619268,2.979059,3.096191,3.213323,3.5373883,3.8614538,4.1894236,4.513489,4.8375545,5.099149,5.3607445,5.6262436,5.8878384,6.1494336,5.8097506,5.4700675,5.1303844,4.7907014,4.4510183,4.552533,4.6540475,4.755562,4.860981,4.9624953,4.806319,4.646239,4.4900627,4.3338866,4.173806,3.7989833,3.4241607,3.049338,2.6745155,2.2996929,2.9868677,3.6740425,4.3612175,5.0483923,5.735567,5.8175592,5.8956475,5.9776397,6.055728,6.13772,6.016684,5.8956475,5.7785153,5.657479,5.5364423,5.4154058,5.2943697,5.169429,5.0483923,4.9234514,4.970304,5.0132523,5.0601053,5.1069584,5.1499066,5.388075,5.630148,5.8683167,6.1103897,6.348558,6.5359693,6.7233806,6.910792,7.098203,7.2856145,7.266093,7.2426662,7.2192397,7.195813,7.1762915,6.969358,6.7663293,6.559396,6.356367,6.1494336,6.2431393,6.336845,6.426646,6.520352,6.6140575,6.9654536,7.3168497,7.6682463,8.023546,8.374943,8.238289,8.101635,7.9610763,7.824422,7.687768,7.7307167,7.7775693,7.824422,7.8673706,7.914223,7.7814736,7.6526284,7.523783,7.3910336,7.262188,7.5862536,7.9064145,8.23048,8.550641,8.874706,8.683391,8.488171,8.296855,8.105539,7.914223,6.676528,5.4427366,4.2089458,2.97125,1.737459,1.5461433,1.358732,1.1674163,0.97610056,0.78868926,0.95657855,1.1205635,1.2884527,1.456342,1.6242313,1.6671798,1.7101282,1.7530766,1.796025,1.8389735,1.5851873,1.3314011,1.0815194,0.8277333,0.57394713,0.5309987,0.48414588,0.44119745,0.39434463,0.3513962,0.46071947,0.57394713,0.6871748,0.80040246,0.9136301,1.1791295,1.4485333,1.7140326,1.9834363,2.2489357,2.2645533,2.280171,2.2957885,2.3114061,2.3231194,2.5612879,2.795552,3.0298162,3.2640803,3.4983444,3.6584249,3.814601,3.970777,4.1308575,4.2870336,4.298747,4.3143644,4.3260775,4.337791,4.349504,3.853645,3.3538816,2.8580225,2.358259,1.8623998,2.1786566,2.4988174,2.815074,3.1313305,3.4514916,4.181615,4.911738,5.6418614,6.36808,7.098203,7.523783,7.9454584,8.367134,8.78881,9.21439,8.628729,8.046973,7.465217,6.883461,6.3017054,5.9073606,5.5169206,5.1225758,4.728231,4.337791,4.884407,5.4310236,5.9815445,6.5281606,7.0747766,7.1450562,7.2153354,7.2856145,7.355894,7.426173,7.309041,7.195813,7.0786815,6.9654536,6.8483214,7.4183645,7.988407,8.55845,9.128492,9.698535,9.288573,8.878611,8.468649,8.058686,7.648724,7.703386,7.7619514,7.816613,7.871275,7.9259367,8.691199,9.460366,10.22563,10.994797,11.763964,13.51704,15.274021,17.027098,18.784079,20.537155,21.43517,22.333181,23.231194,24.129206,25.023314,25.413754,25.804195,26.194635,26.585075,26.975515,26.085312,25.195108,24.304905,23.4147,22.524496,21.021301,19.514202,18.011007,16.503908,15.000713,14.321347,13.645885,12.96652,12.291059,11.611692,11.533605,11.4516115,11.373524,11.291532,11.213444,11.6585455,12.103647,12.548749,12.993851,13.438952,13.368673,13.298394,13.228115,13.157836,13.087557,13.786445,14.481428,15.180316,15.879204,16.574188,16.414106,16.254026,16.093946,15.933866,15.773785,14.797685,13.821584,12.841579,11.8654785,10.889378,10.534078,10.182681,9.8312845,9.475985,9.124588,8.574067,8.019642,7.4691215,6.914696,6.364176,6.165051,5.9659266,5.7707067,5.571582,5.376362,5.2748475,5.173333,5.0757227,4.9742084,4.8765984,5.8800297,6.883461,7.890797,8.894228,9.901564,11.154878,12.408191,13.665408,14.918721,16.175938,17.183275,18.19061,19.197947,20.205282,21.212618,22.016924,22.821232,23.629442,24.43375,25.238056,23.9457,22.653341,21.360985,20.068628,18.77627,17.886066,16.995863,16.10566,15.215456,14.325252,14.567325,14.809398,15.051471,15.293544,15.535617,15.523903,15.51219,15.500477,15.488764,15.473146,19.518106,23.559164,27.604124,31.64518,35.686237,34.530533,33.378735,32.22303,31.06733,29.911625,28.634886,27.358147,26.081408,24.800762,23.524023,22.696291,21.868557,21.040823,20.21309,19.389261,18.151566,16.91387,15.676175,14.438479,13.200784,12.306676,11.416472,10.522364,9.628256,8.738052,8.581876,8.4257,8.273428,8.117252,7.9610763,6.699954,5.4388323,4.173806,2.912684,1.6515622,1.4290112,1.2064602,0.98390937,0.76135844,0.5388075,0.61299115,0.6871748,0.76135844,0.8394465,0.9136301,4.6110992,8.308568,12.006037,15.7035055,19.400974,21.591345,23.785618,25.975988,28.170261,30.360632,26.479656,22.59868,18.7138,14.832824,10.951848,10.147541,9.343235,8.542832,7.7385254,6.9381227,6.8795567,6.8209906,6.7663293,6.707763,6.649197,6.8405128,7.0318284,7.2192397,7.4105554,7.601871,7.230953,6.8639393,6.4969254,6.1299114,5.7628975,5.4388323,5.1108627,4.786797,4.462732,4.138666,3.9942036,3.8458362,3.7013733,3.5569105,3.4124475,3.6740425,3.9356375,4.2011366,4.462732,4.7243266,4.93126,5.138193,5.349031,5.5559645,5.7628975,4.841459,3.9161155,2.9946766,2.0732377,1.1517987,1.1322767,1.116659,1.097137,1.0815194,1.0619974,1.0893283,1.1127546,1.1361811,1.1635119,1.1869383,1.2923572,1.397776,1.5031948,1.6086137,1.7140326,1.5929961,1.4719596,1.3509232,1.2337911,1.1127546,0.92534333,0.737932,0.5505207,0.3631094,0.1756981,0.21474212,0.25378615,0.29673457,0.3357786,0.37482262,0.5583295,0.7418364,0.92143893,1.1049459,1.2884527,1.6593709,2.0263848,2.397303,2.7682211,3.1391394,3.084478,3.0337205,2.979059,2.9283018,2.87364,2.787743,2.7018464,2.612045,2.5261483,2.436347,2.1161861,1.7921207,1.4680552,1.1478943,0.8238289,0.7106012,0.60127795,0.48805028,0.37482262,0.26159495,0.25378615,0.24597734,0.23816854,0.23426414,0.22645533,0.26940376,0.31625658,0.359205,0.40605783,0.44900626,0.5388075,0.62470436,0.7106012,0.80040246,0.8862993,1.1244678,1.3626363,1.6008049,1.8389735,2.0732377,1.8311646,1.5890918,1.3470187,1.1049459,0.8628729,0.7301232,0.59737355,0.46462387,0.3318742,0.19912452,0.1756981,0.15617609,0.13274968,0.10932326,0.08589685,0.078088045,0.07418364,0.06637484,0.058566034,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.046852827,0.039044023,0.03513962,0.031235218,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.2376955,1.116659,0.9956226,0.8784905,0.75745404,0.63641757,0.8706817,1.1088502,1.3431144,1.5773785,1.8116426,1.9092526,2.0029583,2.096664,2.194274,2.2879796,2.639376,2.9868677,3.338264,3.6857557,4.037152,4.5017757,4.9624953,5.423215,5.8878384,6.348558,6.1025805,5.8566036,5.606722,5.3607445,5.1108627,5.2084727,5.3060827,5.4036927,5.5013027,5.5989127,5.395884,5.1889505,4.985922,4.7789884,4.575959,4.087909,3.5998588,3.1118085,2.6237583,2.135708,2.7486992,3.3616903,3.9746814,4.5876727,5.2006636,5.2943697,5.388075,5.4856853,5.579391,5.6730967,5.618435,5.563773,5.5091114,5.45445,5.3997884,5.2865605,5.169429,5.056201,4.939069,4.825841,4.829746,4.83365,4.841459,4.845363,4.8492675,5.1460023,5.446641,5.743376,6.04011,6.336845,6.524256,6.7116675,6.899079,7.08649,7.2739015,7.2348576,7.195813,7.1567693,7.113821,7.0747766,6.9068875,6.735094,6.5633,6.395411,6.223617,6.321227,6.4149327,6.5086384,6.606249,6.699954,6.996689,7.2934237,7.5940623,7.890797,8.187531,8.164105,8.136774,8.113348,8.086017,8.062591,8.117252,8.171914,8.226576,8.281238,8.335898,8.16801,7.996216,7.8283267,7.656533,7.4886436,7.8400397,8.191436,8.546737,8.898132,9.249529,8.679486,8.109444,7.5394006,6.969358,6.3993154,5.423215,4.4432096,3.4671092,2.4910088,1.5110037,1.3782539,1.2415999,1.1088502,0.97219616,0.8394465,0.9956226,1.1517987,1.3118792,1.4680552,1.6242313,1.5969005,1.5656652,1.53443,1.5031948,1.475864,1.2650263,1.0541886,0.8433509,0.63641757,0.42557985,0.43338865,0.44119745,0.44900626,0.45681506,0.46071947,0.5231899,0.58566034,0.6481308,0.7106012,0.77307165,0.92143893,1.0659018,1.2103647,1.3548276,1.4992905,1.5110037,1.5188124,1.5305257,1.5383345,1.5500476,1.8272603,2.1044729,2.3816853,2.6588979,2.9361105,3.018103,3.096191,3.1781836,3.2562714,3.338264,3.435874,3.5373883,3.638903,3.736513,3.8380275,3.4593005,3.0805733,2.7057507,2.3270237,1.9482968,2.2957885,2.639376,2.9868677,3.330455,3.6740425,4.482254,5.290465,6.098676,6.9068875,7.7111945,8.066495,8.4178915,8.769287,9.120684,9.475985,8.921559,8.36323,7.8088045,7.2543793,6.699954,6.1064854,5.5091114,4.9156423,4.318269,3.7247996,4.126953,4.5291066,4.93126,5.3334136,5.735567,5.794133,5.8487945,5.903456,5.958118,6.012779,5.8761253,5.743376,5.606722,5.473972,5.337318,5.9542136,6.571109,7.191909,7.8088045,8.4257,8.171914,7.918128,7.6682463,7.4144597,7.1606736,7.1567693,7.152865,7.1489606,7.141152,7.137247,8.043069,8.952794,9.858616,10.768341,11.674163,13.606842,15.539521,17.4722,19.404879,21.337559,22.37613,23.418604,24.457176,25.495747,26.538221,27.03408,27.533844,28.029703,28.529467,29.025326,28.014086,27.00675,25.99551,24.98427,23.976934,22.391747,20.810465,19.229181,17.643993,16.062712,15.41458,14.766449,14.118319,13.4740925,12.825961,12.743969,12.661977,12.576079,12.494087,12.412095,12.681499,12.946998,13.216402,13.481901,13.751305,13.595129,13.438952,13.286681,13.130505,12.974329,13.614651,14.254972,14.895294,15.535617,16.175938,16.273548,16.371159,16.46877,16.56638,16.663988,15.601992,14.543899,13.481901,12.423808,11.361811,10.826907,10.292005,9.757101,9.2221985,8.687295,8.226576,7.7658563,7.309041,6.8483214,6.387602,6.309514,6.2314262,6.153338,6.0791545,6.001066,5.825368,5.64967,5.473972,5.298274,5.12648,6.0205884,6.914696,7.8088045,8.706817,9.600925,10.8308115,12.064603,13.298394,14.528281,15.762072,16.804546,17.847023,18.889498,19.931974,20.97445,21.634293,22.290232,22.946173,23.606016,24.261955,23.6802,23.098444,22.516687,21.931028,21.349272,19.939783,18.530293,17.120804,15.711315,14.301826,14.69617,15.090515,15.484859,15.879204,16.273548,16.011953,15.750359,15.488764,15.223265,14.96167,18.893402,22.82904,26.760773,30.692507,34.62424,34.49149,34.35874,34.22599,34.09324,33.964394,32.7267,31.492908,30.259117,29.021421,27.78763,26.963802,26.143877,25.32005,24.49622,23.676296,21.849035,20.025679,18.19842,16.375063,14.551707,13.2554455,11.959184,10.666827,9.370565,8.074304,7.656533,7.2348576,6.813182,6.395411,5.9737353,5.001539,4.025439,3.049338,2.0732377,1.1010414,0.96048295,0.8199245,0.679366,0.5388075,0.39824903,0.48805028,0.57394713,0.6637484,0.74964523,0.8394465,5.1772375,9.518932,13.856724,18.19842,22.53621,24.558691,26.577267,28.595842,30.618322,32.636898,28.619268,24.601639,20.58401,16.56638,12.548749,11.990419,11.428185,10.869856,10.311526,9.749292,9.694631,9.639969,9.585307,9.530646,9.475985,9.347139,9.218294,9.093353,8.964508,8.835662,8.203149,7.570636,6.9381227,6.3056097,5.6730967,5.3138914,4.950782,4.5876727,4.224563,3.8614538,3.631094,3.4007344,3.174279,2.9439192,2.7135596,3.174279,3.638903,4.0996222,4.564246,5.024966,4.829746,4.6345253,4.4393053,4.2440853,4.0488653,3.435874,2.8189783,2.2059872,1.5890918,0.97610056,1.0307622,1.0854238,1.1400855,1.1947471,1.2494087,1.3118792,1.3743496,1.43682,1.4992905,1.5617609,1.7062237,1.8506867,1.999054,2.1435168,2.2879796,2.1083772,1.9287747,1.7491722,1.5656652,1.3860629,1.1635119,0.93705654,0.7106012,0.48805028,0.26159495,0.3240654,0.38263142,0.44119745,0.5036679,0.5622339,0.62860876,0.698888,0.76526284,0.8316377,0.9019169,1.3665408,1.8350691,2.3035975,2.7682211,3.2367494,3.0141985,2.7916477,2.5690966,2.3465457,2.1239948,2.135708,2.1513257,2.1630387,2.174752,2.1864653,1.8741131,1.5578566,1.2415999,0.92924774,0.61299115,0.5231899,0.43729305,0.3513962,0.26159495,0.1756981,0.20693332,0.23816854,0.27330816,0.30454338,0.3357786,0.37872702,0.42167544,0.46462387,0.5075723,0.5505207,0.6481308,0.74964523,0.8511597,0.94876975,1.0502841,1.1986516,1.3509232,1.4992905,1.6515622,1.7999294,1.6164225,1.43682,1.2533131,1.0698062,0.8862993,0.76916724,0.6520352,0.5349031,0.41777104,0.30063897,0.26159495,0.21864653,0.1796025,0.14055848,0.10151446,0.093705654,0.08980125,0.08589685,0.078088045,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.96438736,0.8394465,0.71841,0.59346914,0.47243267,0.3513962,0.48024148,0.60908675,0.7418364,0.8706817,0.999527,1.0737107,1.1439898,1.2181735,1.2884527,1.3626363,1.737459,2.1122816,2.4871042,2.8619268,3.2367494,3.900498,4.564246,5.22409,5.8878384,6.551587,6.395411,6.239235,6.083059,5.930787,5.774611,5.8683167,5.958118,6.0518236,6.1455293,6.239235,5.985449,5.7316628,5.481781,5.2279944,4.9742084,4.376835,3.775557,3.174279,2.5769055,1.9756275,2.514435,3.049338,3.5881457,4.126953,4.661856,4.7711797,4.884407,4.9937305,5.1030536,5.212377,5.22409,5.2318993,5.2436123,5.251421,5.263134,5.153811,5.0483923,4.939069,4.83365,4.7243266,4.689187,4.6540475,4.618908,4.5837684,4.548629,4.903929,5.2592297,5.6145306,5.969831,6.3251314,6.5125427,6.699954,6.8873653,7.0747766,7.262188,7.2036223,7.1489606,7.0903945,7.0318284,6.9732623,6.8405128,6.703859,6.571109,6.434455,6.3017054,6.3993154,6.4969254,6.590631,6.688241,6.785851,7.0318284,7.2739015,7.5159745,7.758047,8.00012,8.086017,8.175818,8.261715,8.351517,8.437413,8.503788,8.566258,8.632633,8.699008,8.761478,8.550641,8.343708,8.13287,7.9220324,7.7111945,8.093826,8.476458,8.859089,9.24172,9.6243515,8.675582,7.7307167,6.7819467,5.833177,4.8883114,4.165997,3.4475873,2.7291772,2.0068626,1.2884527,1.2064602,1.1283722,1.0463798,0.96829176,0.8862993,1.0346665,1.183034,1.3314011,1.475864,1.6242313,1.5227169,1.4212024,1.3157835,1.2142692,1.1127546,0.94486535,0.77697605,0.60908675,0.44119745,0.27330816,0.3357786,0.39434463,0.45681506,0.5153811,0.57394713,0.58566034,0.60127795,0.61299115,0.62470436,0.63641757,0.659844,0.6832704,0.7066968,0.7262188,0.74964523,0.75354964,0.76135844,0.76526284,0.76916724,0.77307165,1.0932326,1.4133936,1.7335546,2.0537157,2.3738766,2.377781,2.3816853,2.3816853,2.3855898,2.3855898,2.5769055,2.7643168,2.951728,3.1391394,3.3265507,3.06886,2.8111696,2.5534792,2.2957885,2.0380979,2.4090161,2.7838387,3.154757,3.5256753,3.900498,4.786797,5.6691923,6.5554914,7.4417906,8.324185,8.609207,8.890324,9.171441,9.456462,9.737579,9.2104845,8.683391,8.156297,7.629202,7.098203,6.3017054,5.505207,4.7087092,3.9083066,3.1118085,3.3694992,3.6271896,3.8848803,4.142571,4.4002614,4.4393053,4.478349,4.521298,4.560342,4.5993857,4.4432096,4.290938,4.134762,3.978586,3.8263142,4.4900627,5.153811,5.8214636,6.4852123,7.1489606,7.055255,6.9615493,6.8639393,6.7702336,6.676528,6.610153,6.5437784,6.481308,6.4149327,6.348558,7.3988423,8.445222,9.491602,10.541886,11.588266,13.696643,15.808925,17.917301,20.025679,22.13796,23.320995,24.504028,25.683159,26.866192,28.049225,28.654408,29.25959,29.864773,30.469955,31.075138,29.946766,28.81449,27.686117,26.55384,25.425468,23.766096,22.106726,20.44345,18.784079,17.124708,16.507812,15.890917,15.274021,14.653222,14.036326,13.954333,13.868437,13.78254,13.696643,13.610746,13.704452,13.794253,13.884054,13.973856,14.063657,13.821584,13.583415,13.341343,13.103174,12.861101,13.446761,14.028518,14.610273,15.192029,15.773785,16.129086,16.484386,16.839687,17.194988,17.550287,16.406298,15.266212,14.122223,12.978233,11.838148,11.119738,10.401327,9.686822,8.968412,8.250002,7.882988,7.5159745,7.1489606,6.7780423,6.4110284,6.453977,6.4969254,6.5398736,6.5828223,6.6257706,6.375889,6.126007,5.8761253,5.6262436,5.376362,6.1611466,6.9459314,7.7307167,8.515501,9.300286,10.510651,11.721016,12.93138,14.141745,15.348206,16.42582,17.503435,18.58105,19.658665,20.73628,21.247757,21.759233,22.266806,22.778282,23.285854,23.4147,23.543545,23.668486,23.79733,23.926178,21.993498,20.064724,18.135948,16.20327,14.274494,14.821111,15.371632,15.918248,16.464865,17.01148,16.500004,15.988527,15.473146,14.96167,14.450192,18.272602,22.095013,25.917421,29.739832,33.56224,34.452446,35.342648,36.232853,37.12306,38.01326,36.818512,35.62767,34.43683,33.24208,32.05124,31.231314,30.415293,29.599274,28.779348,27.96333,25.550407,23.137487,20.724567,18.311647,15.8987255,14.204215,12.5058,10.807385,9.108971,7.4105554,6.727285,6.044015,5.35684,4.6735697,3.9863946,3.2992198,2.612045,1.9248703,1.2376955,0.5505207,0.49195468,0.43338865,0.37872702,0.32016098,0.26159495,0.3631094,0.46071947,0.5622339,0.6637484,0.76135844,5.743376,10.729298,15.711315,20.693333,25.67535,27.522131,29.368914,31.215696,33.066383,34.913166,30.75888,26.608501,22.454218,18.303837,14.149553,13.833297,13.513136,13.196879,12.880623,12.564366,12.509705,12.458947,12.404286,12.353529,12.298867,11.8537655,11.408664,10.963562,10.518459,10.073358,9.17925,8.281238,7.3832245,6.4852123,5.5871997,5.1889505,4.786797,4.388548,3.9863946,3.5881457,3.2718892,2.9556324,2.6432803,2.3270237,2.0107672,2.6745155,3.338264,3.998108,4.661856,5.3256044,4.728231,4.1308575,3.533484,2.9361105,2.338737,2.0302892,1.7218413,1.4133936,1.1088502,0.80040246,0.92924774,1.0541886,1.183034,1.3118792,1.43682,1.5383345,1.6359446,1.737459,1.8389735,1.9365835,2.1239948,2.3075018,2.4910088,2.67842,2.8619268,2.6237583,2.3816853,2.1435168,1.901444,1.6632754,1.4016805,1.1361811,0.8745861,0.61299115,0.3513962,0.42948425,0.5114767,0.58956474,0.6715572,0.74964523,0.7027924,0.6559396,0.60908675,0.5583295,0.5114767,1.077615,1.6437533,2.2059872,2.7721257,3.338264,2.9439192,2.5534792,2.1591344,1.7686942,1.3743496,1.4875772,1.6008049,1.7140326,1.8233559,1.9365835,1.6281357,1.3235924,1.0151446,0.7066968,0.39824903,0.3357786,0.27330816,0.21083772,0.14836729,0.08589685,0.16008049,0.23426414,0.30454338,0.37872702,0.44900626,0.49195468,0.5309987,0.5700427,0.60908675,0.6481308,0.76135844,0.8745861,0.9878138,1.1010414,1.2142692,1.2767396,1.33921,1.4016805,1.4641509,1.5266213,1.4016805,1.2806439,1.1557031,1.0346665,0.9136301,0.80821127,0.7066968,0.60518235,0.5036679,0.39824903,0.3435874,0.28502136,0.22645533,0.1717937,0.113227665,0.10932326,0.10932326,0.10541886,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.08980125,0.078088045,0.07027924,0.058566034,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6871748,0.5622339,0.43729305,0.31235218,0.18741131,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.23816854,0.28892577,0.3357786,0.38653582,0.43729305,0.8355421,1.2376955,1.6359446,2.0380979,2.436347,3.2992198,4.1620927,5.024966,5.8878384,6.7507114,6.688241,6.6257706,6.5633,6.5008297,6.4383593,6.524256,6.6140575,6.699954,6.785851,6.8756523,6.575013,6.2743745,5.9737353,5.6730967,5.376362,4.661856,3.951255,3.2367494,2.5261483,1.8116426,2.2762666,2.736986,3.2016098,3.6623292,4.123049,4.251894,4.376835,4.5017757,4.6267166,4.7516575,4.825841,4.900025,4.9742084,5.0483923,5.12648,5.024966,4.9234514,4.825841,4.7243266,4.6267166,4.548629,4.474445,4.4002614,4.3260775,4.251894,4.661856,5.0757227,5.4856853,5.899552,6.3134184,6.5008297,6.688241,6.8756523,7.0630636,7.250475,7.1762915,7.098203,7.0240197,6.949836,6.8756523,6.774138,6.676528,6.575013,6.473499,6.375889,6.473499,6.575013,6.676528,6.774138,6.8756523,7.0630636,7.250475,7.437886,7.6252975,7.812709,8.011833,8.210958,8.413987,8.6131115,8.812236,8.886419,8.960603,9.0386915,9.112875,9.187058,8.937177,8.687295,8.437413,8.187531,7.9376497,8.351517,8.761478,9.175345,9.589212,9.999174,8.675582,7.3519893,6.0244927,4.7009,3.3734035,2.912684,2.4519646,1.9873407,1.5266213,1.0619974,1.038571,1.0112402,0.9878138,0.96438736,0.93705654,1.0737107,1.2142692,1.3509232,1.4875772,1.6242313,1.4485333,1.2767396,1.1010414,0.92534333,0.74964523,0.62470436,0.4997635,0.37482262,0.24988174,0.12494087,0.23816854,0.3513962,0.46071947,0.57394713,0.6871748,0.6481308,0.61299115,0.57394713,0.5388075,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.0,0.0,0.0,0.0,0.0,0.0,0.3631094,0.7262188,1.0893283,1.4485333,1.8116426,1.737459,1.6632754,1.5890918,1.5110037,1.43682,1.7140326,1.9873407,2.260649,2.5378613,2.8111696,2.6745155,2.5378613,2.4012074,2.260649,2.1239948,2.5261483,2.9243972,3.3265507,3.7247996,4.123049,5.087436,6.0518236,7.012306,7.9766936,8.937177,9.151918,9.362757,9.573594,9.788337,9.999174,9.499411,8.999647,8.499884,8.00012,7.5003567,6.5008297,5.5013027,4.5017757,3.4983444,2.4988174,2.612045,2.7252727,2.8385005,2.951728,3.0610514,3.0883822,3.1118085,3.1391394,3.1625657,3.1859922,3.0141985,2.8385005,2.6628022,2.4871042,2.3114061,3.0259118,3.736513,4.4510183,5.1616197,5.8761253,5.938596,6.001066,6.0635366,6.126007,6.1884775,6.0635366,5.938596,5.813655,5.688714,5.563773,6.7507114,7.9376497,9.124588,10.311526,11.498465,13.786445,16.074425,18.362404,20.650383,22.938364,24.261955,25.585548,26.913044,28.236637,29.564135,30.274734,30.98924,31.699842,32.41435,33.12495,31.87554,30.626131,29.376722,28.12341,26.874,25.136541,23.399082,21.661623,19.924164,18.186707,17.601046,17.01148,16.42582,15.836256,15.250595,15.160794,15.074897,14.989,14.899199,14.813302,14.723501,14.637604,14.551707,14.461906,14.376009,14.051944,13.723974,13.399908,13.075843,12.751778,13.274967,13.798158,14.325252,14.848442,15.375536,15.988527,16.601519,17.210606,17.823597,18.436588,17.210606,15.988527,14.762545,13.536563,12.31058,11.412568,10.510651,9.612638,8.710721,7.812709,7.5394006,7.262188,6.98888,6.7116675,6.4383593,6.5984397,6.7624245,6.9264097,7.08649,7.250475,6.9264097,6.5984397,6.2743745,5.950309,5.6262436,6.3017054,6.9732623,7.648724,8.324185,8.999647,10.186585,11.373524,12.564366,13.751305,14.938243,16.050997,17.163752,18.276506,19.389261,20.498112,20.861221,21.22433,21.58744,21.95055,22.31366,23.1492,23.988647,24.82419,25.663635,26.499178,24.051117,21.599154,19.151093,16.69913,14.251068,14.949956,15.648844,16.351637,17.050524,17.749413,16.988054,16.226696,15.461433,14.700074,13.938716,17.651802,21.360985,25.074072,28.787157,32.500244,34.413403,36.326557,38.235813,40.148968,42.062126,40.91423,39.762432,38.610634,37.462738,36.31094,35.498825,34.68671,33.874596,33.062477,32.250362,29.247877,26.249296,23.250715,20.24823,17.24965,15.14908,13.048512,10.951848,8.85128,6.7507114,5.7980375,4.8492675,3.900498,2.951728,1.999054,1.6008049,1.1986516,0.80040246,0.39824903,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.23816854,0.3513962,0.46071947,0.57394713,0.6871748,6.3134184,11.935758,17.562002,23.188246,28.810585,30.489477,32.16056,33.839455,35.514442,37.18943,32.898495,28.61146,24.324427,20.037392,15.750359,15.676175,15.598087,15.523903,15.449719,15.375536,15.324779,15.274021,15.223265,15.176412,15.125654,14.364296,13.599033,12.837675,12.076316,11.311053,10.151445,8.987934,7.824422,6.66091,5.5013027,5.0640097,4.6267166,4.1894236,3.7482262,3.310933,2.912684,2.514435,2.1122816,1.7140326,1.3118792,2.174752,3.0376248,3.900498,4.7633705,5.6262436,4.6267166,3.6232853,2.6237583,1.6242313,0.62470436,0.62470436,0.62470436,0.62470436,0.62470436,0.62470436,0.8238289,1.0268579,1.2259823,1.4251068,1.6242313,1.7608855,1.901444,2.0380979,2.174752,2.3114061,2.5378613,2.7643168,2.9868677,3.213323,3.435874,3.1391394,2.8385005,2.5378613,2.2372224,1.9365835,1.6359446,1.33921,1.038571,0.737932,0.43729305,0.5388075,0.63641757,0.737932,0.8394465,0.93705654,0.77307165,0.61299115,0.44900626,0.28892577,0.12494087,0.78868926,1.4485333,2.1122816,2.77603,3.435874,2.87364,2.3114061,1.7491722,1.1869383,0.62470436,0.8394465,1.0502841,1.261122,1.475864,1.6867018,1.3860629,1.0893283,0.78868926,0.48805028,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.113227665,0.22645533,0.3357786,0.44900626,0.5622339,0.60127795,0.63641757,0.6754616,0.7106012,0.74964523,0.8745861,0.999527,1.1244678,1.2494087,1.3743496,1.3509232,1.3235924,1.3001659,1.2767396,1.2494087,1.1869383,1.1244678,1.0619974,0.999527,0.93705654,0.8511597,0.76135844,0.6754616,0.58566034,0.4997635,0.42557985,0.3513962,0.27330816,0.19912452,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.58566034,0.48024148,0.3709182,0.26549935,0.15617609,0.05075723,0.07027924,0.08980125,0.10932326,0.12884527,0.14836729,0.19131571,0.23035973,0.26940376,0.30844778,0.3513962,0.6715572,0.9917182,1.3118792,1.6281357,1.9482968,2.6432803,3.3343596,4.029343,4.7204223,5.4115014,5.368553,5.3256044,5.2865605,5.2436123,5.2006636,5.270943,5.3451266,5.4193106,5.4895897,5.563773,5.3295093,5.099149,4.8648853,4.630621,4.4002614,3.814601,3.2289407,2.6432803,2.0615244,1.475864,1.8389735,2.2059872,2.5690966,2.9361105,3.2992198,3.4007344,3.4983444,3.5998588,3.7013733,3.7989833,3.8809757,3.959064,4.041056,4.1191444,4.2011366,4.154284,4.1113358,4.0644827,4.0215344,3.9746814,3.998108,4.0215344,4.041056,4.0644827,4.087909,4.357313,4.6267166,4.8961205,5.165524,5.4388323,5.618435,5.801942,5.985449,6.168956,6.348558,6.4305506,6.5164475,6.5984397,6.6804323,6.7624245,6.6960497,6.6257706,6.559396,6.493021,6.426646,6.5554914,6.6843367,6.813182,6.9459314,7.0747766,7.320754,7.570636,7.816613,8.066495,8.312472,8.546737,8.781001,9.019169,9.253433,9.487698,9.425227,9.362757,9.300286,9.237816,9.175345,9.019169,8.859089,8.702912,8.546737,8.386656,8.648251,8.905942,9.167537,9.4291315,9.686822,8.343708,6.996689,5.6535745,4.3065557,2.9634414,2.5573835,2.1513257,1.7491722,1.3431144,0.93705654,0.92924774,0.91753453,0.9058213,0.8980125,0.8862993,0.9956226,1.1088502,1.2181735,1.3274968,1.43682,1.2689307,1.1010414,0.93315214,0.76916724,0.60127795,0.4997635,0.39824903,0.30063897,0.19912452,0.10151446,0.19131571,0.28111696,0.3709182,0.46071947,0.5505207,0.5192855,0.48805028,0.46071947,0.42948425,0.39824903,0.32016098,0.23816854,0.16008049,0.078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.30063897,0.60127795,0.9019169,1.1986516,1.4992905,1.5305257,1.5617609,1.5890918,1.620327,1.6515622,1.8116426,1.9717231,2.1318035,2.2918842,2.4480603,2.366068,2.280171,2.194274,2.1083772,2.0263848,2.3348327,2.6432803,2.9556324,3.2640803,3.5764325,4.3729305,5.169429,5.9659266,6.7663293,7.562827,7.8556576,8.148487,8.441318,8.734148,9.023073,8.777096,8.531119,8.281238,8.03526,7.7892823,6.930314,6.0713453,5.2162814,4.357313,3.4983444,3.4983444,3.4983444,3.4983444,3.4983444,3.4983444,3.6349986,3.7716527,3.9044023,4.041056,4.173806,4.21285,4.251894,4.2870336,4.3260775,4.3612175,4.9234514,5.4856853,6.0518236,6.6140575,7.1762915,7.473026,7.7697606,8.066495,8.36323,8.663869,9.089449,9.511124,9.936704,10.362284,10.787864,11.892809,12.997755,14.102701,15.207646,16.312593,18.90902,21.501543,24.097971,26.694399,29.28692,30.739359,32.187893,33.636425,35.088863,36.537395,36.52178,36.50616,36.49445,36.47883,36.46321,34.585194,32.707176,30.82916,28.951143,27.073126,25.491842,23.906654,22.321468,20.73628,19.151093,18.538101,17.92511,17.31212,16.69913,16.086138,15.844065,15.598087,15.35211,15.1061325,14.864059,14.700074,14.53609,14.376009,14.212025,14.048039,13.770826,13.493614,13.216402,12.939189,12.661977,12.943093,13.228115,13.509232,13.794253,14.07537,14.551707,15.024139,15.500477,15.976814,16.449247,15.543426,14.633699,13.727879,12.818152,11.912332,11.158782,10.401327,9.647778,8.894228,8.136774,7.8517528,7.5667315,7.28171,6.996689,6.7116675,6.8209906,6.9264097,7.0357327,7.141152,7.250475,6.9615493,6.6687193,6.379793,6.0908675,5.801942,6.3915067,6.984976,7.578445,8.171914,8.761478,9.796145,10.826907,11.861574,12.892336,13.923099,14.989,16.054901,17.120804,18.186707,19.248703,19.744562,20.240421,20.73628,21.228235,21.724094,22.594776,23.465458,24.33614,25.206821,26.073599,24.20339,22.333181,20.466877,18.596668,16.72646,16.91387,17.101282,17.288692,17.476105,17.663515,17.058334,16.457056,15.855778,15.250595,14.649317,17.589333,20.529346,23.469362,26.409376,29.349392,30.805735,32.26598,33.72232,35.178665,36.638912,36.14305,35.647194,35.151333,34.655476,34.16352,33.28503,32.40654,31.528048,30.653461,29.774971,27.11217,24.449368,21.786564,19.123762,16.46096,14.805493,13.153932,11.498465,9.8429985,8.187531,7.195813,6.2040954,5.2084727,4.2167544,3.2250361,2.854118,2.4792955,2.1083772,1.7335546,1.3626363,2.069333,2.77603,3.4866312,4.193328,4.900025,4.322173,3.7443218,3.1664703,2.5886188,2.0107672,6.2470436,10.48332,14.7156925,18.95197,23.188246,24.55088,25.913517,27.276154,28.63879,30.001427,26.717825,23.438128,20.158428,16.87873,13.599033,14.352583,15.1061325,15.855778,16.609327,17.362877,16.511717,15.664462,14.813302,13.962143,13.110983,12.306676,11.502369,10.698062,9.893755,9.085544,8.152391,7.2192397,6.282183,5.349031,4.4119744,4.0605783,3.7091823,3.3538816,3.0024853,2.6510892,2.330928,2.0146716,1.698415,1.3782539,1.0619974,1.815547,2.5690966,3.3187418,4.0722914,4.825841,3.9629683,3.1000953,2.2372224,1.3743496,0.5114767,0.5544251,0.59737355,0.64032197,0.6832704,0.7262188,1.1361811,1.5461433,1.9561055,2.366068,2.77603,2.7643168,2.7486992,2.736986,2.7252727,2.7135596,2.7565079,2.795552,2.8385005,2.8814487,2.9243972,2.6588979,2.3933985,2.1318035,1.8663043,1.6008049,1.3509232,1.1010414,0.8511597,0.60127795,0.3513962,0.44119745,0.5309987,0.62079996,0.7106012,0.80040246,0.6637484,0.5231899,0.38653582,0.24988174,0.113227665,0.64032197,1.1674163,1.6945106,2.2216048,2.7486992,2.338737,1.9248703,1.5110037,1.1010414,0.6871748,0.8238289,0.95657855,1.0932326,1.2259823,1.3626363,1.1244678,0.8862993,0.6481308,0.41386664,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.12884527,0.26159495,0.39044023,0.5192855,0.6481308,0.6442264,0.64032197,0.63641757,0.62860876,0.62470436,0.7223144,0.8199245,0.91753453,1.0151446,1.1127546,1.1010414,1.0932326,1.0815194,1.0737107,1.0619974,1.0112402,0.96438736,0.9136301,0.8628729,0.81211567,0.7418364,0.6715572,0.60127795,0.5309987,0.46071947,0.39434463,0.3240654,0.25378615,0.1835069,0.113227665,0.113227665,0.11713207,0.12103647,0.12103647,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12103647,0.12103647,0.11713207,0.113227665,0.113227665,0.21083772,0.31235218,0.41386664,0.5114767,0.61299115,0.49195468,0.3670138,0.24597734,0.12103647,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.12103647,0.093705654,0.06637484,0.039044023,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.13274968,0.12884527,0.12103647,0.11713207,0.113227665,0.09761006,0.08199245,0.06637484,0.05075723,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.48805028,0.39824903,0.30844778,0.21864653,0.12884527,0.039044023,0.05075723,0.06637484,0.08199245,0.09761006,0.113227665,0.14055848,0.1717937,0.20302892,0.23426414,0.26159495,0.5036679,0.7418364,0.98390937,1.2220778,1.4641509,1.9834363,2.5066261,3.0298162,3.5530062,4.0761957,4.0527697,4.029343,4.0059166,3.9863946,3.9629683,4.0215344,4.0761957,4.134762,4.193328,4.251894,4.084005,3.9200199,3.7560349,3.5881457,3.4241607,2.9673457,2.5105307,2.0537157,1.5969005,1.1361811,1.4055848,1.6710842,1.9404879,2.2059872,2.475391,2.5495746,2.6237583,2.7018464,2.77603,2.8502135,2.9361105,3.018103,3.1039999,3.1898966,3.2757936,3.2836022,3.2953155,3.3031244,3.3148375,3.3265507,3.4436827,3.5647192,3.6857557,3.8067923,3.9239242,4.0527697,4.181615,4.3065557,4.435401,4.564246,4.7399445,4.9156423,5.095245,5.270943,5.4505453,5.688714,5.930787,6.168956,6.4110284,6.649197,6.6140575,6.578918,6.5437784,6.5086384,6.473499,6.6335793,6.79366,6.9537406,7.113821,7.2739015,7.5823493,7.890797,8.1992445,8.503788,8.812236,9.081639,9.351044,9.6243515,9.893755,10.163159,9.964035,9.761005,9.561881,9.362757,9.163632,9.097258,9.030883,8.968412,8.902037,8.835662,8.944985,9.054309,9.159728,9.269051,9.37447,8.011833,6.6452928,5.278752,3.9161155,2.5495746,2.2020829,1.8545911,1.5070993,1.1596074,0.81211567,0.8160201,0.8238289,0.8277333,0.8316377,0.8394465,0.92143893,1.0034313,1.0854238,1.1674163,1.2494087,1.0893283,0.92924774,0.76916724,0.60908675,0.44900626,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.14055848,0.21083772,0.27721256,0.3435874,0.41386664,0.39044023,0.3670138,0.3435874,0.3240654,0.30063897,0.23816854,0.1796025,0.12103647,0.058566034,0.0,0.0,0.0,0.0,0.0,0.0,0.23816854,0.47633708,0.7106012,0.94876975,1.1869383,1.3235924,1.456342,1.5929961,1.7257458,1.8623998,1.9092526,1.9522011,1.999054,2.0420024,2.0888553,2.0537157,2.0224805,1.9912452,1.9561055,1.9248703,2.1435168,2.366068,2.5847144,2.803361,3.0259118,3.6584249,4.290938,4.9234514,5.5559645,6.1884775,6.559396,6.9342184,7.3051367,7.676055,8.050878,8.054782,8.058686,8.066495,8.070399,8.074304,7.3597984,6.6452928,5.930787,5.2162814,4.5017757,4.388548,4.2753205,4.1620927,4.0488653,3.9356375,4.181615,4.4275923,4.6735697,4.9156423,5.1616197,5.4115014,5.661383,5.911265,6.1611466,6.4110284,6.824895,7.238762,7.648724,8.062591,8.476458,9.007456,9.538455,10.073358,10.604357,11.139259,12.111456,13.087557,14.063657,15.035853,16.011953,17.034906,18.057861,19.080814,20.103767,21.12672,24.02769,26.928663,29.833538,32.73451,35.63548,37.212856,38.78633,40.363712,41.937183,43.51066,42.76882,42.026985,41.28515,40.543312,39.801476,37.29485,34.788223,32.285503,29.778875,27.276154,25.843239,24.410322,22.977407,21.54449,20.111576,19.475159,18.838741,18.19842,17.562002,16.925583,16.52343,16.121277,15.719124,15.313066,14.9109125,14.676648,14.438479,14.200311,13.962143,13.723974,13.493614,13.263254,13.036799,12.806439,12.576079,12.615124,12.654168,12.693212,12.73616,12.775204,13.110983,13.450665,13.786445,14.126127,14.461906,13.872341,13.282777,12.693212,12.103647,11.514082,10.901091,10.292005,9.682918,9.073831,8.460839,8.16801,7.871275,7.578445,7.28171,6.98888,7.039637,7.094299,7.1450562,7.195813,7.250475,6.996689,6.7389984,6.4852123,6.2314262,5.9737353,6.4852123,6.996689,7.504261,8.015738,8.52331,9.4018,10.280292,11.158782,12.033368,12.911859,13.930907,14.946052,15.965101,16.98415,17.999294,18.627903,19.256512,19.881216,20.509825,21.138433,22.04035,22.942268,23.844185,24.746101,25.651922,24.359566,23.071114,21.778755,20.490303,19.20185,18.87388,18.549814,18.22575,17.901684,17.573715,17.132517,16.69132,16.246218,15.80502,15.363823,17.530766,19.69771,21.864653,24.031595,26.19854,27.201971,28.205402,29.208834,30.20836,31.211792,31.371872,31.531952,31.692034,31.852114,32.012196,31.071234,30.126368,29.185408,28.244446,27.29958,24.976461,22.649437,20.326319,17.999294,15.676175,14.465811,13.2554455,12.045081,10.834716,9.6243515,8.589685,7.5550184,6.520352,5.4856853,4.4510183,4.1035266,3.7599394,3.416352,3.06886,2.7252727,4.11524,5.505207,6.8951745,8.285142,9.675109,8.406178,7.141152,5.872221,4.60329,3.338264,6.184573,9.026978,11.873287,14.719597,17.562002,18.612286,19.662569,20.712854,21.763138,22.813423,20.54106,18.268698,15.996336,13.723974,11.4516115,13.028991,14.610273,16.191557,17.768934,19.350218,17.698656,16.050997,14.399435,12.751778,11.100216,10.25296,9.405705,8.55845,7.7111945,6.8639393,6.153338,5.446641,4.7399445,4.0332475,3.3265507,3.057147,2.7916477,2.522244,2.2567444,1.9873407,1.7530766,1.5188124,1.2806439,1.0463798,0.81211567,1.456342,2.096664,2.7408905,3.3812122,4.025439,3.2992198,2.5769055,1.8506867,1.1244678,0.39824903,0.48414588,0.5700427,0.6559396,0.7418364,0.8238289,1.4446288,2.0654287,2.6862288,3.3031244,3.9239242,3.7638438,3.5998588,3.435874,3.2757936,3.1118085,2.97125,2.8306916,2.6940374,2.5534792,2.4129205,2.182561,1.9522011,1.7218413,1.4914817,1.261122,1.0619974,0.8628729,0.6637484,0.46071947,0.26159495,0.3435874,0.42167544,0.5036679,0.58175594,0.6637484,0.5505207,0.43729305,0.3240654,0.21083772,0.10151446,0.49195468,0.8862993,1.2767396,1.6710842,2.0615244,1.7999294,1.5383345,1.2767396,1.0112402,0.74964523,0.80821127,0.8667773,0.92143893,0.98000497,1.038571,0.8628729,0.6871748,0.5114767,0.3357786,0.1639849,0.12884527,0.09761006,0.06637484,0.031235218,0.0,0.14836729,0.29673457,0.44119745,0.58956474,0.737932,0.6910792,0.6442264,0.59346914,0.5466163,0.4997635,0.5700427,0.64032197,0.7106012,0.78088045,0.8511597,0.8550641,0.8589685,0.8667773,0.8706817,0.8745861,0.8394465,0.80040246,0.76135844,0.7262188,0.6871748,0.63641757,0.58175594,0.5309987,0.47633708,0.42557985,0.359205,0.29673457,0.23035973,0.1639849,0.10151446,0.10541886,0.10932326,0.113227665,0.12103647,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12103647,0.113227665,0.10932326,0.10541886,0.10151446,0.31235218,0.5231899,0.737932,0.94876975,1.1635119,0.92924774,0.698888,0.46462387,0.23426414,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.093705654,0.078088045,0.058566034,0.042948425,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05466163,0.10932326,0.1639849,0.21864653,0.27330816,0.26549935,0.25378615,0.24597734,0.23426414,0.22645533,0.19522011,0.1639849,0.13665408,0.10541886,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.38653582,0.31625658,0.24207294,0.1717937,0.09761006,0.023426414,0.03513962,0.046852827,0.05466163,0.06637484,0.07418364,0.093705654,0.113227665,0.13665408,0.15617609,0.1756981,0.3357786,0.4958591,0.6559396,0.8160201,0.97610056,1.3274968,1.678893,2.0341935,2.3855898,2.736986,2.7330816,2.7330816,2.7291772,2.7291772,2.7252727,2.7682211,2.8111696,2.854118,2.893162,2.9361105,2.8385005,2.7408905,2.6432803,2.5456703,2.4480603,2.1200905,1.7882162,1.4602464,1.1283722,0.80040246,0.96829176,1.1400855,1.3118792,1.4797685,1.6515622,1.698415,1.7491722,1.7999294,1.8506867,1.901444,1.9912452,2.0810463,2.1708477,2.260649,2.35045,2.416825,2.4792955,2.5456703,2.6081407,2.6745155,2.893162,3.1118085,3.3265507,3.5451972,3.7638438,3.7482262,3.7326086,3.716991,3.7013733,3.6857557,3.8614538,4.0332475,4.2050414,4.376835,4.548629,4.9468775,5.3451266,5.743376,6.141625,6.5359693,6.5359693,6.532065,6.5281606,6.5281606,6.524256,6.715572,6.9068875,7.094299,7.2856145,7.47693,7.843944,8.210958,8.577971,8.944985,9.311999,9.616543,9.921086,10.22563,10.534078,10.838621,10.498938,10.163159,9.823476,9.487698,9.151918,9.17925,9.20658,9.2339115,9.261242,9.288573,9.24172,9.198771,9.151918,9.108971,9.062118,7.676055,6.2938967,4.9078336,3.521771,2.135708,1.8467822,1.5578566,1.2689307,0.97610056,0.6871748,0.7066968,0.7262188,0.74574083,0.76916724,0.78868926,0.8433509,0.8980125,0.95267415,1.0073358,1.0619974,0.9097257,0.75745404,0.60518235,0.45291066,0.30063897,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.093705654,0.14055848,0.1835069,0.23035973,0.27330816,0.26159495,0.24597734,0.23035973,0.21474212,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.1756981,0.3513962,0.5231899,0.698888,0.8745861,1.116659,1.3548276,1.5969005,1.8350691,2.0732377,2.0068626,1.9365835,1.8663043,1.796025,1.7257458,1.7452679,1.7647898,1.7843118,1.8038338,1.8233559,1.9561055,2.084951,2.2137961,2.3465457,2.475391,2.9439192,3.408543,3.8770714,4.3455997,4.814128,5.263134,5.716045,6.168956,6.621866,7.0747766,7.3324676,7.590158,7.8478484,8.105539,8.36323,7.7892823,7.2192397,6.6452928,6.0713453,5.5013027,5.2748475,5.0483923,4.825841,4.5993857,4.376835,4.728231,5.083532,5.4388323,5.794133,6.1494336,6.6140575,7.0747766,7.5394006,8.00012,8.460839,8.726339,8.987934,9.249529,9.511124,9.776623,10.541886,11.311053,12.076316,12.845484,13.610746,15.137367,16.663988,18.186707,19.713327,21.236044,22.177006,23.117966,24.058928,24.995983,25.936945,29.146362,32.35578,35.569103,38.778522,41.98794,43.686356,45.388676,47.08709,48.78941,50.487827,49.015865,47.54781,46.07585,44.607796,43.135838,40.004505,36.873177,33.741844,30.60661,27.475279,26.194635,24.91399,23.633347,22.356607,21.075964,20.412214,19.748466,19.088623,18.424873,17.761126,17.202797,16.644466,16.082233,15.523903,14.96167,14.649317,14.336966,14.024612,13.712261,13.399908,13.216402,13.036799,12.853292,12.6697855,12.486279,12.28325,12.084125,11.881096,11.678067,11.475039,11.674163,11.873287,12.076316,12.27544,12.4745655,12.201257,11.931853,11.6585455,11.385237,11.111929,10.647305,10.182681,9.718058,9.253433,8.78881,8.484266,8.175818,7.871275,7.5667315,7.262188,7.2582836,7.2582836,7.2543793,7.2543793,7.250475,7.0318284,6.8092775,6.590631,6.36808,6.1494336,6.578918,7.0044975,7.433982,7.859562,8.289046,9.01136,9.733675,10.455989,11.178304,11.900618,12.86891,13.841106,14.809398,15.781594,16.749886,17.511244,18.268698,19.030056,19.791414,20.548868,21.485926,22.419077,23.356134,24.289286,25.226343,24.515741,23.805141,23.09454,22.383938,21.673336,20.837795,19.998348,19.162806,18.32336,17.487818,17.206701,16.921679,16.640562,16.359446,16.074425,17.468296,18.866072,20.259943,21.653814,23.05159,23.598207,24.144823,24.69144,25.238056,25.788576,26.600693,27.416712,28.232733,29.048752,29.860868,28.853533,27.846197,26.838861,25.831526,24.82419,22.83685,20.849508,18.862167,16.874826,14.8874855,14.122223,13.35696,12.591698,11.826434,11.061172,9.983557,8.905942,7.8283267,6.7507114,5.6730967,5.35684,5.040583,4.7243266,4.4041657,4.087909,6.1611466,8.234385,10.303718,12.376955,14.450192,12.494087,10.534078,8.577971,6.621866,4.661856,6.1181984,7.570636,9.026978,10.48332,11.935758,12.67369,13.411622,14.149553,14.8874855,15.625418,14.360392,13.095366,11.8303385,10.565312,9.300286,11.709302,14.114414,16.52343,18.928543,21.337559,18.885593,16.437534,13.985569,11.537509,9.085544,8.1992445,7.309041,6.4188375,5.5286336,4.6384296,4.1581883,3.677947,3.1977055,2.717464,2.2372224,2.0537157,1.8741131,1.6906061,1.5070993,1.3235924,1.1713207,1.0190489,0.8667773,0.7145056,0.5622339,1.0932326,1.6281357,2.1591344,2.6940374,3.2250361,2.639376,2.0498111,1.4641509,0.8745861,0.28892577,0.41386664,0.5427119,0.6715572,0.79649806,0.92534333,1.756981,2.5847144,3.416352,4.2440853,5.0757227,4.7633705,4.4510183,4.138666,3.8263142,3.513962,3.1898966,2.8658314,2.5456703,2.2216048,1.901444,1.7062237,1.5110037,1.3157835,1.1205635,0.92534333,0.77307165,0.62470436,0.47633708,0.3240654,0.1756981,0.24597734,0.31625658,0.38653582,0.45681506,0.5231899,0.43729305,0.3513962,0.26159495,0.1756981,0.08589685,0.3435874,0.60127795,0.8589685,1.116659,1.3743496,1.261122,1.1517987,1.038571,0.92534333,0.81211567,0.79259366,0.77307165,0.75354964,0.7340276,0.7106012,0.60127795,0.48805028,0.37482262,0.26159495,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.1639849,0.3318742,0.4958591,0.659844,0.8238289,0.7340276,0.6442264,0.5544251,0.46462387,0.37482262,0.41777104,0.46071947,0.5036679,0.5466163,0.58566034,0.60908675,0.62860876,0.6481308,0.6676528,0.6871748,0.6637484,0.63641757,0.61299115,0.58566034,0.5622339,0.5270943,0.49195468,0.45681506,0.42167544,0.38653582,0.3279698,0.26940376,0.20693332,0.14836729,0.08589685,0.093705654,0.10151446,0.10932326,0.11713207,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.11713207,0.10932326,0.10151446,0.093705654,0.08589685,0.41386664,0.737932,1.0619974,1.3860629,1.7140326,1.3704453,1.0268579,0.6832704,0.3435874,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.06637484,0.058566034,0.05075723,0.046852827,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08199245,0.1639849,0.24597734,0.3318742,0.41386664,0.39824903,0.38263142,0.3670138,0.3513962,0.3357786,0.29283017,0.24597734,0.20302892,0.15617609,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28892577,0.23426414,0.1756981,0.12103647,0.06637484,0.011713207,0.015617609,0.023426414,0.027330816,0.031235218,0.039044023,0.046852827,0.058566034,0.06637484,0.078088045,0.08589685,0.1678893,0.24597734,0.3279698,0.40605783,0.48805028,0.6715572,0.8511597,1.0346665,1.2181735,1.4016805,1.4172981,1.43682,1.4524376,1.4680552,1.4875772,1.5149081,1.542239,1.5695697,1.5969005,1.6242313,1.5969005,1.5656652,1.53443,1.5031948,1.475864,1.2728351,1.0698062,0.8667773,0.6637484,0.46071947,0.5349031,0.60908675,0.679366,0.75354964,0.8238289,0.8511597,0.8745861,0.9019169,0.92534333,0.94876975,1.0463798,1.1400855,1.2337911,1.3314011,1.4251068,1.5461433,1.6632754,1.7843118,1.9053483,2.0263848,2.338737,2.6549935,2.97125,3.2836022,3.5998588,3.4436827,3.2836022,3.1274261,2.97125,2.8111696,2.979059,3.1469483,3.3148375,3.4827268,3.6506162,4.2050414,4.759466,5.3138914,5.8683167,6.426646,6.453977,6.4852123,6.5164475,6.5437784,6.575013,6.79366,7.016211,7.2348576,7.453504,7.676055,8.101635,8.531119,8.956698,9.386183,9.811763,10.151445,10.491129,10.8308115,11.174399,11.514082,11.037745,10.561408,10.088976,9.612638,9.136301,9.257338,9.378374,9.499411,9.616543,9.737579,9.538455,9.343235,9.14411,8.94889,8.749765,7.3441806,5.938596,4.533011,3.1313305,1.7257458,1.4914817,1.261122,1.0268579,0.79649806,0.5622339,0.59737355,0.63251317,0.6676528,0.7027924,0.737932,0.76526284,0.79259366,0.8199245,0.8472553,0.8745861,0.7301232,0.58566034,0.44119745,0.29673457,0.14836729,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.046852827,0.07027924,0.093705654,0.113227665,0.13665408,0.12884527,0.12103647,0.113227665,0.10932326,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.113227665,0.22645533,0.3357786,0.44900626,0.5622339,0.9058213,1.2533131,1.5969005,1.9443923,2.2879796,2.1005683,1.9170616,1.7335546,1.5461433,1.3626363,1.43682,1.5070993,1.5812829,1.6515622,1.7257458,1.7647898,1.8038338,1.8467822,1.8858263,1.9248703,2.2294137,2.5300527,2.8306916,3.135235,3.435874,3.970777,4.5017757,5.036679,5.5676775,6.098676,6.610153,7.1216297,7.629202,8.140678,8.648251,8.218767,7.7892823,7.3597984,6.930314,6.5008297,6.1611466,5.825368,5.4856853,5.1499066,4.814128,5.278752,5.743376,6.2079997,6.6726236,7.137247,7.812709,8.488171,9.163632,9.839094,10.510651,10.6238785,10.737106,10.850334,10.963562,11.076789,12.076316,13.079747,14.0831785,15.086611,16.086138,18.163279,20.236517,22.31366,24.386896,26.464039,27.319103,28.178072,29.037039,29.892103,30.751072,34.26894,37.786804,41.300766,44.818634,48.3365,50.16376,51.987118,53.814377,55.637733,57.461086,55.266815,53.068634,50.870457,48.67228,46.4741,42.71416,38.95422,35.194283,31.434343,27.674404,26.54603,25.421562,24.29319,23.164818,22.036446,21.349272,20.662096,19.974922,19.287746,18.600573,17.882162,17.163752,16.449247,15.730837,15.012426,14.625891,14.239355,13.848915,13.462379,13.075843,12.939189,12.806439,12.6697855,12.533132,12.400381,11.955279,11.510178,11.065076,10.619974,10.174872,10.237343,10.299813,10.362284,10.424754,10.487225,10.534078,10.577025,10.6238785,10.666827,10.71368,10.393518,10.073358,9.753197,9.433036,9.112875,8.796618,8.484266,8.16801,7.8517528,7.5394006,7.480835,7.422269,7.363703,7.309041,7.250475,7.0630636,6.8795567,6.6960497,6.5086384,6.3251314,6.6687193,7.016211,7.3597984,7.703386,8.050878,8.617016,9.183154,9.753197,10.319335,10.889378,11.810817,12.732256,13.653695,14.579038,15.500477,16.39068,17.284788,18.178898,19.069101,19.96321,20.931501,21.895887,22.86418,23.832472,24.800762,24.671917,24.539167,24.410322,24.281477,24.148727,22.801708,21.450787,20.099863,18.74894,17.40192,17.27698,17.155943,17.031002,16.909966,16.788929,17.409729,18.030529,18.655233,19.276033,19.900738,19.99054,20.084246,20.177952,20.271656,20.361458,21.833418,23.301472,24.773432,26.241488,27.713448,26.639736,25.566027,24.49622,23.422508,22.348799,20.701141,19.049578,17.398016,15.750359,14.098797,13.778636,13.458474,13.138313,12.818152,12.501896,11.381332,10.260769,9.140205,8.019642,6.899079,6.610153,6.321227,6.028397,5.7394714,5.4505453,8.207053,10.959657,13.716166,16.46877,19.225277,16.578093,13.930907,11.283723,8.636538,5.989353,6.0518236,6.1181984,6.180669,6.2470436,6.3134184,6.7389984,7.1606736,7.5862536,8.011833,8.437413,8.179723,7.9220324,7.6643414,7.406651,7.1489606,10.38571,13.618555,16.855305,20.08815,23.3249,20.076437,16.82407,13.575606,10.323239,7.0747766,6.141625,5.2084727,4.279225,3.3460727,2.4129205,2.1591344,1.9092526,1.6554666,1.4016805,1.1517987,1.0541886,0.95657855,0.8589685,0.76135844,0.6637484,0.59346914,0.5231899,0.45291066,0.38263142,0.31235218,0.7340276,1.1557031,1.5812829,2.0029583,2.4246337,1.9756275,1.5266213,1.0737107,0.62470436,0.1756981,0.3435874,0.5153811,0.6832704,0.8550641,1.0268579,2.0654287,3.1039999,4.1464753,5.185046,6.223617,5.7628975,5.298274,4.8375545,4.376835,3.912211,3.408543,2.900971,2.397303,1.893635,1.3860629,1.2259823,1.0659018,0.9058213,0.74574083,0.58566034,0.48805028,0.38653582,0.28892577,0.18741131,0.08589685,0.14836729,0.20693332,0.26940376,0.3279698,0.38653582,0.3240654,0.26159495,0.19912452,0.13665408,0.07418364,0.19912452,0.32016098,0.44119745,0.5661383,0.6871748,0.7262188,0.76135844,0.80040246,0.8394465,0.8745861,0.77697605,0.679366,0.58175594,0.48414588,0.38653582,0.3357786,0.28892577,0.23816854,0.18741131,0.13665408,0.10932326,0.08199245,0.05466163,0.027330816,0.0,0.1835069,0.3631094,0.5466163,0.7301232,0.9136301,0.78088045,0.6481308,0.5153811,0.38263142,0.24988174,0.26549935,0.28111696,0.29673457,0.30844778,0.3240654,0.359205,0.39434463,0.42948425,0.46462387,0.4997635,0.48805028,0.47633708,0.46071947,0.44900626,0.43729305,0.42167544,0.40215343,0.38653582,0.3670138,0.3513962,0.29673457,0.23816854,0.1835069,0.12884527,0.07418364,0.08589685,0.093705654,0.10541886,0.113227665,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.113227665,0.10541886,0.093705654,0.08589685,0.07418364,0.5114767,0.94876975,1.3860629,1.8233559,2.260649,1.8116426,1.358732,0.9058213,0.45291066,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.039044023,0.042948425,0.046852827,0.046852827,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10932326,0.21864653,0.3318742,0.44119745,0.5505207,0.5309987,0.5114767,0.48805028,0.46852827,0.44900626,0.39044023,0.3318742,0.26940376,0.21083772,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.10151446,0.13665408,0.1756981,0.21083772,0.24988174,0.26159495,0.27330816,0.28892577,0.30063897,0.31235218,0.3513962,0.38653582,0.42557985,0.46071947,0.4997635,0.42557985,0.3513962,0.27330816,0.19912452,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.6754616,0.8511597,1.0268579,1.1986516,1.3743496,1.7882162,2.1981785,2.612045,3.0259118,3.435874,3.1391394,2.8385005,2.5378613,2.2372224,1.9365835,2.1005683,2.260649,2.4246337,2.5886188,2.7486992,3.4632049,4.173806,4.8883114,5.5989127,6.3134184,6.375889,6.4383593,6.5008297,6.5633,6.6257706,6.8756523,7.125534,7.375416,7.6252975,7.8751793,8.36323,8.85128,9.339331,9.823476,10.311526,10.686349,11.061172,11.435994,11.810817,12.185639,11.576552,10.963562,10.350571,9.737579,9.124588,9.339331,9.550168,9.761005,9.975748,10.186585,9.839094,9.487698,9.136301,8.78881,8.437413,7.012306,5.5871997,4.1620927,2.736986,1.3118792,1.1361811,0.96438736,0.78868926,0.61299115,0.43729305,0.48805028,0.5388075,0.58566034,0.63641757,0.6871748,0.6871748,0.6871748,0.6871748,0.6871748,0.6871748,0.5505207,0.41386664,0.27330816,0.13665408,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.698888,1.1517987,1.6008049,2.0498111,2.4988174,2.1981785,1.901444,1.6008049,1.3001659,0.999527,1.1244678,1.2494087,1.3743496,1.4992905,1.6242313,1.5734742,1.5266213,1.475864,1.4251068,1.3743496,1.5110037,1.6515622,1.7882162,1.9248703,2.0615244,2.6745155,3.2875066,3.900498,4.513489,5.12648,5.8878384,6.649197,7.4144597,8.175818,8.937177,8.648251,8.36323,8.074304,7.7892823,7.5003567,7.0513506,6.5984397,6.1494336,5.700427,5.251421,5.825368,6.3993154,6.9732623,7.551114,8.125061,9.01136,9.901564,10.787864,11.674163,12.564366,12.525322,12.486279,12.4511385,12.412095,12.373051,13.610746,14.848442,16.086138,17.323833,18.56153,21.189192,23.81295,26.436708,29.064371,31.68813,32.4612,33.23818,34.01125,34.788223,35.561295,39.38761,43.213924,47.036335,50.862648,54.68896,56.63726,58.585556,60.537758,62.486053,64.438255,61.51386,58.58946,55.66116,52.736763,49.812363,45.423817,41.039173,36.650623,32.262077,27.873528,26.90133,25.925232,24.949131,23.976934,23.000834,22.286327,21.575727,20.861221,20.15062,19.436115,18.56153,17.686943,16.812357,15.93777,15.063184,14.59856,14.13784,13.673217,13.212498,12.751778,12.661977,12.576079,12.486279,12.400381,12.31058,11.623405,10.936231,10.249056,9.561881,8.874706,8.800523,8.726339,8.648251,8.574067,8.499884,8.862993,9.226103,9.589212,9.948417,10.311526,10.135828,9.964035,9.788337,9.612638,9.43694,9.112875,8.78881,8.460839,8.136774,7.812709,7.699481,7.5862536,7.47693,7.363703,7.250475,7.098203,6.949836,6.801469,6.649197,6.5008297,6.7624245,7.0240197,7.2856145,7.551114,7.812709,8.226576,8.636538,9.050405,9.464272,9.874233,10.748819,11.623405,12.501896,13.376482,14.251068,15.274021,16.300879,17.323833,18.35069,19.373644,20.37317,21.376602,22.37613,23.375656,24.375183,24.82419,25.273195,25.726107,26.175114,26.624119,24.761719,22.899319,21.036919,19.174519,17.31212,17.351164,17.386303,17.425346,17.464392,17.49953,17.351164,17.198893,17.050524,16.898252,16.749886,16.386776,16.023666,15.660558,15.3013525,14.938243,17.062239,19.186234,21.314133,23.438128,25.562122,24.425941,23.285854,22.149673,21.013493,19.873407,18.56153,17.24965,15.93777,14.625891,13.314012,13.438952,13.563893,13.688834,13.813775,13.938716,12.775204,11.611692,10.44818,9.288573,8.125061,7.8634663,7.601871,7.336372,7.0747766,6.813182,10.249056,13.688834,17.124708,20.564487,24.00036,20.662096,17.323833,13.985569,10.651209,7.3129454,5.989353,4.661856,3.338264,2.0107672,0.6871748,0.80040246,0.9136301,1.0268579,1.1361811,1.2494087,1.999054,2.7486992,3.4983444,4.251894,5.001539,9.062118,13.1266,17.18718,21.251661,25.31224,21.263374,17.21451,13.16174,9.112875,5.0640097,4.087909,3.1118085,2.135708,1.1635119,0.18741131,0.1639849,0.13665408,0.113227665,0.08589685,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.37482262,0.6871748,0.999527,1.3118792,1.6242313,1.3118792,0.999527,0.6871748,0.37482262,0.062470436,0.27330816,0.48805028,0.698888,0.9136301,1.1244678,2.3738766,3.6232853,4.8765984,6.126007,7.375416,6.7624245,6.1494336,5.5364423,4.9234514,4.3143644,3.6232853,2.9361105,2.2489357,1.5617609,0.8745861,0.74964523,0.62470436,0.4997635,0.37482262,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.21083772,0.1756981,0.13665408,0.10151446,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.18741131,0.37482262,0.5622339,0.74964523,0.93705654,0.76135844,0.58566034,0.41386664,0.23816854,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.19912452,0.39824903,0.60127795,0.80040246,0.999527,0.8238289,0.6481308,0.47633708,0.30063897,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.113227665,0.1639849,0.21083772,0.26159495,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.61299115,1.1635119,1.7140326,2.260649,2.8111696,2.2489357,1.6867018,1.1244678,0.5622339,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13665408,0.27330816,0.41386664,0.5505207,0.6871748,0.6637484,0.63641757,0.61299115,0.58566034,0.5622339,0.48805028,0.41386664,0.3357786,0.26159495,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.078088045,0.10932326,0.14055848,0.1717937,0.19912452,0.21083772,0.21864653,0.23035973,0.23816854,0.24988174,0.28111696,0.30844778,0.339683,0.3709182,0.39824903,0.339683,0.28111696,0.21864653,0.16008049,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,0.5583295,0.71841,0.8784905,1.038571,1.1986516,1.5969005,1.9951496,2.3933985,2.7916477,3.1859922,2.9361105,2.6862288,2.436347,2.1864653,1.9365835,2.0927596,2.2489357,2.4012074,2.5573835,2.7135596,3.357786,4.0020123,4.646239,5.2943697,5.938596,6.0713453,6.2079997,6.3407493,6.477403,6.6140575,6.8287997,7.043542,7.2582836,7.473026,7.687768,8.066495,8.449126,8.827853,9.20658,9.589212,9.905469,10.221725,10.541886,10.858143,11.174399,10.709775,10.2451515,9.780528,9.315904,8.85128,9.081639,9.308095,9.538455,9.768814,9.999174,9.60483,9.2104845,8.81614,8.421796,8.023546,6.707763,5.3919797,4.0722914,2.7565079,1.43682,1.261122,1.0815194,0.9058213,0.7262188,0.5505207,0.5661383,0.58566034,0.60127795,0.62079996,0.63641757,0.62079996,0.60127795,0.58566034,0.5661383,0.5505207,0.44119745,0.3318742,0.21864653,0.10932326,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.093705654,0.14055848,0.19131571,0.23816854,0.61689556,0.9956226,1.3782539,1.756981,2.135708,1.9561055,1.7765031,1.5969005,1.4172981,1.2376955,1.3314011,1.4212024,1.5149081,1.6086137,1.698415,1.6671798,1.6359446,1.6008049,1.5695697,1.5383345,1.7218413,1.901444,2.084951,2.2684577,2.4519646,3.049338,3.6506162,4.251894,4.8492675,5.4505453,6.098676,6.7507114,7.3988423,8.050878,8.699008,8.367134,8.03526,7.703386,7.3715115,7.0357327,6.7624245,6.4891167,6.211904,5.938596,5.661383,6.3134184,6.9615493,7.6135845,8.261715,8.913751,9.679013,10.444276,11.205634,11.970898,12.73616,12.96652,13.192975,13.419431,13.645885,13.8762455,15.566852,17.261362,18.95197,20.646479,22.337086,24.289286,26.241488,28.19369,30.14589,32.09809,33.351402,34.604717,35.858032,37.111343,38.360752,42.36667,46.372585,50.3785,54.38442,58.386433,60.151222,61.912106,63.676895,65.43778,67.19867,63.98925,60.775925,57.562603,54.34928,51.135956,46.786453,42.436947,38.087444,33.73794,29.388435,28.291298,27.198067,26.10093,25.007696,23.914463,23.012547,22.11063,21.212618,20.310701,19.412687,18.249176,17.085665,15.926057,14.762545,13.599033,13.087557,12.576079,12.0606985,11.549222,11.037745,11.014318,10.990892,10.971371,10.947944,10.924518,10.370092,9.815667,9.261242,8.706817,8.148487,8.140678,8.136774,8.128965,8.121157,8.113348,8.413987,8.710721,9.01136,9.311999,9.612638,9.413514,9.21439,9.01136,8.812236,8.6131115,8.320281,8.027451,7.734621,7.4417906,7.1489606,7.168483,7.1841,7.2036223,7.2192397,7.238762,7.08649,6.9342184,6.7780423,6.6257706,6.473499,6.5945354,6.715572,6.8366084,6.9537406,7.0747766,7.6409154,8.203149,8.769287,9.335425,9.901564,10.87376,11.845957,12.818152,13.790349,14.762545,15.7035055,16.64837,17.589333,18.534197,19.475159,20.416119,21.360985,22.301945,23.24681,24.187773,24.574308,24.95694,25.343475,25.726107,26.112642,24.507933,22.903223,21.298513,19.693806,18.089096,18.007103,17.929016,17.847023,17.768934,17.686943,17.378494,17.073952,16.765503,16.457056,16.148607,15.781594,15.410676,15.039758,14.668839,14.301826,15.953387,17.608854,19.26432,20.919786,22.575254,22.001307,21.431265,20.857317,20.28337,19.713327,18.475632,17.237936,16.00024,14.762545,13.524849,14.17298,14.821111,15.469242,16.113468,16.761599,15.410676,14.063657,12.712734,11.361811,10.010887,9.999174,9.987461,9.975748,9.964035,9.948417,12.240301,14.528281,16.820166,19.108145,21.400028,18.440493,15.480955,12.521418,9.557977,6.5984397,5.6730967,4.743849,3.8185053,2.8892577,1.9639144,1.796025,1.6320401,1.4680552,1.3040704,1.1361811,2.0107672,2.8892577,3.7638438,4.6384296,5.5130157,8.577971,11.642927,14.707883,17.772839,20.837795,17.905588,14.977287,12.0489855,9.116779,6.1884775,5.138193,4.087909,3.0376248,1.9873407,0.93705654,0.94096094,0.94876975,0.95267415,0.95657855,0.96438736,0.9058213,0.8511597,0.79649806,0.7418364,0.6871748,1.2845483,1.8819219,2.4792955,3.076669,3.6740425,3.513962,3.349977,3.1859922,3.0259118,2.8619268,3.1703746,3.4788225,3.7833657,4.0918136,4.4002614,3.970777,3.5451972,3.1157131,2.690133,2.260649,2.9907722,3.7208953,4.4510183,5.181142,5.911265,5.4193106,4.927356,4.435401,3.9434462,3.4514916,3.0922866,2.7330816,2.377781,2.018576,1.6632754,1.5851873,1.5070993,1.4290112,1.3509232,1.2767396,1.0307622,0.78868926,0.5466163,0.30454338,0.062470436,0.08980125,0.11713207,0.14446288,0.1717937,0.19912452,0.1756981,0.14836729,0.12494087,0.10151446,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.19131571,0.37872702,0.5700427,0.76135844,0.94876975,0.77307165,0.59346914,0.41777104,0.23816854,0.062470436,0.07027924,0.078088045,0.08589685,0.093705654,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.3318742,0.6637484,0.9956226,1.3314011,1.6632754,1.3938715,1.1283722,0.8589685,0.59346914,0.3240654,0.26940376,0.21474212,0.16008049,0.10541886,0.05075723,0.08980125,0.12884527,0.1717937,0.21083772,0.24988174,0.3279698,0.40605783,0.48414588,0.5583295,0.63641757,0.57785153,0.5192855,0.45681506,0.39824903,0.3357786,0.3513962,0.3670138,0.38263142,0.39824903,0.41386664,0.5700427,0.7262188,0.8862993,1.0424755,1.1986516,1.1517987,1.1010414,1.0502841,0.999527,0.94876975,0.9058213,0.8667773,0.8238289,0.78088045,0.737932,1.0463798,1.358732,1.6671798,1.9756275,2.2879796,1.8506867,1.4172981,0.98390937,0.5466163,0.113227665,0.11713207,0.12103647,0.12884527,0.13274968,0.13665408,0.21474212,0.29283017,0.3709182,0.44900626,0.5231899,0.5114767,0.4997635,0.48805028,0.47633708,0.46071947,0.5114767,0.5583295,0.60518235,0.6520352,0.698888,0.6559396,0.61689556,0.57394713,0.5309987,0.48805028,0.5192855,0.5544251,0.58566034,0.61689556,0.6481308,0.61299115,0.57394713,0.5388075,0.4997635,0.46071947,0.46852827,0.47243267,0.47633708,0.48414588,0.48805028,0.40605783,0.3279698,0.24597734,0.1678893,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.093705654,0.16008049,0.22645533,0.29673457,0.3631094,0.30063897,0.24207294,0.1835069,0.12103647,0.062470436,0.12103647,0.1835069,0.24207294,0.30063897,0.3631094,0.30844778,0.25378615,0.19912452,0.14446288,0.08589685,0.12103647,0.15227169,0.1835069,0.21864653,0.24988174,0.22645533,0.20693332,0.1835069,0.16008049,0.13665408,0.10932326,0.08199245,0.05466163,0.027330816,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.058566034,0.08199245,0.10541886,0.12884527,0.14836729,0.15617609,0.1639849,0.1717937,0.1796025,0.18741131,0.21083772,0.23426414,0.25378615,0.27721256,0.30063897,0.25378615,0.21083772,0.1639849,0.12103647,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.44510186,0.58956474,0.7340276,0.8784905,1.0268579,1.4055848,1.7882162,2.1708477,2.5534792,2.9361105,2.736986,2.5378613,2.338737,2.135708,1.9365835,2.084951,2.233318,2.3816853,2.5261483,2.6745155,3.252367,3.8302186,4.40807,4.985922,5.563773,5.7707067,5.9776397,6.184573,6.3915067,6.5984397,6.7819467,6.9615493,7.141152,7.320754,7.5003567,7.773665,8.043069,8.316377,8.589685,8.862993,9.120684,9.382278,9.643873,9.901564,10.163159,9.846903,9.526741,9.2104845,8.894228,8.574067,8.823949,9.069926,9.315904,9.565785,9.811763,9.370565,8.933272,8.492075,8.050878,7.6135845,6.4032197,5.192855,3.9824903,2.7721257,1.5617609,1.3821584,1.2025559,1.0229534,0.8433509,0.6637484,0.6481308,0.63251317,0.61689556,0.60127795,0.58566034,0.5544251,0.5192855,0.48414588,0.44900626,0.41386664,0.3318742,0.24597734,0.1639849,0.08199245,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.046852827,0.08980125,0.13665408,0.1796025,0.22645533,0.5349031,0.8433509,1.1557031,1.4641509,1.7765031,1.7140326,1.6554666,1.5969005,1.53443,1.475864,1.53443,1.5969005,1.6554666,1.7140326,1.7765031,1.7608855,1.7452679,1.7296503,1.7140326,1.698415,1.9287747,2.15523,2.3816853,2.6081407,2.8385005,3.4241607,4.0137253,4.5993857,5.1889505,5.774611,6.3134184,6.8483214,7.387129,7.9259367,8.460839,8.086017,7.70729,7.328563,6.9537406,6.575013,6.473499,6.375889,6.2743745,6.1767645,6.0752497,6.801469,7.523783,8.250002,8.976221,9.698535,10.342762,10.983084,11.62731,12.271536,12.911859,13.403813,13.895767,14.391626,14.883581,15.375536,17.522957,19.670378,21.8178,23.965221,26.112642,27.393286,28.673931,29.95067,31.231314,32.51196,34.241608,35.971256,37.70091,39.430557,41.164112,45.345726,49.531246,53.716766,57.902287,62.087803,63.661278,65.238655,66.81213,68.385605,69.96298,66.46073,62.96239,59.464046,55.961796,52.46345,48.14909,43.838627,39.524265,35.213802,30.899439,29.685171,28.470901,27.256632,26.038458,24.82419,23.738766,22.649437,21.564014,20.474686,19.389261,17.936825,16.48829,15.035853,13.58732,12.138786,11.576552,11.014318,10.44818,9.885946,9.323712,9.366661,9.40961,9.452558,9.495506,9.538455,9.116779,8.691199,8.269524,7.8478484,7.426173,7.4847393,7.5433054,7.605776,7.6643414,7.726812,7.9610763,8.1992445,8.437413,8.675582,8.913751,8.687295,8.460839,8.238289,8.011833,7.7892823,7.5276875,7.266093,7.008402,6.746807,6.4891167,6.6335793,6.7819467,6.930314,7.0786815,7.223144,7.0708723,6.914696,6.75852,6.606249,6.4500723,6.426646,6.4032197,6.3836975,6.3602715,6.336845,7.055255,7.773665,8.488171,9.20658,9.924991,10.994797,12.064603,13.134409,14.204215,15.274021,16.136894,16.995863,17.854832,18.7138,19.576674,20.459068,21.345367,22.231667,23.114061,24.00036,24.320522,24.640682,24.960844,25.281004,25.601166,24.254147,22.903223,21.556206,20.209187,18.862167,18.663042,18.467823,18.268698,18.073479,17.874353,17.409729,16.945107,16.480482,16.015858,15.551234,15.172507,14.79378,14.418958,14.040231,13.661504,14.848442,16.031475,17.218414,18.401447,19.588387,19.580578,19.57277,19.56496,19.557152,19.549341,18.38583,17.226223,16.062712,14.899199,13.735687,14.907008,16.07833,17.245745,18.417065,19.588387,18.05005,16.511717,14.973383,13.438952,11.900618,12.138786,12.373051,12.611219,12.849388,13.087557,14.231546,15.371632,16.515621,17.655706,18.799696,16.218887,13.634172,11.053363,8.468649,5.8878384,5.35684,4.825841,4.298747,3.767748,3.2367494,2.795552,2.3543546,1.9092526,1.4680552,1.0268579,2.0263848,3.0259118,4.025439,5.024966,6.0244927,8.093826,10.159255,12.228588,14.294017,16.36335,14.551707,12.743969,10.932326,9.120684,7.3129454,6.1884775,5.0640097,3.9356375,2.8111696,1.6867018,1.7218413,1.756981,1.7921207,1.8272603,1.8623998,1.7647898,1.6671798,1.5695697,1.4719596,1.3743496,2.5573835,3.7404175,4.9234514,6.1064854,7.2856145,6.649197,6.012779,5.376362,4.73604,4.0996222,5.02887,5.9542136,6.883461,7.8088045,8.738052,7.6682463,6.602344,5.5364423,4.466636,3.4007344,3.611572,3.8185053,4.029343,4.240181,4.4510183,4.0761957,3.7052777,3.3343596,2.959537,2.5886188,2.5612879,2.533957,2.5066261,2.4792955,2.4480603,2.4207294,2.3894942,2.358259,2.330928,2.2996929,1.8663043,1.4290112,0.9956226,0.5583295,0.12494087,0.12884527,0.13665408,0.14055848,0.14446288,0.14836729,0.13665408,0.12494087,0.113227665,0.10151446,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.19131571,0.38653582,0.57785153,0.76916724,0.96438736,0.78088045,0.60127795,0.42167544,0.24207294,0.062470436,0.06637484,0.06637484,0.07027924,0.07418364,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.46462387,0.92924774,1.3938715,1.8584955,2.3231194,1.9639144,1.6047094,1.2455044,0.8862993,0.5231899,0.42557985,0.3318742,0.23426414,0.13665408,0.039044023,0.06637484,0.09761006,0.12884527,0.15617609,0.18741131,0.3435874,0.4958591,0.6520352,0.80821127,0.96438736,0.8433509,0.7223144,0.60127795,0.48414588,0.3631094,0.44119745,0.5231899,0.60127795,0.6832704,0.76135844,1.0659018,1.3665408,1.6710842,1.9717231,2.2762666,2.174752,2.0732377,1.9756275,1.8741131,1.7765031,1.7023194,1.6281357,1.5578566,1.4836729,1.4133936,1.4836729,1.5539521,1.6242313,1.6906061,1.7608855,1.456342,1.1478943,0.8394465,0.5309987,0.22645533,0.23426414,0.24597734,0.25378615,0.26549935,0.27330816,0.41777104,0.5583295,0.7027924,0.8433509,0.9878138,0.97610056,0.96438736,0.94876975,0.93705654,0.92534333,1.0190489,1.116659,1.2103647,1.3040704,1.4016805,1.3157835,1.2298868,1.1439898,1.0580931,0.97610056,0.9019169,0.8316377,0.75745404,0.6832704,0.61299115,0.5622339,0.5114767,0.46071947,0.41386664,0.3631094,0.44900626,0.5309987,0.61689556,0.7027924,0.78868926,0.6637484,0.5427119,0.42167544,0.29673457,0.1756981,0.14836729,0.12494087,0.10151446,0.07418364,0.05075723,0.1835069,0.32016098,0.45681506,0.58956474,0.7262188,0.60518235,0.48414588,0.3631094,0.24597734,0.12494087,0.24597734,0.3631094,0.48414588,0.60518235,0.7262188,0.61689556,0.5036679,0.39434463,0.28502136,0.1756981,0.23816854,0.30454338,0.3709182,0.43338865,0.4997635,0.45681506,0.40996224,0.3631094,0.32016098,0.27330816,0.21864653,0.1639849,0.10932326,0.05466163,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.039044023,0.05466163,0.07027924,0.08589685,0.10151446,0.10541886,0.10932326,0.113227665,0.12103647,0.12494087,0.14055848,0.15617609,0.1717937,0.1835069,0.19912452,0.1717937,0.14055848,0.10932326,0.078088045,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.3318742,0.46071947,0.58956474,0.71841,0.8511597,1.2181735,1.5851873,1.9522011,2.3192148,2.6862288,2.5378613,2.3855898,2.2372224,2.0888553,1.9365835,2.077142,2.2177005,2.358259,2.4988174,2.639376,3.1469483,3.6584249,4.165997,4.677474,5.1889505,5.466163,5.74728,6.028397,6.3056097,6.5867267,6.7311897,6.8756523,7.0240197,7.168483,7.3129454,7.47693,7.6409154,7.8088045,7.9727893,8.136774,8.339804,8.542832,8.745861,8.94889,9.151918,8.980125,8.8083315,8.640442,8.468649,8.300759,8.566258,8.831758,9.093353,9.358852,9.6243515,9.140205,8.65606,8.171914,7.6838636,7.1997175,6.098676,4.9937305,3.892689,2.7916477,1.6867018,1.5031948,1.3235924,1.1400855,0.95657855,0.77307165,0.7262188,0.679366,0.63251317,0.58566034,0.5388075,0.48414588,0.43338865,0.37872702,0.3279698,0.27330816,0.21864653,0.1639849,0.10932326,0.05466163,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.042948425,0.08589685,0.12884527,0.1717937,0.21083772,0.45291066,0.6910792,0.93315214,1.1713207,1.4133936,1.4719596,1.53443,1.5929961,1.6515622,1.7140326,1.7413634,1.7686942,1.796025,1.8233559,1.8506867,1.8506867,1.8545911,1.8584955,1.8584955,1.8623998,2.135708,2.4090161,2.67842,2.951728,3.2250361,3.7989833,4.376835,4.950782,5.5247293,6.098676,6.524256,6.949836,7.375416,7.800996,8.226576,7.800996,7.37932,6.957645,6.5359693,6.114294,6.1884775,6.262661,6.336845,6.4110284,6.4891167,7.2856145,8.086017,8.886419,9.686822,10.487225,11.00651,11.525795,12.0489855,12.568271,13.087557,13.845011,14.602465,15.359919,16.117373,16.874826,19.479063,22.079395,24.683632,27.283962,29.888199,30.493382,31.102468,31.711555,32.31674,32.925823,35.131813,37.3417,39.54769,41.753677,43.96357,48.32869,52.693813,57.058933,61.424057,65.78918,67.17524,68.5613,69.95127,71.33733,72.7234,68.93613,65.14886,61.361588,57.574314,53.787045,49.511726,45.236404,40.961082,36.685764,32.41435,31.079042,29.743736,28.40843,27.073126,25.73782,24.46108,23.188246,21.911505,20.63867,19.36193,17.624472,15.8870125,14.149553,12.412095,10.674636,10.061645,9.448653,8.835662,8.226576,7.6135845,7.719003,7.8283267,7.9337454,8.043069,8.148487,7.859562,7.570636,7.28171,6.98888,6.699954,6.8287997,6.9537406,7.082586,7.211431,7.336372,7.5120697,7.687768,7.8634663,8.039165,8.210958,7.9610763,7.7111945,7.461313,7.211431,6.9615493,6.735094,6.5086384,6.278279,6.0518236,5.825368,6.1025805,6.379793,6.657006,6.9342184,7.211431,7.055255,6.899079,6.7389984,6.5828223,6.426646,6.2587566,6.094772,5.930787,5.7668023,5.5989127,6.4695945,7.3402762,8.210958,9.081639,9.948417,11.115833,12.28325,13.450665,14.618082,15.789403,16.56638,17.343355,18.12033,18.897306,19.674282,20.502016,21.32975,22.157482,22.985216,23.81295,24.066736,24.324427,24.578213,24.831999,25.085785,23.996456,22.907127,21.8178,20.728472,19.639143,19.322887,19.00663,18.694279,18.378021,18.061766,17.440966,16.816261,16.195461,15.570756,14.949956,14.56342,14.180789,13.794253,13.411622,13.025085,13.739592,14.454097,15.168603,15.883108,16.601519,17.155943,17.714273,18.272602,18.830933,19.389261,18.299932,17.210606,16.125181,15.035853,13.950429,15.641035,17.335546,19.026152,20.720663,22.411268,20.689428,18.963682,17.237936,15.51219,13.786445,14.274494,14.762545,15.250595,15.738646,16.226696,16.218887,16.214983,16.211079,16.20327,16.199366,13.993378,11.791295,9.585307,7.37932,5.173333,5.040583,4.911738,4.7789884,4.646239,4.513489,3.7911747,3.0727646,2.3543546,1.6320401,0.9136301,2.0380979,3.1625657,4.2870336,5.4115014,6.5359693,7.605776,8.675582,9.749292,10.819098,11.888905,11.197825,10.506746,9.815667,9.128492,8.437413,7.238762,6.036206,4.8375545,3.638903,2.436347,2.5027218,2.5690966,2.631567,2.697942,2.7643168,2.6237583,2.4831998,2.3426414,2.2020829,2.0615244,3.8302186,5.5989127,7.363703,9.132397,10.901091,9.788337,8.675582,7.562827,6.4500723,5.337318,6.883461,8.433509,9.979652,11.525795,13.075843,11.365715,9.659492,7.9532676,6.2431393,4.5369153,4.2284675,3.9161155,3.6076677,3.2992198,2.9868677,2.7330816,2.4831998,2.2294137,1.9756275,1.7257458,2.0263848,2.330928,2.631567,2.9361105,3.2367494,3.2562714,3.2718892,3.2914112,3.3070288,3.3265507,2.697942,2.069333,1.4407244,0.8160201,0.18741131,0.1717937,0.15227169,0.13665408,0.11713207,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.19522011,0.39044023,0.58566034,0.78088045,0.97610056,0.79259366,0.60908675,0.42557985,0.24597734,0.062470436,0.058566034,0.058566034,0.05466163,0.05075723,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.59737355,1.1947471,1.7921207,2.3894942,2.9868677,2.533957,2.0810463,1.6281357,1.1791295,0.7262188,0.58566034,0.44510186,0.30454338,0.1639849,0.023426414,0.046852827,0.06637484,0.08589685,0.10541886,0.12494087,0.359205,0.58956474,0.8238289,1.0541886,1.2884527,1.1088502,0.92924774,0.74574083,0.5661383,0.38653582,0.5309987,0.679366,0.8238289,0.96829176,1.1127546,1.5617609,2.0068626,2.455869,2.900971,3.349977,3.2016098,3.049338,2.900971,2.7486992,2.6003318,2.4988174,2.3933985,2.2918842,2.1903696,2.0888553,1.9170616,1.7491722,1.5773785,1.4055848,1.2376955,1.0580931,0.8784905,0.698888,0.5192855,0.3357786,0.3513962,0.3670138,0.38263142,0.39824903,0.41386664,0.62079996,0.8277333,1.0346665,1.2415999,1.4485333,1.43682,1.4251068,1.4133936,1.4016805,1.3860629,1.5305257,1.6710842,1.815547,1.9561055,2.1005683,1.9717231,1.8467822,1.717937,1.5890918,1.4641509,1.2845483,1.1088502,0.92924774,0.75354964,0.57394713,0.5114767,0.44900626,0.38653582,0.3240654,0.26159495,0.42557985,0.59346914,0.75745404,0.92143893,1.0893283,0.92143893,0.75745404,0.59346914,0.42557985,0.26159495,0.22645533,0.18741131,0.14836729,0.113227665,0.07418364,0.27721256,0.48024148,0.6832704,0.8862993,1.0893283,0.9058213,0.7262188,0.5466163,0.3670138,0.18741131,0.3670138,0.5466163,0.7262188,0.9058213,1.0893283,0.92143893,0.75745404,0.59346914,0.42557985,0.26159495,0.359205,0.45681506,0.5544251,0.6520352,0.74964523,0.6832704,0.61689556,0.5466163,0.48024148,0.41386664,0.3318742,0.24597734,0.1639849,0.08199245,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.019522011,0.027330816,0.03513962,0.042948425,0.05075723,0.05075723,0.05466163,0.058566034,0.058566034,0.062470436,0.07027924,0.078088045,0.08589685,0.093705654,0.10151446,0.08589685,0.07027924,0.05466163,0.039044023,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.21474212,0.3318742,0.44510186,0.5583295,0.6754616,1.0268579,1.3782539,1.7335546,2.084951,2.436347,2.338737,2.2372224,2.135708,2.0380979,1.9365835,2.069333,2.2020829,2.3348327,2.4675822,2.6003318,3.0415294,3.4866312,3.9278288,4.369026,4.814128,5.165524,5.5169206,5.8683167,6.223617,6.575013,6.6843367,6.79366,6.9068875,7.016211,7.125534,7.1841,7.238762,7.297328,7.355894,7.4105554,7.558923,7.703386,7.8478484,7.9923115,8.136774,8.113348,8.093826,8.070399,8.046973,8.023546,8.308568,8.589685,8.870802,9.155824,9.43694,8.905942,8.378847,7.8478484,7.3168497,6.785851,5.794133,4.7985106,3.802888,2.8072653,1.8116426,1.6281357,1.4407244,1.2572175,1.0737107,0.8862993,0.80821127,0.7262188,0.6481308,0.5661383,0.48805028,0.41777104,0.3474918,0.27721256,0.20693332,0.13665408,0.10932326,0.08199245,0.05466163,0.027330816,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.3709182,0.5388075,0.7106012,0.8784905,1.0502841,1.2298868,1.4094892,1.5890918,1.7686942,1.9482968,1.9443923,1.9404879,1.9365835,1.9287747,1.9248703,1.9443923,1.9639144,1.9834363,2.0068626,2.0263848,2.3426414,2.6588979,2.979059,3.2953155,3.611572,4.173806,4.73604,5.298274,5.8644123,6.426646,6.7389984,7.0513506,7.363703,7.676055,7.988407,7.519879,7.0513506,6.5867267,6.1181984,5.64967,5.899552,6.1494336,6.3993154,6.649197,6.899079,7.773665,8.648251,9.526741,10.401327,11.275913,11.674163,12.068507,12.466757,12.8650055,13.263254,14.286208,15.309161,16.32821,17.351164,18.374117,21.431265,24.48841,27.549461,30.60661,33.663757,33.59738,33.531006,33.468536,33.40216,33.335785,36.022015,38.708244,41.394474,44.076797,46.763027,51.30775,55.852474,60.397198,64.941925,69.48665,70.6892,71.887856,73.0865,74.28906,75.48772,71.411514,67.339226,63.26303,59.186832,55.110638,50.874363,46.638084,42.40181,38.16163,33.92535,32.46901,31.016571,29.56023,28.103888,26.65145,25.1873,23.723148,22.262901,20.79875,19.338505,17.31212,15.285735,13.263254,11.23687,9.21439,8.550641,7.8868923,7.223144,6.5633,5.899552,6.0713453,6.2431393,6.4188375,6.590631,6.7624245,6.606249,6.446168,6.289992,6.133816,5.9737353,6.168956,6.364176,6.559396,6.754616,6.949836,7.0630636,7.1762915,7.2856145,7.3988423,7.5120697,7.238762,6.9615493,6.688241,6.4110284,6.13772,5.9425,5.74728,5.55206,5.35684,5.1616197,5.571582,5.9776397,6.3836975,6.79366,7.1997175,7.039637,6.8795567,6.719476,6.559396,6.3993154,6.0908675,5.786324,5.477876,5.169429,4.860981,5.883934,6.9068875,7.929841,8.952794,9.975748,11.240774,12.5058,13.770826,15.035853,16.300879,16.995863,17.690847,18.38583,19.080814,19.775797,20.544964,21.314133,22.0833,22.85637,23.625538,23.816854,24.004265,24.195581,24.386896,24.574308,23.74267,22.911032,22.079395,21.243853,20.412214,19.978827,19.549341,19.115953,18.682566,18.249176,17.468296,16.69132,15.9104395,15.129559,14.348679,13.958238,13.563893,13.173453,12.779109,12.388668,12.630741,12.8767185,13.122696,13.368673,13.610746,14.735214,15.855778,16.980246,18.10081,19.225277,18.214037,17.198893,16.187653,15.176412,14.161267,16.378967,18.592764,20.80656,23.02426,25.238056,23.3249,21.411741,19.498585,17.589333,15.676175,16.414106,17.148134,17.886066,18.623999,19.36193,18.210133,17.058334,15.906535,14.750832,13.599033,11.771772,9.944512,8.117252,6.289992,4.462732,4.728231,4.9937305,5.2592297,5.520825,5.786324,4.7907014,3.7911747,2.795552,1.796025,0.80040246,2.0498111,3.2992198,4.548629,5.801942,7.0513506,7.1216297,7.195813,7.266093,7.3402762,7.4105554,7.843944,8.273428,8.702912,9.132397,9.561881,8.289046,7.012306,5.735567,4.462732,3.1859922,3.2836022,3.377308,3.4710135,3.5686235,3.6623292,3.4788225,3.2992198,3.1157131,2.9322062,2.7486992,5.1030536,7.453504,9.807858,12.158309,14.512663,12.923572,11.338385,9.749292,8.164105,6.575013,8.741957,10.9089,13.075843,15.246691,17.413633,15.063184,12.716639,10.370092,8.023546,5.6730967,4.845363,4.0137253,3.1859922,2.3543546,1.5266213,1.3938715,1.261122,1.1283722,0.9956226,0.8628729,1.4953861,2.1278992,2.7604125,3.3929255,4.025439,4.0918136,4.154284,4.220659,4.283129,4.349504,3.5295796,2.7096553,1.8897307,1.0698062,0.24988174,0.21083772,0.1717937,0.12884527,0.08980125,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.19912452,0.39434463,0.59346914,0.78868926,0.9878138,0.80430686,0.61689556,0.43338865,0.24597734,0.062470436,0.05466163,0.046852827,0.039044023,0.031235218,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.7301232,1.4602464,2.1903696,2.920493,3.6506162,3.1039999,2.5612879,2.0146716,1.4680552,0.92534333,0.7418364,0.5583295,0.37872702,0.19522011,0.011713207,0.023426414,0.031235218,0.042948425,0.05075723,0.062470436,0.3709182,0.6832704,0.9917182,1.3040704,1.6125181,1.3743496,1.1322767,0.8941081,0.6520352,0.41386664,0.62079996,0.8316377,1.0424755,1.2533131,1.4641509,2.0537157,2.6471848,3.240654,3.8341231,4.423688,4.224563,4.025439,3.8263142,3.6232853,3.4241607,3.2914112,3.1586614,3.0259118,2.893162,2.7643168,2.3543546,1.9443923,1.53443,1.1244678,0.7106012,0.659844,0.60908675,0.5544251,0.5036679,0.44900626,0.46852827,0.48805028,0.5114767,0.5309987,0.5505207,0.8238289,1.0932326,1.3665408,1.639849,1.9131571,1.901444,1.8858263,1.8741131,1.8623998,1.8506867,2.0380979,2.2294137,2.4207294,2.6081407,2.7994564,2.631567,2.4597735,2.2918842,2.1200905,1.9482968,1.6671798,1.3860629,1.1010414,0.8199245,0.5388075,0.46071947,0.38653582,0.31235218,0.23816854,0.1639849,0.40605783,0.6520352,0.8980125,1.1439898,1.3860629,1.1791295,0.97219616,0.76526284,0.5583295,0.3513962,0.30063897,0.24988174,0.19912452,0.14836729,0.10151446,0.3709182,0.64032197,0.9097257,1.1791295,1.4485333,1.2103647,0.96829176,0.7301232,0.49195468,0.24988174,0.49195468,0.7301232,0.96829176,1.2103647,1.4485333,1.2298868,1.0112402,0.78868926,0.5700427,0.3513962,0.48024148,0.60908675,0.7418364,0.8706817,0.999527,0.9097257,0.8199245,0.7301232,0.64032197,0.5505207,0.44119745,0.3318742,0.21864653,0.10932326,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.8394465,1.175225,1.5110037,1.8506867,2.1864653,2.135708,2.0888553,2.0380979,1.9873407,1.9365835,2.0615244,2.1864653,2.3114061,2.436347,2.5612879,2.9361105,3.310933,3.6857557,4.0605783,4.4393053,4.860981,5.2865605,5.7121406,6.13772,6.5633,6.6374836,6.7116675,6.785851,6.8639393,6.9381227,6.8873653,6.8366084,6.785851,6.7389984,6.688241,6.774138,6.8639393,6.949836,7.0357327,7.125534,7.250475,7.375416,7.5003567,7.6252975,7.7502384,8.050878,8.351517,8.648251,8.94889,9.249529,8.675582,8.101635,7.523783,6.949836,6.375889,5.4856853,4.5993857,3.7130866,2.8267872,1.9365835,1.7491722,1.5617609,1.3743496,1.1869383,0.999527,0.8862993,0.77307165,0.6637484,0.5505207,0.43729305,0.3513962,0.26159495,0.1756981,0.08589685,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.28892577,0.38653582,0.48805028,0.58566034,0.6871748,0.9878138,1.2884527,1.5890918,1.8858263,2.1864653,2.1513257,2.1122816,2.0732377,2.0380979,1.999054,2.0380979,2.0732377,2.1122816,2.1513257,2.1864653,2.5495746,2.912684,3.2757936,3.638903,3.998108,4.548629,5.099149,5.64967,6.2001905,6.7507114,6.949836,7.1489606,7.348085,7.551114,7.7502384,7.238762,6.7233806,6.211904,5.700427,5.1889505,5.610626,6.036206,6.461786,6.8873653,7.3129454,8.261715,9.21439,10.163159,11.111929,12.0606985,12.337912,12.611219,12.888432,13.16174,13.438952,14.723501,16.011953,17.300406,18.58886,19.873407,23.38737,26.90133,30.411388,33.92535,37.439312,36.70138,35.963448,35.225517,34.487587,33.749653,36.91222,40.074783,43.23735,46.399918,49.56248,54.286808,59.011135,63.73937,68.46369,73.18802,74.19926,75.2144,76.22565,77.236885,78.24812,73.88691,69.52569,65.16057,60.79935,56.438133,52.237,48.035862,43.838627,39.637493,35.436356,33.86288,32.289406,30.712029,29.138554,27.561176,25.913517,24.261955,22.614298,20.962736,19.311174,16.999767,14.688361,12.373051,10.061645,7.7502384,7.0357327,6.3251314,5.610626,4.900025,4.1894236,4.423688,4.661856,4.900025,5.138193,5.376362,5.349031,5.3256044,5.298274,5.2748475,5.251421,5.5130157,5.774611,6.036206,6.3017054,6.5633,6.6140575,6.66091,6.7116675,6.7624245,6.813182,6.5125427,6.211904,5.911265,5.610626,5.3138914,5.1499066,4.985922,4.825841,4.661856,4.5017757,5.036679,5.575486,6.114294,6.649197,7.1880045,7.0240197,6.8639393,6.699954,6.5359693,6.375889,5.9268827,5.473972,5.024966,4.575959,4.123049,5.298274,6.473499,7.648724,8.823949,9.999174,11.361811,12.724447,14.087084,15.449719,16.812357,17.425346,18.038338,18.651329,19.26432,19.873407,20.587914,21.298513,22.01302,22.723621,23.438128,23.563068,23.68801,23.81295,23.937891,24.062832,23.488884,22.911032,22.337086,21.763138,21.189192,20.63867,20.08815,19.537628,18.987108,18.436588,17.49953,16.562475,15.625418,14.688361,13.751305,13.349152,12.950902,12.548749,12.150499,11.748346,11.525795,11.29934,11.076789,10.850334,10.6238785,12.314485,14.001186,15.687888,17.37459,19.061293,18.124235,17.18718,16.250122,15.313066,14.376009,17.112995,19.849981,22.586967,25.323954,28.06094,25.964275,23.863707,21.763138,19.662569,17.562002,18.549814,19.537628,20.525442,21.513256,22.50107,20.201378,17.901684,15.598087,13.298394,10.998701,9.550168,8.101635,6.649197,5.2006636,3.7482262,4.4119744,5.0757227,5.7394714,6.3993154,7.0630636,5.786324,4.513489,3.2367494,1.9639144,0.6871748,2.0615244,3.435874,4.814128,6.1884775,7.562827,6.6374836,5.7121406,4.786797,3.8614538,2.9361105,4.4861584,6.036206,7.5862536,9.136301,10.686349,9.339331,7.988407,6.6374836,5.2865605,3.9356375,4.0605783,4.1894236,4.3143644,4.4393053,4.564246,4.337791,4.1113358,3.8887846,3.6623292,3.435874,6.375889,9.311999,12.252014,15.188125,18.124235,16.062712,14.001186,11.935758,9.874233,7.812709,10.600452,13.388195,16.175938,18.963682,21.751425,18.760653,15.773785,12.786918,9.80005,6.813182,5.462259,4.1113358,2.7643168,1.4133936,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.96438736,1.9248703,2.8892577,3.8497405,4.814128,4.9234514,5.036679,5.1499066,5.263134,5.376362,4.3612175,3.349977,2.338737,1.3235924,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.19912452,0.39824903,0.60127795,0.80040246,0.999527,0.81211567,0.62470436,0.43729305,0.24988174,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.8628729,1.7257458,2.5886188,3.4514916,4.3143644,3.6740425,3.0376248,2.4012074,1.7608855,1.1244678,0.9019169,0.6754616,0.44900626,0.22645533,0.0,0.0,0.0,0.0,0.0,0.0,0.38653582,0.77307165,1.1635119,1.5500476,1.9365835,1.6359446,1.33921,1.038571,0.737932,0.43729305,0.7106012,0.9878138,1.261122,1.5383345,1.8116426,2.5495746,3.2875066,4.025439,4.7633705,5.5013027,5.251421,5.001539,4.7516575,4.5017757,4.251894,4.087909,3.9239242,3.7638438,3.5998588,3.435874,2.787743,2.135708,1.4875772,0.8394465,0.18741131,0.26159495,0.3357786,0.41386664,0.48805028,0.5622339,0.58566034,0.61299115,0.63641757,0.6637484,0.6871748,1.0268579,1.3626363,1.698415,2.0380979,2.3738766,2.3621633,2.35045,2.338737,2.3231194,2.3114061,2.5495746,2.787743,3.0259118,3.2640803,3.4983444,3.2875066,3.076669,2.8619268,2.6510892,2.436347,2.0498111,1.6632754,1.2767396,0.8862993,0.4997635,0.41386664,0.3240654,0.23816854,0.14836729,0.062470436,0.38653582,0.7106012,1.038571,1.3626363,1.6867018,1.43682,1.1869383,0.93705654,0.6871748,0.43729305,0.37482262,0.31235218,0.24988174,0.18741131,0.12494087,0.46071947,0.80040246,1.1361811,1.475864,1.8116426,1.5110037,1.2142692,0.9136301,0.61299115,0.31235218,0.61299115,0.9136301,1.2142692,1.5110037,1.8116426,1.5383345,1.261122,0.9878138,0.7106012,0.43729305,0.60127795,0.76135844,0.92534333,1.0893283,1.2494087,1.1361811,1.0268579,0.9136301,0.80040246,0.6871748,0.5505207,0.41386664,0.27330816,0.13665408,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09761006,0.19522011,0.29283017,0.39044023,0.48805028,0.79649806,1.1088502,1.4172981,1.7257458,2.0380979,2.0380979,2.0380979,2.0380979,2.0380979,2.0380979,2.15523,2.2723622,2.3894942,2.5066261,2.6237583,2.9634414,3.3031244,3.6467118,3.9863946,4.3260775,4.7243266,5.1186714,5.5169206,5.9151692,6.3134184,6.336845,6.364176,6.387602,6.4110284,6.4383593,6.329036,6.223617,6.114294,6.008875,5.899552,6.168956,6.434455,6.703859,6.969358,7.238762,7.4417906,7.6409154,7.843944,8.046973,8.250002,8.378847,8.511597,8.640442,8.769287,8.898132,8.19534,7.4886436,6.785851,6.0791545,5.376362,4.6345253,3.8965936,3.154757,2.416825,1.6749885,1.5110037,1.3509232,1.1869383,1.0268579,0.8628729,0.76135844,0.6559396,0.5544251,0.45291066,0.3513962,0.28111696,0.21083772,0.14055848,0.07027924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.06637484,0.09761006,0.12884527,0.1639849,0.28111696,0.39824903,0.5153811,0.63251317,0.74964523,1.0346665,1.319688,1.6047094,1.8897307,2.174752,2.2567444,2.3348327,2.416825,2.494913,2.5769055,2.6667068,2.7604125,2.854118,2.9439192,3.0376248,3.3265507,3.611572,3.900498,4.1894236,4.474445,4.9468775,5.4154058,5.883934,6.356367,6.824895,7.113821,7.3988423,7.687768,7.9766936,8.261715,7.8205175,7.37932,6.9342184,6.493021,6.0518236,6.2938967,6.5359693,6.7780423,7.0201154,7.262188,8.113348,8.960603,9.811763,10.662923,11.514082,11.861574,12.212971,12.564366,12.911859,13.263254,14.426766,15.586374,16.749886,17.913397,19.073006,22.196527,25.32005,28.443571,31.563189,34.68671,34.046387,33.40216,32.757935,32.117615,31.473387,33.944874,36.41636,38.88394,41.35543,43.82301,47.727413,51.62791,55.532314,59.43281,63.33721,64.34846,65.35579,66.36703,67.37827,68.385605,64.91459,61.443577,57.96866,54.497646,51.022728,47.579044,44.13146,40.683872,37.236286,33.788696,32.30893,30.82916,29.345488,27.865719,26.38595,24.476698,22.563541,20.650383,18.737226,16.82407,15.035853,13.243732,11.455516,9.663396,7.8751793,7.3441806,6.813182,6.2860875,5.755089,5.22409,5.2436123,5.2592297,5.278752,5.2943697,5.3138914,5.35684,5.395884,5.4388323,5.481781,5.5247293,5.84489,6.165051,6.4852123,6.805373,7.125534,7.0591593,6.996689,6.930314,6.8639393,6.801469,6.524256,6.250948,5.9737353,5.700427,5.423215,5.2475166,5.0718184,4.892216,4.716518,4.5369153,4.970304,5.4036927,5.833177,6.266566,6.699954,6.5554914,6.4110284,6.266566,6.1181984,5.9737353,5.7668023,5.559869,5.3529353,5.1460023,4.939069,6.04011,7.141152,8.246098,9.347139,10.44818,11.732729,13.013372,14.297921,15.578565,16.863113,17.511244,18.163279,18.81141,19.463446,20.111576,21.013493,21.911505,22.813423,23.711435,24.613352,24.949131,25.281004,25.616783,25.952562,26.28834,25.690968,25.097498,24.504028,23.906654,23.313187,22.337086,21.360985,20.388788,19.412687,18.436588,17.26917,16.101755,14.934339,13.766922,12.599506,12.212971,11.8303385,11.443803,11.061172,10.674636,10.612165,10.549695,10.487225,10.424754,10.362284,11.584361,12.802535,14.020708,15.242786,16.46096,15.914344,15.367727,14.821111,14.27059,13.723974,16.43363,19.13938,21.849035,24.554787,27.260536,24.980366,22.696291,20.416119,18.132044,15.847969,16.788929,17.72989,18.67085,19.611813,20.548868,18.631807,16.714746,14.797685,12.880623,10.963562,10.139732,9.315904,8.495979,7.6721506,6.8483214,6.8209906,6.79366,6.7663293,6.7389984,6.7116675,5.911265,5.1069584,4.3065557,3.5022488,2.7018464,4.2167544,5.7316628,7.2465706,8.761478,10.276386,8.769287,7.2582836,5.7511845,4.2440853,2.736986,4.73604,6.7389984,8.738052,10.737106,12.73616,12.127073,11.514082,10.901091,10.2881,9.675109,8.519405,7.3597984,6.2040954,5.044488,3.8887846,3.8380275,3.78727,3.736513,3.6857557,3.638903,5.9815445,8.32809,10.670732,13.017277,15.363823,13.575606,11.787391,9.999174,8.210958,6.426646,8.823949,11.221252,13.618555,16.015858,18.41316,16.09785,13.786445,11.475039,9.163632,6.8483214,5.6809053,4.5095844,3.338264,2.1708477,0.999527,1.077615,1.1557031,1.2337911,1.3118792,1.3860629,1.9404879,2.4910088,3.0454338,3.5959544,4.1503797,4.181615,4.2167544,4.2479897,4.279225,4.3143644,3.5608149,2.8072653,2.0537157,1.3040704,0.5505207,0.7262188,0.9019169,1.0737107,1.2494087,1.4251068,1.3782539,1.3314011,1.2806439,1.2337911,1.1869383,1.4133936,1.6437533,1.8702087,2.096664,2.3270237,2.5300527,2.736986,2.9400148,3.1469483,3.349977,3.1391394,2.9243972,2.7135596,2.4988174,2.2879796,2.233318,2.182561,2.1318035,2.077142,2.0263848,1.7804074,1.53443,1.2884527,1.0463798,0.80040246,1.4446288,2.0888553,2.7330816,3.3812122,4.025439,3.4983444,2.97125,2.4441557,1.9131571,1.3860629,1.1439898,0.8980125,0.6520352,0.40605783,0.1639849,0.29673457,0.42557985,0.5583295,0.6910792,0.8238289,1.0698062,1.3157835,1.5617609,1.8038338,2.0498111,1.8467822,1.6437533,1.4407244,1.2415999,1.038571,1.5656652,2.096664,2.6276627,3.1586614,3.6857557,4.298747,4.911738,5.5247293,6.13772,6.7507114,6.239235,5.7316628,5.2201858,4.7087092,4.2011366,4.0918136,3.9863946,3.8770714,3.7716527,3.6623292,3.1430438,2.6276627,2.1083772,1.5929961,1.0737107,1.0268579,0.97610056,0.92534333,0.8745861,0.8238289,0.8589685,0.8941081,0.92924774,0.96438736,0.999527,1.5773785,2.15523,2.7330816,3.310933,3.8887846,3.951255,4.01763,4.084005,4.1464753,4.21285,4.173806,4.138666,4.0996222,4.0644827,4.025439,3.8302186,3.6349986,3.4397783,3.2445583,3.049338,2.7643168,2.475391,2.1864653,1.901444,1.6125181,1.5110037,1.4094892,1.3040704,1.2025559,1.1010414,1.261122,1.4251068,1.5890918,1.7491722,1.9131571,1.6593709,1.4055848,1.1557031,0.9019169,0.6481308,0.57785153,0.5036679,0.43338865,0.359205,0.28892577,0.5231899,0.76135844,0.999527,1.2376955,1.475864,1.2337911,0.9917182,0.74574083,0.5036679,0.26159495,0.5036679,0.74574083,0.9917182,1.2337911,1.475864,1.2533131,1.0307622,0.80821127,0.58566034,0.3631094,0.4958591,0.62860876,0.76135844,0.8941081,1.0268579,0.93315214,0.8433509,0.75354964,0.6637484,0.57394713,0.46071947,0.3513962,0.23816854,0.12494087,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.093705654,0.19131571,0.28502136,0.37872702,0.47633708,0.75745404,1.038571,1.3235924,1.6047094,1.8858263,1.9365835,1.9873407,2.0380979,2.0888553,2.135708,2.2489357,2.358259,2.4675822,2.5769055,2.6862288,2.9907722,3.2992198,3.6037633,3.9083066,4.21285,4.5837684,4.950782,5.3217,5.6926184,6.0635366,6.036206,6.012779,5.989353,5.9620223,5.938596,5.7707067,5.606722,5.4427366,5.278752,5.1108627,5.559869,6.008875,6.453977,6.902983,7.348085,7.629202,7.910319,8.191436,8.468649,8.749765,8.710721,8.671678,8.628729,8.589685,8.550641,7.715099,6.8795567,6.044015,5.2084727,4.376835,3.7833657,3.1898966,2.5964274,2.0068626,1.4133936,1.2767396,1.1361811,0.999527,0.8628729,0.7262188,0.63251317,0.5388075,0.44900626,0.3553006,0.26159495,0.21083772,0.15617609,0.10541886,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.027330816,0.05466163,0.08199245,0.10932326,0.13665408,0.27330816,0.40605783,0.5427119,0.679366,0.81211567,1.0815194,1.3509232,1.6242313,1.893635,2.1630387,2.358259,2.5573835,2.7565079,2.951728,3.1508527,3.2992198,3.4436827,3.59205,3.7404175,3.8887846,4.0996222,4.3143644,4.5252023,4.73604,4.950782,5.3412223,5.7316628,6.1181984,6.5086384,6.899079,7.2739015,7.648724,8.023546,8.398369,8.773191,8.402273,8.031356,7.656533,7.2856145,6.910792,6.9732623,7.0318284,7.094299,7.152865,7.211431,7.9610763,8.710721,9.464272,10.213917,10.963562,11.389141,11.810817,12.236397,12.661977,13.087557,14.126127,15.160794,16.199366,17.237936,18.276506,21.005684,23.738766,26.471848,29.20493,31.938011,31.391394,30.840874,30.294256,29.74764,29.201025,30.977528,32.754032,34.53444,36.31094,38.087444,41.16802,44.248592,47.329163,50.409737,53.48641,54.493744,55.50108,56.508415,57.519653,58.52699,55.942276,53.361465,50.776752,48.195942,45.61123,42.91719,40.223152,37.529114,34.831173,32.137135,30.751072,29.368914,27.982851,26.596788,25.210726,23.035973,20.861221,18.68647,16.511717,14.336966,13.0719385,11.803008,10.534078,9.269051,8.00012,7.6526284,7.3051367,6.957645,6.610153,6.262661,6.0596323,5.8566036,5.6535745,5.4505453,5.251421,5.3607445,5.4700675,5.579391,5.688714,5.801942,6.1767645,6.5554914,6.9342184,7.309041,7.687768,7.5081654,7.328563,7.1489606,6.969358,6.785851,6.5359693,6.2860875,6.036206,5.786324,5.5364423,5.3451266,5.153811,4.958591,4.7672753,4.575959,4.903929,5.2318993,5.5559645,5.883934,6.211904,6.083059,5.958118,5.8292727,5.704332,5.575486,5.610626,5.645766,5.6809053,5.716045,5.7511845,6.7819467,7.8088045,8.839567,9.870329,10.901091,12.103647,13.306203,14.508759,15.711315,16.91387,17.601046,18.28822,18.975395,19.662569,20.349745,21.439074,22.524496,23.613825,24.69925,25.788576,26.33129,26.877905,27.420616,27.967234,28.51385,27.896954,27.283962,26.667067,26.054077,25.437181,24.0355,22.637724,21.236044,19.838268,18.436588,17.03881,15.641035,14.243259,12.849388,11.4516115,11.080693,10.709775,10.338858,9.971844,9.600925,9.698535,9.80005,9.901564,9.999174,10.100689,10.8542385,11.603884,12.357433,13.110983,13.860628,13.704452,13.548276,13.388195,13.232019,13.075843,15.754263,18.42878,21.107199,23.785618,26.464039,23.996456,21.532778,19.069101,16.601519,14.13784,15.031949,15.9221525,16.816261,17.706465,18.600573,17.066143,15.531713,13.993378,12.458947,10.924518,10.729298,10.534078,10.338858,10.143637,9.948417,9.2339115,8.515501,7.7970915,7.0786815,6.364176,6.0323014,5.704332,5.3724575,5.040583,4.7126136,6.36808,8.023546,9.679013,11.330575,12.986042,10.897186,8.8083315,6.715572,4.6267166,2.5378613,4.985922,7.437886,9.885946,12.337912,14.785972,14.9109125,15.035853,15.160794,15.285735,15.410676,12.970425,10.534078,8.093826,5.6535745,3.213323,3.338264,3.4632049,3.5881457,3.7130866,3.8380275,5.591104,7.3441806,9.093353,10.84643,12.599506,11.088503,9.573594,8.062591,6.551587,5.036679,7.043542,9.054309,11.061172,13.068034,15.074897,13.438952,11.799104,10.163159,8.52331,6.8873653,5.8956475,4.9078336,3.9161155,2.9283018,1.9365835,2.1044729,2.2723622,2.4402514,2.6081407,2.77603,2.9165885,3.0610514,3.2016098,3.3460727,3.4866312,3.4397783,3.3929255,3.3460727,3.2992198,3.2484627,2.7565079,2.2645533,1.7725986,1.2806439,0.78868926,1.1986516,1.6125181,2.0263848,2.436347,2.8502135,2.7291772,2.6081407,2.4910088,2.3699722,2.2489357,2.7291772,3.2094188,3.68966,4.169902,4.650143,4.860981,5.0718184,5.278752,5.4895897,5.700427,5.462259,5.22409,4.985922,4.7516575,4.513489,4.4197836,4.3260775,4.2362766,4.142571,4.0488653,3.5608149,3.06886,2.5808098,2.0888553,1.6008049,2.0263848,2.455869,2.8814487,3.310933,3.736513,3.3187418,2.900971,2.4831998,2.069333,1.6515622,1.3860629,1.1205635,0.8550641,0.58956474,0.3240654,0.58956474,0.8550641,1.1205635,1.3860629,1.6515622,1.7530766,1.8545911,1.9561055,2.0615244,2.1630387,2.05762,1.9522011,1.8467822,1.7413634,1.6359446,2.4207294,3.2055142,3.9942036,4.7789884,5.563773,6.0518236,6.5359693,7.0240197,7.5120697,8.00012,7.230953,6.461786,5.688714,4.919547,4.1503797,4.095718,4.044961,3.9942036,3.9395418,3.8887846,3.5022488,3.1157131,2.7330816,2.3465457,1.9639144,1.7882162,1.6125181,1.43682,1.261122,1.0893283,1.1322767,1.1791295,1.2220778,1.2689307,1.3118792,2.1318035,2.9478238,3.7638438,4.5837684,5.3997884,5.5442514,5.6848097,5.8292727,5.969831,6.114294,5.7980375,5.4856853,5.173333,4.860981,4.548629,4.3729305,4.193328,4.01763,3.8419318,3.6623292,3.474918,3.2875066,3.1000953,2.912684,2.7252727,2.6081407,2.4910088,2.3738766,2.2567444,2.135708,2.135708,2.135708,2.135708,2.135708,2.135708,1.8819219,1.6281357,1.3743496,1.116659,0.8628729,0.78088045,0.698888,0.61689556,0.5309987,0.44900626,0.58566034,0.7262188,0.8628729,0.999527,1.1361811,0.95267415,0.76916724,0.58175594,0.39824903,0.21083772,0.39824903,0.58175594,0.76916724,0.95267415,1.1361811,0.96829176,0.79649806,0.62860876,0.45681506,0.28892577,0.39044023,0.49195468,0.59346914,0.698888,0.80040246,0.7340276,0.6637484,0.59737355,0.5309987,0.46071947,0.37482262,0.28892577,0.19912452,0.113227665,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.14836729,0.14836729,0.14836729,0.14836729,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.093705654,0.1835069,0.27721256,0.3709182,0.46071947,0.71841,0.97219616,1.2259823,1.4836729,1.737459,1.8389735,1.9365835,2.0380979,2.135708,2.2372224,2.338737,2.4441557,2.5456703,2.6471848,2.7486992,3.018103,3.2914112,3.5608149,3.8302186,4.0996222,4.4432096,4.786797,5.12648,5.4700675,5.813655,5.735567,5.661383,5.5871997,5.5130157,5.4388323,5.2162814,4.9937305,4.7711797,4.548629,4.3260775,4.950782,5.579391,6.2079997,6.8366084,7.461313,7.8205175,8.175818,8.535024,8.894228,9.249529,9.0386915,8.831758,8.62092,8.410083,8.1992445,7.2348576,6.27047,5.3060827,4.3416953,3.3734035,2.9283018,2.4831998,2.0380979,1.5969005,1.1517987,1.038571,0.92534333,0.81211567,0.698888,0.58566034,0.5036679,0.42167544,0.339683,0.25769055,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.26549935,0.41777104,0.5700427,0.7223144,0.8745861,1.1283722,1.3860629,1.639849,1.893635,2.1513257,2.463678,2.7799344,3.096191,3.408543,3.7247996,3.9278288,4.1308575,4.3338866,4.5369153,4.73604,4.8765984,5.0132523,5.1499066,5.2865605,5.423215,5.735567,6.044015,6.356367,6.6648145,6.9732623,7.437886,7.898606,8.36323,8.823949,9.288573,8.98403,8.683391,8.378847,8.078208,7.773665,7.6526284,7.531592,7.406651,7.2856145,7.1606736,7.812709,8.460839,9.112875,9.761005,10.413041,10.912805,11.412568,11.912332,12.412095,12.911859,13.825488,14.739119,15.648844,16.562475,17.476105,19.818747,22.161386,24.504028,26.84667,29.189312,28.7364,28.28349,27.83058,27.377668,26.924759,28.010181,29.095606,30.18103,31.266453,32.347973,34.60862,36.865368,39.122112,41.378857,43.6356,44.642937,45.646366,46.6537,47.657135,48.660564,46.96996,45.275448,43.584843,41.89033,40.199726,38.25924,36.314846,34.370453,32.429966,30.485573,29.19712,27.908667,26.61631,25.327858,24.039404,21.599154,19.162806,16.72646,14.286208,11.849861,11.10412,10.358379,9.616543,8.870802,8.125061,7.9610763,7.793187,7.629202,7.465217,7.3012323,6.8756523,6.453977,6.0323014,5.610626,5.1889505,5.364649,5.5442514,5.7199492,5.8956475,6.0752497,6.5086384,6.9459314,7.37932,7.816613,8.250002,7.9532676,7.660437,7.363703,7.0708723,6.774138,6.551587,6.3251314,6.098676,5.8761253,5.64967,5.4427366,5.2358036,5.02887,4.8219366,4.6110992,4.83365,5.056201,5.278752,5.5013027,5.7238536,5.6145306,5.505207,5.395884,5.2865605,5.173333,5.45445,5.7316628,6.008875,6.2860875,6.5633,7.519879,8.476458,9.43694,10.393518,11.350098,12.470661,13.595129,14.7156925,15.84016,16.960724,17.686943,18.41316,19.13938,19.861694,20.587914,21.860748,23.137487,24.414227,25.687063,26.963802,27.717352,28.470901,29.228355,29.981905,30.739359,30.102942,29.466524,28.834011,28.197594,27.561176,25.73782,23.914463,22.087204,20.263847,18.436588,16.808453,15.18422,13.556085,11.927949,10.299813,9.944512,9.589212,9.2339115,8.878611,8.52331,8.78881,9.050405,9.311999,9.573594,9.839094,10.124115,10.409137,10.694158,10.979179,11.2642,11.49456,11.728825,11.959184,12.193448,12.423808,15.070992,17.718178,20.369267,23.01645,25.663635,23.01645,20.369267,17.718178,15.070992,12.423808,13.271063,14.114414,14.96167,15.80502,16.64837,15.4965725,14.344774,13.192975,12.041177,10.889378,11.318862,11.752251,12.185639,12.619028,13.048512,11.642927,10.2334385,8.827853,7.4183645,6.012779,6.153338,6.297801,6.4383593,6.5828223,6.7233806,8.519405,10.315431,12.111456,13.903577,15.699601,13.028991,10.354475,7.6838636,5.009348,2.338737,5.2358036,8.136774,11.037745,13.938716,16.835783,17.698656,18.56153,19.4244,20.287273,21.150146,17.429253,13.704452,9.983557,6.2587566,2.5378613,2.8385005,3.1391394,3.435874,3.736513,4.037152,5.196759,6.356367,7.5159745,8.675582,9.839094,8.601398,7.363703,6.126007,4.8883114,3.6506162,5.267039,6.883461,8.503788,10.120211,11.736633,10.77615,9.811763,8.85128,7.8868923,6.9264097,6.114294,5.3060827,4.493967,3.6857557,2.87364,3.1313305,3.3890212,3.6467118,3.9044023,4.1620927,3.8965936,3.6271896,3.3616903,3.0922866,2.8267872,2.697942,2.5690966,2.4441557,2.3153105,2.1864653,1.9561055,1.7218413,1.4914817,1.2572175,1.0268579,1.6749885,2.3231194,2.9751544,3.6232853,4.2753205,4.084005,3.8887846,3.697469,3.506153,3.310933,4.044961,4.7789884,5.5091114,6.2431393,6.9732623,7.191909,7.406651,7.621393,7.8361354,8.050878,7.7892823,7.523783,7.262188,7.000593,6.7389984,6.606249,6.473499,6.3407493,6.2079997,6.0752497,5.3412223,4.60329,3.8692627,3.135235,2.4012074,2.6081407,2.8189783,3.0298162,3.240654,3.4514916,3.1430438,2.8345962,2.5261483,2.2216048,1.9131571,1.6281357,1.3431144,1.0580931,0.77307165,0.48805028,0.8862993,1.2806439,1.678893,2.077142,2.475391,2.436347,2.3933985,2.3543546,2.3153105,2.2762666,2.2684577,2.260649,2.25284,2.2450314,2.2372224,3.2757936,4.318269,5.35684,6.3993154,7.437886,7.800996,8.164105,8.52331,8.886419,9.249529,8.218767,7.191909,6.1611466,5.1303844,4.0996222,4.1035266,4.1035266,4.1074314,4.1113358,4.1113358,3.8614538,3.6076677,3.3538816,3.1039999,2.8502135,2.5495746,2.2489357,1.9482968,1.6515622,1.3509232,1.4055848,1.4602464,1.5149081,1.5695697,1.6242313,2.6823244,3.7404175,4.7985106,5.8566036,6.910792,7.1333427,7.3519893,7.570636,7.793187,8.011833,7.426173,6.8366084,6.250948,5.661383,5.0757227,4.9156423,4.755562,4.5954814,4.435401,4.2753205,4.1894236,4.0996222,4.0137253,3.9239242,3.8380275,3.7052777,3.5725281,3.4397783,3.3070288,3.174279,3.0141985,2.8502135,2.6862288,2.5261483,2.3621633,2.1044729,1.8467822,1.5890918,1.3314011,1.0737107,0.98390937,0.8902037,0.79649806,0.7066968,0.61299115,0.6481308,0.6871748,0.7262188,0.76135844,0.80040246,0.6715572,0.5466163,0.41777104,0.28892577,0.1639849,0.28892577,0.41777104,0.5466163,0.6715572,0.80040246,0.6832704,0.5661383,0.44900626,0.3318742,0.21083772,0.28502136,0.359205,0.42948425,0.5036679,0.57394713,0.5309987,0.48414588,0.44119745,0.39434463,0.3513962,0.28892577,0.22645533,0.1639849,0.10151446,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.19912452,0.19912452,0.19912452,0.19912452,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08980125,0.1796025,0.26940376,0.359205,0.44900626,0.679366,0.9058213,1.1322767,1.358732,1.5890918,1.737459,1.8858263,2.0380979,2.1864653,2.338737,2.4324427,2.5261483,2.6237583,2.717464,2.8111696,3.049338,3.2836022,3.5178664,3.7521305,3.9863946,4.3026514,4.618908,4.93126,5.2475166,5.563773,5.4388323,5.3138914,5.1889505,5.0640097,4.939069,4.657952,4.376835,4.095718,3.8185053,3.5373883,4.3455997,5.153811,5.958118,6.7663293,7.57454,8.011833,8.445222,8.878611,9.315904,9.749292,9.370565,8.991838,8.609207,8.23048,7.8517528,6.754616,5.661383,4.564246,3.4710135,2.3738766,2.077142,1.7804074,1.4836729,1.1869383,0.8862993,0.80040246,0.7106012,0.62470436,0.5388075,0.44900626,0.37872702,0.30454338,0.23426414,0.16008049,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.03513962,0.05075723,0.07027924,0.08589685,0.25769055,0.42557985,0.59737355,0.76916724,0.93705654,1.1791295,1.4172981,1.6593709,1.8975395,2.135708,2.5690966,3.0024853,3.435874,3.8692627,4.298747,4.5564375,4.814128,5.0718184,5.3295093,5.5871997,5.64967,5.7121406,5.774611,5.8370814,5.899552,6.1299114,6.3602715,6.590631,6.8209906,7.0513506,7.601871,8.148487,8.699008,9.249529,9.80005,9.565785,9.335425,9.101162,8.870802,8.636538,8.331994,8.027451,7.7229075,7.4183645,7.113821,7.6643414,8.210958,8.761478,9.311999,9.86252,10.436467,11.014318,11.588266,12.162213,12.73616,13.524849,14.313539,15.098324,15.8870125,16.675701,18.627903,20.580105,22.532305,24.484507,26.436708,26.081408,25.722202,25.366901,25.007696,24.64849,25.042835,25.433277,25.827621,26.218061,26.612406,28.049225,29.482141,30.91896,32.351875,33.788696,34.788223,35.791656,36.795086,37.79852,38.798046,37.997643,37.193336,36.392933,35.588627,34.788223,33.59738,32.40654,31.215696,30.028757,28.837915,27.643167,26.448421,25.253674,24.058928,22.86418,20.162333,17.464392,14.762545,12.0606985,9.362757,9.140205,8.917655,8.695104,8.472553,8.250002,8.265619,8.285142,8.300759,8.320281,8.335898,7.6955767,7.0513506,6.4110284,5.7668023,5.12648,5.368553,5.6145306,5.860508,6.1064854,6.348558,6.844417,7.336372,7.8283267,8.320281,8.812236,8.402273,7.9923115,7.5823493,7.172387,6.7624245,6.5633,6.364176,6.1611466,5.9620223,5.7628975,5.5403466,5.3177958,5.095245,4.872694,4.650143,4.7672753,4.884407,5.001539,5.1186714,5.2358036,5.1460023,5.0522966,4.958591,4.8687897,4.775084,5.2943697,5.813655,6.336845,6.8561306,7.375416,8.261715,9.14411,10.03041,10.916709,11.799104,12.841579,13.884054,14.92653,15.969006,17.01148,17.776743,18.538101,19.29946,20.06082,20.826082,22.286327,23.750479,25.210726,26.674877,28.139027,29.103415,30.067802,31.032188,31.996576,32.960964,32.30893,31.652988,30.99705,30.34111,29.689075,27.436235,25.1873,22.938364,20.685524,18.436588,16.578093,14.723501,12.8650055,11.00651,9.151918,8.8083315,8.468649,8.128965,7.7892823,7.4495993,7.8751793,8.300759,8.726339,9.151918,9.573594,9.393991,9.2104845,9.026978,8.843472,8.663869,9.284669,9.909373,10.530173,11.150972,11.775677,14.391626,17.01148,19.62743,22.24338,24.863234,22.032541,19.20185,16.371159,13.544372,10.71368,11.510178,12.306676,13.103174,13.903577,14.700074,13.930907,13.16174,12.388668,11.619501,10.850334,11.908427,12.970425,14.028518,15.090515,16.148607,14.051944,11.955279,9.858616,7.758047,5.661383,6.278279,6.89127,7.5081654,8.121157,8.738052,10.670732,12.607315,14.543899,16.476578,18.41316,15.15689,11.904523,8.648251,5.3919797,2.135708,5.4895897,8.835662,12.189544,15.539521,18.885593,20.486399,22.087204,23.68801,25.288813,26.885714,21.884174,16.87873,11.873287,6.8678436,1.8623998,2.338737,2.8111696,3.2875066,3.7638438,4.2362766,4.806319,5.3724575,5.938596,6.5086384,7.0747766,6.114294,5.1499066,4.185519,3.2250361,2.260649,3.4905357,4.716518,5.9464045,7.172387,8.398369,8.113348,7.824422,7.5394006,7.250475,6.9615493,6.3329406,5.704332,5.0718184,4.4432096,3.8106966,4.1581883,4.50568,4.853172,5.2006636,5.548156,4.872694,4.193328,3.5178664,2.8385005,2.1630387,1.9561055,1.7491722,1.5383345,1.3314011,1.1244678,1.1517987,1.1791295,1.2064602,1.2337911,1.261122,2.1513257,3.0376248,3.9239242,4.814128,5.700427,5.434928,5.169429,4.903929,4.6384296,4.376835,5.3607445,6.3446536,7.328563,8.316377,9.300286,9.518932,9.741484,9.96013,10.178777,10.401327,10.112402,9.823476,9.538455,9.249529,8.960603,8.78881,8.617016,8.445222,8.273428,8.101635,7.1216297,6.141625,5.1616197,4.181615,3.2016098,3.193801,3.1859922,3.1781836,3.1703746,3.1625657,2.9634414,2.7682211,2.5690966,2.3738766,2.174752,1.8702087,1.5656652,1.261122,0.95657855,0.6481308,1.1791295,1.7101282,2.241127,2.7682211,3.2992198,3.1157131,2.9361105,2.7526035,2.5690966,2.3855898,2.4792955,2.5690966,2.6588979,2.7486992,2.8385005,4.1308575,5.4271193,6.7233806,8.015738,9.311999,9.550168,9.788337,10.0265045,10.260769,10.498938,9.2104845,7.918128,6.629675,5.3412223,4.0488653,4.1074314,4.165997,4.220659,4.279225,4.337791,4.2167544,4.095718,3.978586,3.8575494,3.736513,3.310933,2.8892577,2.463678,2.0380979,1.6125181,1.678893,1.7413634,1.8077383,1.8741131,1.9365835,3.2367494,4.533011,5.8292727,7.125534,8.4257,8.722435,9.019169,9.315904,9.616543,9.913278,9.050405,8.187531,7.3246584,6.461786,5.5989127,5.4583545,5.3138914,5.173333,5.02887,4.8883114,4.900025,4.911738,4.9234514,4.939069,4.950782,4.802415,4.6540475,4.50568,4.3612175,4.21285,3.8887846,3.5608149,3.2367494,2.912684,2.5886188,2.3270237,2.069333,1.8077383,1.5461433,1.2884527,1.1869383,1.0815194,0.98000497,0.8784905,0.77307165,0.7106012,0.6481308,0.58566034,0.5231899,0.46071947,0.39434463,0.3240654,0.25378615,0.1835069,0.113227665,0.1835069,0.25378615,0.3240654,0.39434463,0.46071947,0.39824903,0.3318742,0.26940376,0.20302892,0.13665408,0.1796025,0.22255093,0.26549935,0.30844778,0.3513962,0.3279698,0.30454338,0.28111696,0.26159495,0.23816854,0.19912452,0.1639849,0.12494087,0.08589685,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.63641757,0.8355421,1.038571,1.2376955,1.43682,1.6359446,1.8389735,2.0380979,2.2372224,2.436347,2.5261483,2.612045,2.7018464,2.787743,2.87364,3.076669,3.2757936,3.474918,3.6740425,3.873167,4.1620927,4.4510183,4.73604,5.024966,5.3138914,5.138193,4.9624953,4.786797,4.6110992,4.4393053,4.0996222,3.7638438,3.4241607,3.0883822,2.7486992,3.736513,4.7243266,5.7121406,6.699954,7.687768,8.1992445,8.710721,9.226103,9.737579,10.249056,9.698535,9.151918,8.601398,8.050878,7.5003567,6.2743745,5.0483923,3.8263142,2.6003318,1.3743496,1.2259823,1.0737107,0.92534333,0.77307165,0.62470436,0.5622339,0.4997635,0.43729305,0.37482262,0.31235218,0.24988174,0.18741131,0.12494087,0.062470436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.24988174,0.43729305,0.62470436,0.81211567,0.999527,1.2259823,1.4485333,1.6749885,1.901444,2.1239948,2.6745155,3.2250361,3.775557,4.3260775,4.8765984,5.1889505,5.5013027,5.813655,6.126007,6.4383593,6.426646,6.4110284,6.3993154,6.387602,6.375889,6.524256,6.676528,6.824895,6.9732623,7.125534,7.7619514,8.398369,9.0386915,9.675109,10.311526,10.151445,9.987461,9.823476,9.663396,9.499411,9.01136,8.52331,8.039165,7.551114,7.0630636,7.5120697,7.9610763,8.413987,8.862993,9.311999,9.964035,10.612165,11.2642,11.912332,12.564366,13.224211,13.887959,14.551707,15.211552,15.875299,17.437061,18.998821,20.564487,22.126247,23.68801,23.426414,23.160913,22.899319,22.637724,22.37613,22.07549,21.77485,21.474213,21.173573,20.876839,21.485926,22.098917,22.711908,23.3249,23.937891,24.937418,25.936945,26.936472,27.935999,28.93943,29.025326,29.111223,29.201025,29.28692,29.376722,28.93943,28.498232,28.06094,27.623646,27.186354,26.089216,24.988174,23.887133,22.78609,21.688955,18.725513,15.762072,12.798631,9.839094,6.8756523,7.1762915,7.47693,7.773665,8.074304,8.374943,8.574067,8.773191,8.976221,9.175345,9.37447,8.511597,7.648724,6.785851,5.9268827,5.0640097,5.376362,5.688714,6.001066,6.3134184,6.6257706,7.1762915,7.726812,8.273428,8.823949,9.37447,8.85128,8.324185,7.800996,7.2739015,6.7507114,6.575013,6.3993154,6.223617,6.0518236,5.8761253,5.6379566,5.3997884,5.1616197,4.9234514,4.689187,4.7009,4.7126136,4.7243266,4.73604,4.7516575,4.6735697,4.5993857,4.5252023,4.4510183,4.376835,5.138193,5.899552,6.66091,7.426173,8.187531,8.999647,9.811763,10.6238785,11.435994,12.24811,13.212498,14.176885,15.137367,16.101755,17.062239,17.86264,18.663042,19.463446,20.263847,21.06425,22.711908,24.36347,26.011127,27.66269,29.314253,30.489477,31.660797,32.83602,34.01125,35.186474,34.511013,33.839455,33.163994,32.488533,31.81307,29.138554,26.464039,23.785618,21.111103,18.436588,16.351637,14.262781,12.173926,10.088976,8.00012,7.676055,7.348085,7.0240197,6.699954,6.375889,6.9615493,7.551114,8.136774,8.726339,9.311999,8.663869,8.011833,7.363703,6.7116675,6.0635366,7.0747766,8.086017,9.101162,10.112402,11.123642,13.712261,16.300879,18.889498,21.474213,24.062832,21.048632,18.038338,15.024139,12.013845,8.999647,9.749292,10.498938,11.248583,11.998228,12.751778,12.361338,11.974802,11.588266,11.20173,10.81129,12.501896,14.188598,15.875299,17.562002,19.248703,16.46096,13.673217,10.885473,8.101635,5.3138914,6.3993154,7.4886436,8.574067,9.663396,10.748819,12.825961,14.899199,16.976341,19.049578,21.12672,17.288692,13.450665,9.612638,5.774611,1.9365835,5.7394714,9.538455,13.337439,17.136421,20.93931,23.274141,25.612879,27.951616,30.286448,32.625187,26.335194,20.049105,13.763018,7.473026,1.1869383,1.8389735,2.4871042,3.1391394,3.78727,4.4393053,4.4119744,4.388548,4.3612175,4.337791,4.3143644,3.6232853,2.9361105,2.2489357,1.5617609,0.8745861,1.7140326,2.5495746,3.3890212,4.224563,5.0640097,5.4505453,5.8370814,6.223617,6.6140575,7.000593,6.551587,6.098676,5.64967,5.2006636,4.7516575,5.1889505,5.6262436,6.0635366,6.5008297,6.9381227,5.8487945,4.7633705,3.6740425,2.5886188,1.4992905,1.2142692,0.92534333,0.63641757,0.3513962,0.062470436,0.3513962,0.63641757,0.92534333,1.2142692,1.4992905,2.6237583,3.7482262,4.8765984,6.001066,7.125534,6.785851,6.4500723,6.114294,5.774611,5.4388323,6.676528,7.914223,9.151918,10.38571,11.623405,11.849861,12.076316,12.298867,12.525322,12.751778,12.439425,12.123169,11.810817,11.498465,11.186112,10.975275,10.764437,10.549695,10.338858,10.124115,8.898132,7.676055,6.4500723,5.22409,3.998108,3.775557,3.5491016,3.3265507,3.1000953,2.87364,2.787743,2.7018464,2.612045,2.5261483,2.436347,2.1122816,1.7882162,1.4641509,1.1361811,0.81211567,1.475864,2.135708,2.7994564,3.4632049,4.123049,3.7989833,3.474918,3.1508527,2.8267872,2.4988174,2.6862288,2.87364,3.0610514,3.2484627,3.435874,4.985922,6.5359693,8.086017,9.636065,11.186112,11.29934,11.412568,11.525795,11.639023,11.748346,10.198298,8.648251,7.098203,5.548156,3.998108,4.1113358,4.224563,4.337791,4.4510183,4.564246,4.575959,4.5876727,4.5993857,4.6110992,4.6267166,4.0761957,3.5256753,2.9751544,2.4246337,1.8741131,1.9482968,2.0263848,2.1005683,2.174752,2.2489357,3.78727,5.3256044,6.8639393,8.398369,9.936704,10.311526,10.686349,11.061172,11.435994,11.810817,10.674636,9.538455,8.398369,7.262188,6.126007,6.001066,5.8761253,5.7511845,5.6262436,5.5013027,5.610626,5.7238536,5.8370814,5.950309,6.0635366,5.899552,5.735567,5.575486,5.4115014,5.251421,4.7633705,4.2753205,3.78727,3.2992198,2.8111696,2.5495746,2.2879796,2.0263848,1.7608855,1.4992905,1.3860629,1.2767396,1.1635119,1.0502841,0.93705654,0.77307165,0.61299115,0.44900626,0.28892577,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.19912452,0.19912452,0.19912452,0.19912452,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08199245,0.1639849,0.24597734,0.3318742,0.41386664,0.60127795,0.78868926,0.97610056,1.1635119,1.3509232,1.5851873,1.8194515,2.0537157,2.2918842,2.5261483,2.6354716,2.7447948,2.854118,2.9634414,3.076669,3.2367494,3.39683,3.5569105,3.7130866,3.873167,4.087909,4.298747,4.513489,4.7243266,4.939069,4.802415,4.6657605,4.533011,4.396357,4.263607,4.01763,3.7716527,3.5256753,3.2836022,3.0376248,3.9317331,4.8219366,5.716045,6.606249,7.5003567,8.105539,8.710721,9.315904,9.921086,10.526268,9.721962,8.913751,8.109444,7.3051367,6.5008297,5.4700675,4.4393053,3.408543,2.3816853,1.3509232,1.1986516,1.0463798,0.8941081,0.7418364,0.58566034,0.5231899,0.46071947,0.39824903,0.3357786,0.27330816,0.21864653,0.1639849,0.10932326,0.05466163,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.21083772,0.3709182,0.5309987,0.6910792,0.8511597,1.0502841,1.2494087,1.4485333,1.6515622,1.8506867,2.3894942,2.9283018,3.4710135,4.009821,4.548629,4.9781127,5.4036927,5.833177,6.2587566,6.688241,6.66091,6.6374836,6.6140575,6.5867267,6.5633,6.6335793,6.707763,6.7819467,6.852226,6.9264097,7.3715115,7.8205175,8.265619,8.714626,9.163632,9.105066,9.0465,8.991838,8.933272,8.874706,8.531119,8.191436,7.8478484,7.504261,7.1606736,7.535496,7.9064145,8.281238,8.652155,9.023073,9.554072,10.081166,10.608261,11.135355,11.66245,12.330102,12.997755,13.665408,14.33306,15.000713,16.33602,17.675228,19.010534,20.349745,21.688955,21.466404,21.243853,21.021301,20.79875,20.5762,20.556679,20.54106,20.521538,20.50592,20.486399,21.220427,21.95055,22.684578,23.418604,24.148727,24.82419,25.495747,26.167303,26.838861,27.514322,27.623646,27.736874,27.850101,27.96333,28.076557,28.197594,28.31863,28.443571,28.564608,28.685644,27.729065,26.768581,25.8081,24.847616,23.887133,21.20481,18.522484,15.84016,13.157836,10.475512,10.416945,10.358379,10.303718,10.2451515,10.186585,10.03041,9.874233,9.714153,9.557977,9.4018,8.741957,8.086017,7.426173,6.7702336,6.114294,6.446168,6.7819467,7.1177254,7.453504,7.7892823,8.226576,8.667773,9.108971,9.546264,9.987461,9.6243515,9.261242,8.898132,8.538928,8.175818,7.843944,7.5159745,7.1841,6.8561306,6.524256,6.329036,6.133816,5.938596,5.743376,5.548156,5.548156,5.5442514,5.5442514,5.5403466,5.5364423,5.5403466,5.5442514,5.5442514,5.548156,5.548156,6.2860875,7.0240197,7.7619514,8.499884,9.237816,10.010887,10.787864,11.560935,12.337912,13.110983,13.958238,14.809398,15.656653,16.503908,17.351164,18.089096,18.823124,19.561056,20.298986,21.036919,22.508879,23.976934,25.448895,26.916948,28.388908,29.536802,30.680794,31.828688,32.97658,34.124477,33.468536,32.8165,32.16056,31.504622,30.848682,28.466997,26.085312,23.703627,21.318037,18.936352,16.82407,14.707883,12.591698,10.479416,8.36323,7.871275,7.3832245,6.89127,6.4032197,5.911265,6.5086384,7.1060123,7.703386,8.300759,8.898132,8.433509,7.9649806,7.4964523,7.0318284,6.5633,7.2543793,7.941554,8.632633,9.323712,10.010887,12.064603,14.118319,16.168129,18.221846,20.27556,17.956347,15.633226,13.314012,10.994797,8.675582,9.253433,9.835189,10.413041,10.994797,11.576552,11.393045,11.209538,11.0260315,10.84643,10.662923,12.197352,13.731783,15.266212,16.800642,18.338978,16.093946,13.852819,11.611692,9.366661,7.125534,7.70729,8.289046,8.870802,9.456462,10.0382185,11.6702585,13.302299,14.934339,16.56638,18.19842,15.078801,11.955279,8.831758,5.708236,2.5886188,5.5832953,8.581876,11.580457,14.579038,17.573715,19.49468,21.415646,23.336613,25.253674,27.17464,22.21605,17.253553,12.294963,7.336372,2.3738766,2.8502135,3.3265507,3.7989833,4.2753205,4.7516575,4.8375545,4.9234514,5.0132523,5.099149,5.1889505,4.349504,3.513962,2.6745155,1.8389735,0.999527,2.0927596,3.1859922,4.279225,5.368553,6.461786,6.5008297,6.5359693,6.575013,6.6140575,6.649197,6.2353306,5.8214636,5.4036927,4.989826,4.575959,4.950782,5.3295093,5.708236,6.083059,6.461786,5.575486,4.6930914,3.8067923,2.9243972,2.0380979,1.7843118,1.53443,1.2806439,1.0268579,0.77697605,0.94876975,1.1205635,1.2923572,1.4641509,1.6359446,2.7994564,3.959064,5.1186714,6.278279,7.437886,7.0357327,6.6335793,6.2314262,5.8292727,5.423215,6.6843367,7.941554,9.198771,10.455989,11.713207,12.146595,12.576079,13.009468,13.442857,13.8762455,13.677121,13.481901,13.282777,13.083652,12.888432,12.751778,12.611219,12.4745655,12.337912,12.201257,10.77615,9.354948,7.9337454,6.5086384,5.087436,4.8883114,4.689187,4.4861584,4.2870336,4.087909,4.0918136,4.0918136,4.095718,4.095718,4.0996222,3.8614538,3.6232853,3.3890212,3.1508527,2.912684,3.5100577,4.1074314,4.704805,5.3021784,5.899552,5.477876,5.056201,4.6345253,4.2089458,3.78727,3.7599394,3.7326086,3.7052777,3.677947,3.6506162,5.0757227,6.504734,7.9337454,9.358852,10.787864,10.67854,10.569217,10.455989,10.346666,10.237343,9.175345,8.113348,7.0513506,5.989353,4.9234514,4.989826,5.056201,5.1186714,5.185046,5.251421,5.532538,5.813655,6.098676,6.379793,6.66091,6.3134184,5.9620223,5.6145306,5.263134,4.911738,4.572055,4.2323723,3.892689,3.5530062,3.213323,4.251894,5.2865605,6.3251314,7.363703,8.398369,8.710721,9.023073,9.339331,9.651682,9.964035,9.019169,8.078208,7.1333427,6.192382,5.251421,5.196759,5.1460023,5.0913405,5.040583,4.985922,5.099149,5.212377,5.3256044,5.4388323,5.548156,5.35684,5.165524,4.9742084,4.7789884,4.5876727,4.251894,3.912211,3.5764325,3.2367494,2.900971,2.5964274,2.2957885,1.9912452,1.6906061,1.3860629,1.3314011,1.2728351,1.2142692,1.1557031,1.1010414,0.9136301,0.7262188,0.5388075,0.3513962,0.1639849,0.15617609,0.15227169,0.14836729,0.14055848,0.13665408,0.13274968,0.12884527,0.12103647,0.11713207,0.113227665,0.12884527,0.14836729,0.1639849,0.1835069,0.19912452,0.19131571,0.1835069,0.1756981,0.1717937,0.1639849,0.15227169,0.14055848,0.13274968,0.12103647,0.113227665,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.14836729,0.14836729,0.14836729,0.14836729,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.078088045,0.15617609,0.23426414,0.30844778,0.38653582,0.5622339,0.737932,0.9136301,1.0893283,1.261122,1.53443,1.8038338,2.0732377,2.3426414,2.612045,2.7447948,2.8775444,3.0102942,3.1430438,3.2757936,3.39683,3.513962,3.6349986,3.7560349,3.873167,4.0137253,4.1503797,4.2870336,4.423688,4.564246,4.466636,4.3729305,4.279225,4.181615,4.087909,3.9356375,3.7833657,3.631094,3.4788225,3.3265507,4.123049,4.919547,5.716045,6.5164475,7.3129454,8.011833,8.706817,9.405705,10.100689,10.799577,9.741484,8.679486,7.621393,6.559396,5.5013027,4.6657605,3.8302186,2.9946766,2.1591344,1.3235924,1.1713207,1.0151446,0.8589685,0.7066968,0.5505207,0.48805028,0.42557985,0.3631094,0.30063897,0.23816854,0.19131571,0.14055848,0.093705654,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.1717937,0.30063897,0.43338865,0.5661383,0.698888,0.8745861,1.0502841,1.2259823,1.4016805,1.5734742,2.1044729,2.6354716,3.1664703,3.6935644,4.224563,4.7672753,5.309987,5.852699,6.395411,6.9381227,6.899079,6.8639393,6.824895,6.785851,6.7507114,6.746807,6.7389984,6.735094,6.7311897,6.7233806,6.9810715,7.238762,7.4964523,7.7541428,8.011833,8.058686,8.109444,8.156297,8.203149,8.250002,8.050878,7.8556576,7.656533,7.461313,7.262188,7.558923,7.8517528,8.148487,8.441318,8.738052,9.14411,9.546264,9.952321,10.358379,10.764437,11.435994,12.107552,12.779109,13.450665,14.126127,15.238882,16.351637,17.464392,18.573242,19.685997,19.506393,19.322887,19.13938,18.955873,18.77627,19.041769,19.303364,19.568865,19.834364,20.099863,20.951023,21.806087,22.657246,23.508406,24.36347,24.707058,25.050644,25.398136,25.741724,26.089216,26.22587,26.362524,26.499178,26.635832,26.77639,27.455757,28.139027,28.822298,29.505568,30.188839,29.368914,28.548988,27.729065,26.90914,26.089216,23.684105,21.282896,18.88169,16.476578,14.07537,13.661504,13.243732,12.829865,12.415999,11.998228,11.486752,10.971371,10.455989,9.940608,9.425227,8.972317,8.519405,8.066495,7.6135845,7.1606736,7.519879,7.8790836,8.234385,8.59359,8.94889,9.280765,9.608734,9.940608,10.268578,10.600452,10.401327,10.198298,9.999174,9.80005,9.600925,9.116779,8.628729,8.144583,7.660437,7.1762915,7.0240197,6.871748,6.715572,6.5633,6.4110284,6.395411,6.375889,6.3602715,6.3407493,6.3251314,6.4032197,6.4852123,6.5633,6.6452928,6.7233806,7.437886,8.148487,8.862993,9.573594,10.2881,11.0260315,11.763964,12.501896,13.235924,13.973856,14.707883,15.441911,16.172033,16.906061,17.636185,18.311647,18.987108,19.662569,20.338032,21.013493,22.301945,23.594303,24.882755,26.171207,27.463566,28.58413,29.700788,30.821352,31.941916,33.062477,32.42606,31.793547,31.15713,30.520712,29.888199,27.799343,25.706585,23.61773,21.528873,19.436115,17.296501,15.152986,13.009468,10.865952,8.726339,8.070399,7.4144597,6.75852,6.1064854,5.4505453,6.055728,6.6648145,7.2739015,7.8790836,8.488171,8.203149,7.918128,7.633106,7.348085,7.0630636,7.4300776,7.7970915,8.164105,8.531119,8.898132,10.416945,11.935758,13.45457,14.969479,16.48829,14.860155,13.232019,11.603884,9.975748,8.351517,8.761478,9.171441,9.581403,9.991365,10.401327,10.42085,10.444276,10.467703,10.491129,10.510651,11.896713,13.2788725,14.661031,16.043188,17.425346,15.726933,14.028518,12.334006,10.6355915,8.937177,9.0152645,9.093353,9.171441,9.245625,9.323712,10.514555,11.705398,12.89624,14.0831785,15.274021,12.86891,10.459893,8.050878,5.645766,3.2367494,5.4310236,7.629202,9.823476,12.01775,14.212025,15.7152195,17.218414,18.72161,20.2209,21.724094,18.093,14.461906,10.826907,7.195813,3.5608149,3.8614538,4.1620927,4.462732,4.7633705,5.0640097,5.263134,5.462259,5.661383,5.8644123,6.0635366,5.0757227,4.087909,3.1000953,2.1122816,1.1244678,2.4714866,3.8185053,5.169429,6.5164475,7.8634663,7.551114,7.238762,6.9264097,6.6140575,6.3017054,5.919074,5.5403466,5.1616197,4.7789884,4.4002614,4.716518,5.036679,5.3529353,5.6691923,5.989353,5.3060827,4.6228123,3.9395418,3.2562714,2.5769055,2.358259,2.1396124,1.9209659,1.7062237,1.4875772,1.5461433,1.6008049,1.6593709,1.717937,1.7765031,2.97125,4.165997,5.3607445,6.5554914,7.7502384,7.28171,6.813182,6.348558,5.8800297,5.4115014,6.688241,7.968885,9.245625,10.522364,11.799104,12.439425,13.079747,13.72007,14.360392,15.000713,14.918721,14.836729,14.750832,14.668839,14.586847,14.524376,14.461906,14.399435,14.336966,14.274494,12.654168,11.033841,9.413514,7.793187,6.1767645,6.001066,5.825368,5.64967,5.473972,5.298274,5.3919797,5.4856853,5.579391,5.6691923,5.7628975,5.610626,5.462259,5.3138914,5.1616197,5.0132523,5.5442514,6.0791545,6.610153,7.141152,7.676055,7.1567693,6.6335793,6.114294,5.5950084,5.0757227,4.83365,4.591577,4.3455997,4.1035266,3.8614538,5.169429,6.473499,7.7775693,9.081639,10.38571,10.053836,9.721962,9.390087,9.058213,8.726339,8.148487,7.57454,7.000593,6.426646,5.8487945,5.8683167,5.883934,5.903456,5.919074,5.938596,6.4891167,7.043542,7.5940623,8.148487,8.699008,8.550641,8.398369,8.250002,8.101635,7.9493628,7.195813,6.4383593,5.6848097,4.93126,4.173806,4.7126136,5.251421,5.786324,6.3251314,6.8639393,7.113821,7.363703,7.6135845,7.8634663,8.113348,7.363703,6.617962,5.8683167,5.1225758,4.376835,4.396357,4.415879,4.435401,4.454923,4.474445,4.5876727,4.7009,4.814128,4.9234514,5.036679,4.814128,4.591577,4.369026,4.1464753,3.9239242,3.736513,3.5491016,3.3616903,3.174279,2.9868677,2.6432803,2.3035975,1.9600099,1.6164225,1.2767396,1.2728351,1.2689307,1.2689307,1.2650263,1.261122,1.0502841,0.8355421,0.62470436,0.41386664,0.19912452,0.20302892,0.20693332,0.20693332,0.21083772,0.21083772,0.19131571,0.1678893,0.14446288,0.12103647,0.10151446,0.14836729,0.19522011,0.24207294,0.28892577,0.3357786,0.30844778,0.28111696,0.25378615,0.22645533,0.19912452,0.1796025,0.16008049,0.14055848,0.12103647,0.10151446,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14446288,0.21864653,0.28892577,0.3631094,0.5231899,0.6871748,0.8511597,1.0112402,1.175225,1.4797685,1.7843118,2.0888553,2.3933985,2.7018464,2.854118,3.0102942,3.1664703,3.3187418,3.474918,3.5569105,3.6349986,3.7130866,3.795079,3.873167,3.9356375,3.998108,4.0605783,4.123049,4.1894236,4.1308575,4.0761957,4.0215344,3.9668727,3.912211,3.853645,3.7911747,3.7326086,3.6740425,3.611572,4.3143644,5.017157,5.7199492,6.422742,7.125534,7.914223,8.706817,9.495506,10.284196,11.076789,9.761005,8.445222,7.1294384,5.813655,4.5017757,3.8614538,3.2211318,2.5808098,1.9404879,1.3001659,1.1439898,0.98390937,0.8277333,0.6715572,0.5114767,0.44900626,0.38653582,0.3240654,0.26159495,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.12884527,0.23426414,0.339683,0.44510186,0.5505207,0.698888,0.8511597,0.999527,1.1517987,1.3001659,1.8194515,2.338737,2.8619268,3.3812122,3.900498,4.5564375,5.2162814,5.872221,6.5281606,7.1880045,7.137247,7.08649,7.0357327,6.98888,6.9381227,6.8561306,6.774138,6.688241,6.606249,6.524256,6.590631,6.66091,6.727285,6.79366,6.8639393,7.016211,7.168483,7.320754,7.473026,7.6252975,7.570636,7.519879,7.4691215,7.4144597,7.363703,7.578445,7.7970915,8.015738,8.234385,8.449126,8.734148,9.0152645,9.296382,9.581403,9.86252,10.541886,11.217348,11.896713,12.572175,13.251541,14.13784,15.024139,15.914344,16.800642,17.686943,17.546383,17.40192,17.261362,17.1169,16.976341,17.522957,18.069574,18.61619,19.16671,19.713327,20.685524,21.657719,22.629915,23.602112,24.574308,24.59383,24.609447,24.62897,24.644587,24.664108,24.82419,24.988174,25.148254,25.31224,25.476225,26.717825,27.959425,29.201025,30.44653,31.68813,31.008762,30.329397,29.646126,28.96676,28.287394,26.163399,24.043308,21.919313,19.799223,17.675228,16.902157,16.129086,15.356014,14.586847,13.813775,12.939189,12.068507,11.193921,10.323239,9.448653,9.202676,8.956698,8.706817,8.460839,8.210958,8.59359,8.972317,9.351044,9.733675,10.112402,10.331048,10.553599,10.772245,10.990892,11.213444,11.174399,11.139259,11.100216,11.061172,11.0260315,10.38571,9.745388,9.105066,8.464745,7.824422,7.715099,7.605776,7.4964523,7.3832245,7.2739015,7.2426662,7.211431,7.1762915,7.1450562,7.113821,7.269997,7.426173,7.5862536,7.7424297,7.898606,8.58578,9.276859,9.964035,10.651209,11.338385,12.037272,12.73616,13.438952,14.13784,14.836729,15.453624,16.074425,16.69132,17.308216,17.92511,18.538101,19.151093,19.764084,20.37317,20.986162,22.098917,23.207767,24.316618,25.429373,26.538221,27.631454,28.720783,29.814016,30.907248,32.00048,31.383585,30.770594,30.153698,29.540707,28.923813,27.127787,25.331762,23.531832,21.735807,19.935879,17.768934,15.598087,13.427239,11.256392,9.089449,8.265619,7.445695,6.6257706,5.805846,4.985922,5.606722,6.223617,6.8405128,7.4574084,8.074304,7.9727893,7.871275,7.7658563,7.6643414,7.562827,7.605776,7.6526284,7.6955767,7.7424297,7.7892823,8.769287,9.753197,10.733202,11.717112,12.70102,11.763964,10.8308115,9.893755,8.960603,8.023546,8.265619,8.503788,8.745861,8.98403,9.226103,9.452558,9.679013,9.909373,10.135828,10.362284,11.592171,12.822057,14.051944,15.281831,16.511717,15.359919,14.208119,13.056321,11.900618,10.748819,10.323239,9.893755,9.468176,9.0386915,8.6131115,9.358852,10.108498,10.8542385,11.603884,12.349625,10.6590185,8.964508,7.2739015,5.579391,3.8887846,5.278752,6.6726236,8.066495,9.456462,10.850334,11.935758,13.021181,14.106606,15.188125,16.273548,13.969952,11.666354,9.358852,7.055255,4.7516575,4.8765984,5.001539,5.12648,5.251421,5.376362,5.688714,6.001066,6.3134184,6.6257706,6.9381227,5.7980375,4.661856,3.5256753,2.3855898,1.2494087,2.854118,4.454923,6.055728,7.660437,9.261242,8.601398,7.9376497,7.2739015,6.6140575,5.950309,5.606722,5.2592297,4.9156423,4.5681505,4.224563,4.482254,4.7399445,4.997635,5.2553253,5.5130157,5.0327744,4.552533,4.0722914,3.59205,3.1118085,2.9283018,2.7486992,2.5651922,2.3816853,2.1981785,2.1435168,2.084951,2.0263848,1.9717231,1.9131571,3.1430438,4.3729305,5.602817,6.832704,8.062591,7.531592,6.996689,6.46569,5.930787,5.3997884,6.6960497,7.996216,9.292478,10.588739,11.888905,12.73616,13.583415,14.430671,15.277926,16.125181,16.156416,16.191557,16.222792,16.254026,16.289165,16.300879,16.312593,16.324306,16.33602,16.351637,14.532186,12.716639,10.897186,9.081639,7.262188,7.113821,6.9615493,6.813182,6.66091,6.5125427,6.6960497,6.8756523,7.0591593,7.2426662,7.426173,7.363703,7.3012323,7.238762,7.1762915,7.113821,7.578445,8.046973,8.515501,8.98403,9.448653,8.831758,8.214863,7.5979667,6.9810715,6.364176,5.903456,5.446641,4.989826,4.533011,4.0761957,5.2592297,6.4383593,7.621393,8.804427,9.987461,9.433036,8.878611,8.324185,7.7658563,7.211431,7.125534,7.0357327,6.949836,6.8639393,6.774138,6.746807,6.715572,6.6843367,6.6531014,6.6257706,7.445695,8.269524,9.093353,9.913278,10.737106,10.787864,10.838621,10.889378,10.936231,10.986988,9.815667,8.648251,7.47693,6.309514,5.138193,5.173333,5.212377,5.251421,5.2865605,5.3256044,5.5130157,5.700427,5.8878384,6.0752497,6.262661,5.708236,5.1577153,4.60329,4.0527697,3.4983444,3.59205,3.6857557,3.775557,3.8692627,3.9629683,4.0761957,4.1894236,4.298747,4.4119744,4.5252023,4.271416,4.0215344,3.767748,3.513962,3.2640803,3.2250361,3.1859922,3.1508527,3.1118085,3.076669,2.6940374,2.3114061,1.9287747,1.5461433,1.1635119,1.2142692,1.2689307,1.319688,1.3743496,1.4251068,1.1869383,0.94876975,0.7106012,0.47633708,0.23816854,0.24597734,0.25769055,0.26940376,0.27721256,0.28892577,0.24597734,0.20693332,0.1678893,0.12884527,0.08589685,0.1639849,0.24207294,0.32016098,0.39824903,0.47633708,0.42557985,0.37872702,0.3318742,0.28502136,0.23816854,0.20693332,0.1756981,0.14836729,0.11713207,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06637484,0.13665408,0.20302892,0.26940376,0.3357786,0.48805028,0.63641757,0.78868926,0.93705654,1.0893283,1.4290112,1.7686942,2.1083772,2.4480603,2.787743,2.9634414,3.1430438,3.3187418,3.4983444,3.6740425,3.7130866,3.7560349,3.795079,3.8341231,3.873167,3.8614538,3.8497405,3.8380275,3.8263142,3.8106966,3.7989833,3.7833657,3.767748,3.7521305,3.736513,3.7716527,3.802888,3.8341231,3.8692627,3.900498,4.50568,5.114767,5.7238536,6.329036,6.9381227,7.8205175,8.702912,9.585307,10.467703,11.350098,9.780528,8.210958,6.6413884,5.0718184,3.4983444,3.0532427,2.6081407,2.1630387,1.7218413,1.2767396,1.116659,0.95657855,0.79649806,0.63641757,0.47633708,0.41386664,0.3513962,0.28892577,0.22645533,0.1639849,0.12884527,0.09761006,0.06637484,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.08980125,0.1678893,0.24597734,0.3240654,0.39824903,0.5231899,0.6481308,0.77307165,0.9019169,1.0268579,1.53443,2.0459068,2.5534792,3.0649557,3.5764325,4.3455997,5.1186714,5.891743,6.6648145,7.437886,7.375416,7.3129454,7.250475,7.1880045,7.125534,6.9654536,6.805373,6.6452928,6.4852123,6.3251314,6.2040954,6.0791545,5.958118,5.833177,5.7121406,5.969831,6.2275214,6.4852123,6.7429028,7.000593,7.094299,7.1841,7.277806,7.3715115,7.461313,7.601871,7.7424297,7.882988,8.023546,8.164105,8.324185,8.484266,8.644346,8.804427,8.960603,9.643873,10.327144,11.010414,11.693685,12.373051,13.036799,13.700547,14.364296,15.024139,15.687888,15.586374,15.480955,15.37944,15.277926,15.176412,16.004145,16.835783,17.663515,18.495153,19.326792,20.416119,21.509352,22.602585,23.695818,24.78905,24.476698,24.16825,23.855898,23.54745,23.239002,23.426414,23.613825,23.801235,23.988647,24.17606,25.975988,27.779821,29.583656,31.383585,33.18742,32.648613,32.1059,31.567093,31.028284,30.489477,28.646599,26.803722,24.960844,23.117966,21.275087,20.146715,19.014439,17.886066,16.75379,15.625418,14.395531,13.165645,11.935758,10.705871,9.475985,9.433036,9.390087,9.347139,9.304191,9.261242,9.663396,10.069453,10.471607,10.87376,11.275913,11.385237,11.49456,11.603884,11.713207,11.826434,11.951375,12.076316,12.201257,12.326198,12.4511385,11.654641,10.858143,10.065549,9.269051,8.476458,8.406178,8.339804,8.273428,8.203149,8.136774,8.089922,8.043069,7.996216,7.9493628,7.898606,8.136774,8.371038,8.605303,8.839567,9.073831,9.737579,10.401327,11.061172,11.72492,12.388668,13.048512,13.712261,14.376009,15.035853,15.699601,16.20327,16.706938,17.206701,17.71037,18.214037,18.760653,19.311174,19.861694,20.412214,20.962736,21.891983,22.821232,23.754383,24.683632,25.612879,26.678782,27.740778,28.80668,29.872581,30.938484,30.34111,29.74764,29.154171,28.556799,27.96333,26.45623,24.953035,23.445936,21.942741,20.435642,18.241367,16.043188,13.845011,11.6468315,9.448653,8.464745,7.480835,6.493021,5.5091114,4.5252023,5.153811,5.7785153,6.407124,7.0357327,7.6643414,7.7424297,7.824422,7.90251,7.9805984,8.062591,7.785378,7.5081654,7.230953,6.9537406,6.676528,7.1216297,7.570636,8.015738,8.464745,8.913751,8.671678,8.4257,8.183627,7.941554,7.699481,7.7697606,7.8400397,7.910319,7.9805984,8.050878,8.484266,8.913751,9.347139,9.780528,10.213917,11.291532,12.369146,13.446761,14.524376,15.598087,14.992905,14.383818,13.778636,13.169549,12.564366,11.631214,10.698062,9.76491,8.831758,7.898606,8.203149,8.511597,8.81614,9.120684,9.425227,8.449126,7.4691215,6.493021,5.5169206,4.5369153,5.12648,5.716045,6.3056097,6.899079,7.4886436,8.156297,8.823949,9.491602,10.159255,10.823003,9.846903,8.870802,7.890797,6.914696,5.938596,5.8878384,5.8370814,5.786324,5.735567,5.688714,6.114294,6.5359693,6.9615493,7.387129,7.812709,6.524256,5.2358036,3.951255,2.6628022,1.3743496,3.232845,5.0913405,6.9459314,8.804427,10.662923,9.651682,8.636538,7.6252975,6.6140575,5.5989127,5.290465,4.9781127,4.6696653,4.3612175,4.0488653,4.2479897,4.4432096,4.6423345,4.841459,5.036679,4.759466,4.482254,4.2050414,3.9278288,3.6506162,3.5022488,3.3538816,3.2094188,3.0610514,2.912684,2.7408905,2.5690966,2.3933985,2.2216048,2.0498111,3.3148375,4.579864,5.84489,7.1099167,8.374943,7.7775693,7.180196,6.5828223,5.985449,5.388075,6.703859,8.023546,9.339331,10.6590185,11.974802,13.028991,14.0831785,15.141272,16.195461,17.24965,17.398016,17.546383,17.690847,17.839214,17.987581,18.073479,18.163279,18.249176,18.338978,18.424873,16.410202,14.395531,12.380859,10.366188,8.351517,8.226576,8.101635,7.9766936,7.8517528,7.726812,7.996216,8.269524,8.542832,8.81614,9.089449,9.112875,9.136301,9.163632,9.187058,9.21439,9.616543,10.018696,10.42085,10.823003,11.225157,10.510651,9.796145,9.081639,8.36323,7.648724,6.9771667,6.3056097,5.6340523,4.958591,4.2870336,5.349031,6.407124,7.4691215,8.527214,9.589212,8.8083315,8.031356,7.2543793,6.477403,5.700427,6.098676,6.5008297,6.899079,7.3012323,7.699481,7.621393,7.5433054,7.4691215,7.3910336,7.3129454,8.406178,9.499411,10.588739,11.681972,12.775204,13.025085,13.274967,13.524849,13.774731,14.024612,12.439425,10.8542385,9.269051,7.6838636,6.098676,5.6379566,5.173333,4.7126136,4.251894,3.78727,3.912211,4.037152,4.1620927,4.2870336,4.4119744,4.056674,3.697469,3.338264,2.9829633,2.6237583,2.7916477,2.9556324,3.1196175,3.2836022,3.4514916,3.5608149,3.6740425,3.78727,3.900498,4.0137253,3.7287042,3.4475873,3.1664703,2.8814487,2.6003318,2.7135596,2.8267872,2.9361105,3.049338,3.1625657,2.7408905,2.3192148,1.893635,1.4719596,1.0502841,1.1557031,1.2650263,1.3743496,1.4797685,1.5890918,1.3235924,1.0619974,0.80040246,0.5388075,0.27330816,0.29283017,0.30844778,0.3279698,0.3435874,0.3631094,0.30454338,0.24597734,0.19131571,0.13274968,0.07418364,0.1835069,0.28892577,0.39824903,0.5036679,0.61299115,0.5466163,0.47633708,0.40996224,0.3435874,0.27330816,0.23426414,0.19522011,0.15617609,0.113227665,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.44900626,0.58566034,0.7262188,0.8628729,0.999527,1.3743496,1.7491722,2.1239948,2.4988174,2.87364,3.076669,3.2757936,3.474918,3.6740425,3.873167,3.873167,3.873167,3.873167,3.873167,3.873167,3.78727,3.7013733,3.611572,3.5256753,3.435874,3.4632049,3.4866312,3.513962,3.5373883,3.5608149,3.6857557,3.8106966,3.9356375,4.0605783,4.1894236,4.7009,5.212377,5.7238536,6.239235,6.7507114,7.726812,8.699008,9.675109,10.651209,11.623405,9.80005,7.9766936,6.1494336,4.3260775,2.4988174,2.2489357,1.999054,1.7491722,1.4992905,1.2494087,1.0893283,0.92534333,0.76135844,0.60127795,0.43729305,0.37482262,0.31235218,0.24988174,0.18741131,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.3513962,0.44900626,0.5505207,0.6481308,0.74964523,1.2494087,1.7491722,2.2489357,2.7486992,3.2484627,4.138666,5.024966,5.911265,6.801469,7.687768,7.6135845,7.5394006,7.461313,7.387129,7.3129454,7.0747766,6.8366084,6.5984397,6.364176,6.126007,5.813655,5.5013027,5.1889505,4.8765984,4.564246,4.9234514,5.2865605,5.64967,6.012779,6.375889,6.6140575,6.8483214,7.08649,7.3246584,7.562827,7.6252975,7.687768,7.7502384,7.812709,7.8751793,7.914223,7.9493628,7.988407,8.023546,8.062591,8.749765,9.43694,10.124115,10.81129,11.498465,11.935758,12.373051,12.814248,13.251541,13.688834,13.626364,13.563893,13.501423,13.438952,13.376482,14.489237,15.598087,16.710842,17.823597,18.936352,20.15062,21.360985,22.575254,23.785618,24.999887,24.36347,23.723148,23.086731,22.450314,21.813896,22.024733,22.23557,22.450314,22.66115,22.875893,25.238056,27.60022,29.962383,32.324547,34.68671,34.28846,33.886307,33.48806,33.085903,32.687656,31.125895,29.564135,27.998468,26.436708,24.874947,23.38737,21.899792,20.412214,18.924637,17.437061,15.851873,14.262781,12.67369,11.088503,9.499411,9.663396,9.823476,9.987461,10.151445,10.311526,10.737106,11.162686,11.588266,12.013845,12.439425,12.439425,12.439425,12.439425,12.439425,12.439425,12.724447,13.013372,13.298394,13.58732,13.8762455,12.923572,11.974802,11.0260315,10.073358,9.124588,9.101162,9.073831,9.050405,9.023073,8.999647,8.937177,8.874706,8.812236,8.749765,8.687295,8.999647,9.311999,9.6243515,9.936704,10.249056,10.889378,11.525795,12.162213,12.798631,13.438952,14.063657,14.688361,15.313066,15.93777,16.562475,16.94901,17.335546,17.725986,18.112522,18.499058,18.987108,19.475159,19.96321,20.45126,20.93931,21.688955,22.4386,23.188246,23.937891,24.687536,25.726107,26.760773,27.799343,28.837915,29.876486,29.298634,28.724688,28.15074,27.576794,26.998941,25.788576,24.574308,23.363943,22.149673,20.93931,18.7138,16.48829,14.262781,12.037272,9.811763,8.663869,7.5120697,6.364176,5.212377,4.0605783,4.7009,5.337318,5.9737353,6.6140575,7.250475,7.5120697,7.773665,8.039165,8.300759,8.562354,7.9610763,7.363703,6.7624245,6.1611466,5.563773,5.473972,5.388075,5.298274,5.212377,5.12648,5.575486,6.0244927,6.473499,6.9264097,7.375416,7.2739015,7.1762915,7.0747766,6.9732623,6.8756523,7.5120697,8.148487,8.78881,9.425227,10.061645,10.986988,11.912332,12.837675,13.763018,14.688361,14.625891,14.56342,14.50095,14.438479,14.376009,12.939189,11.498465,10.061645,8.624825,7.1880045,7.0513506,6.910792,6.774138,6.6374836,6.5008297,6.239235,5.9737353,5.7121406,5.4505453,5.1889505,4.9742084,4.7633705,4.548629,4.337791,4.123049,4.376835,4.6267166,4.8765984,5.12648,5.376362,5.7238536,6.0752497,6.426646,6.774138,7.125534,6.899079,6.676528,6.4500723,6.223617,6.001066,6.5359693,7.0747766,7.6135845,8.148487,8.687295,7.250475,5.813655,4.376835,2.9361105,1.4992905,3.611572,5.7238536,7.8361354,9.948417,12.0606985,10.698062,9.339331,7.9766936,6.6140575,5.251421,4.9742084,4.7009,4.423688,4.1503797,3.873167,4.0137253,4.1503797,4.2870336,4.423688,4.564246,4.4861584,4.4119744,4.337791,4.263607,4.1894236,4.0761957,3.9629683,3.8497405,3.736513,3.6232853,3.338264,3.049338,2.7643168,2.475391,2.1864653,3.4866312,4.786797,6.086963,7.387129,8.687295,8.023546,7.363703,6.699954,6.036206,5.376362,6.7116675,8.050878,9.386183,10.725393,12.0606985,13.325725,14.586847,15.851873,17.112995,18.374117,18.635712,18.90121,19.162806,19.4244,19.685997,19.849981,20.013966,20.174046,20.338032,20.498112,18.28822,16.074425,13.860628,11.650736,9.43694,9.339331,9.237816,9.136301,9.0386915,8.937177,9.300286,9.663396,10.0265045,10.38571,10.748819,10.862047,10.975275,11.088503,11.20173,11.311053,11.650736,11.986515,12.326198,12.661977,13.001659,12.185639,11.373524,10.561408,9.749292,8.937177,8.050878,7.1606736,6.2743745,5.388075,4.5017757,5.4388323,6.375889,7.3129454,8.250002,9.187058,8.187531,7.1880045,6.1884775,5.1889505,4.1894236,5.0757227,5.9620223,6.8483214,7.7385254,8.624825,8.499884,8.374943,8.250002,8.125061,8.00012,9.362757,10.725393,12.08803,13.450665,14.813302,15.262308,15.711315,16.164225,16.613232,17.062239,15.063184,13.06413,11.061172,9.062118,7.0630636,6.098676,5.138193,4.173806,3.213323,2.2489357,2.3114061,2.3738766,2.436347,2.4988174,2.5612879,2.4012074,2.2372224,2.0732377,1.9131571,1.7491722,1.9873407,2.2255092,2.463678,2.7018464,2.9361105,3.049338,3.1625657,3.2757936,3.3890212,3.4983444,3.1859922,2.87364,2.5612879,2.2489357,1.9365835,2.1981785,2.463678,2.7252727,2.9868677,3.2484627,2.787743,2.3231194,1.8623998,1.4016805,0.93705654,1.1010414,1.261122,1.4251068,1.5890918,1.7491722,1.4641509,1.175225,0.8862993,0.60127795,0.31235218,0.3357786,0.3631094,0.38653582,0.41386664,0.43729305,0.3631094,0.28892577,0.21083772,0.13665408,0.062470436,0.19912452,0.3357786,0.47633708,0.61299115,0.74964523,0.6637484,0.57394713,0.48805028,0.39824903,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10541886,0.15617609,0.21083772,0.26159495,0.39044023,0.5192855,0.6442264,0.77307165,0.9019169,1.2767396,1.6515622,2.0263848,2.4012074,2.77603,2.9556324,3.1391394,3.3226464,3.506153,3.6857557,3.6935644,3.697469,3.7013733,3.7091823,3.7130866,3.5959544,3.4827268,3.3655949,3.252367,3.1391394,3.154757,3.174279,3.1898966,3.2094188,3.2250361,3.4788225,3.7287042,3.9824903,4.2362766,4.4861584,4.860981,5.2318993,5.606722,5.9776397,6.348558,7.28171,8.214863,9.148014,10.081166,11.014318,9.405705,7.7970915,6.1884775,4.5837684,2.9751544,2.6940374,2.416825,2.135708,1.8545911,1.5734742,1.3314011,1.0854238,0.8394465,0.59346914,0.3513962,0.30063897,0.24988174,0.19912452,0.14836729,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.07418364,0.12103647,0.1678893,0.21474212,0.26159495,0.3513962,0.44119745,0.5309987,0.62079996,0.7106012,1.2806439,1.8467822,2.416825,2.9829633,3.5491016,4.169902,4.7907014,5.4115014,6.028397,6.649197,6.5867267,6.524256,6.461786,6.3993154,6.336845,6.1767645,6.016684,5.8566036,5.6965227,5.5364423,5.298274,5.0640097,4.825841,4.5876727,4.349504,4.7009,5.056201,5.407597,5.758993,6.114294,6.2353306,6.356367,6.481308,6.602344,6.7233806,6.7311897,6.735094,6.7389984,6.746807,6.7507114,6.774138,6.801469,6.824895,6.8483214,6.8756523,7.3910336,7.910319,8.4257,8.944985,9.464272,9.999174,10.537982,11.076789,11.611692,12.150499,12.2559185,12.365242,12.470661,12.579984,12.689307,13.626364,14.56342,15.500477,16.437534,17.37459,18.506866,19.639143,20.77142,21.903696,23.035973,22.813423,22.586967,22.360512,22.13796,21.911505,22.46593,23.01645,23.570877,24.121397,24.675823,26.874,29.076084,31.274261,33.476345,35.674522,35.63548,35.596436,35.553486,35.514442,35.4754,34.17133,32.863354,31.559284,30.255213,28.951143,27.34253,25.733915,24.129206,22.520592,20.911978,19.678188,18.444397,17.206701,15.97291,14.739119,14.633699,14.528281,14.422862,14.317443,14.212025,14.750832,15.293544,15.832351,16.371159,16.91387,16.343828,15.77769,15.211552,14.641508,14.07537,13.973856,13.868437,13.766922,13.665408,13.563893,12.665881,11.771772,10.877665,9.983557,9.089449,8.995743,8.905942,8.81614,8.726339,8.636538,8.601398,8.562354,8.52331,8.488171,8.449126,8.781001,9.108971,9.440845,9.768814,10.100689,10.81129,11.525795,12.236397,12.950902,13.661504,14.348679,15.031949,15.719124,16.402393,17.085665,17.288692,17.491722,17.694752,17.89778,18.10081,18.631807,19.158901,19.689901,20.2209,20.751898,21.306324,21.864653,22.422981,22.981312,23.535736,24.507933,25.476225,26.448421,27.416712,28.388908,28.158548,27.92819,27.69783,27.46747,27.23711,26.112642,24.988174,23.863707,22.739239,21.610867,19.381453,17.148134,14.914817,12.681499,10.44818,9.288573,8.128965,6.969358,5.8097506,4.650143,5.22409,5.794133,6.36808,6.9381227,7.5120697,7.715099,7.918128,8.121157,8.324185,8.52331,7.910319,7.2934237,6.6804323,6.0635366,5.4505453,5.3841705,5.3217,5.2553253,5.1889505,5.12648,5.55206,5.9815445,6.407124,6.8366084,7.262188,7.2192397,7.1762915,7.1333427,7.094299,7.0513506,7.5276875,8.0040245,8.484266,8.960603,9.43694,10.38571,11.330575,12.2793455,13.228115,14.176885,14.376009,14.579038,14.782067,14.985096,15.188125,13.645885,12.107552,10.569217,9.026978,7.4886436,7.480835,7.47693,7.473026,7.4691215,7.461313,7.531592,7.601871,7.6721506,7.7424297,7.812709,7.289519,6.7624245,6.239235,5.7121406,5.1889505,5.2045684,5.22409,5.239708,5.2592297,5.2748475,5.4973984,5.7199492,5.9425,6.165051,6.387602,6.114294,5.840986,5.571582,5.298274,5.024966,5.423215,5.8214636,6.2158084,6.6140575,7.012306,5.989353,4.9663997,3.9434462,2.9243972,1.901444,3.541293,5.185046,6.8287997,8.468649,10.112402,9.14411,8.171914,7.2036223,6.2314262,5.263134,5.0483923,4.8375545,4.6267166,4.4119744,4.2011366,4.365122,4.5291066,4.6930914,4.860981,5.024966,5.0640097,5.1069584,5.1460023,5.185046,5.22409,5.0796275,4.9351645,4.7907014,4.646239,4.5017757,4.267512,4.0332475,3.802888,3.5686235,3.338264,4.396357,5.45445,6.5086384,7.5667315,8.624825,8.101635,7.57454,7.0513506,6.524256,6.001066,7.195813,8.39056,9.585307,10.780055,11.974802,12.939189,13.899672,14.864059,15.824542,16.788929,17.1169,17.448774,17.776743,18.108618,18.436588,18.538101,18.64352,18.745035,18.84655,18.948065,17.019289,15.090515,13.16174,11.229061,9.300286,9.261242,9.218294,9.17925,9.140205,9.101162,9.573594,10.049932,10.526268,10.998701,11.475039,11.45942,11.443803,11.428185,11.416472,11.400854,11.740538,12.08022,12.419904,12.759586,13.09927,12.31058,11.525795,10.737106,9.948417,9.163632,8.421796,7.676055,6.9342184,6.192382,5.4505453,6.3134184,7.1762915,8.039165,8.898132,9.761005,8.972317,8.183627,7.3910336,6.602344,5.813655,6.364176,6.918601,7.4691215,8.023546,8.574067,8.218767,7.859562,7.504261,7.1450562,6.785851,7.8556576,8.921559,9.991365,11.057267,12.123169,12.470661,12.818152,13.165645,13.513136,13.860628,12.400381,10.944039,9.483793,8.023546,6.5633,5.8761253,5.1889505,4.5017757,3.8106966,3.1235218,3.2016098,3.279698,3.357786,3.435874,3.513962,3.4280653,3.3421683,3.2562714,3.174279,3.0883822,3.2836022,3.4788225,3.6740425,3.8692627,4.0644827,4.0644827,4.068387,4.068387,4.0722914,4.0761957,3.9239242,3.775557,3.6232853,3.474918,3.3265507,3.5725281,3.8185053,4.068387,4.3143644,4.564246,4.0332475,3.506153,2.979059,2.4519646,1.9248703,1.9951496,2.0654287,2.135708,2.2059872,2.2762666,2.0380979,1.7999294,1.5617609,1.3235924,1.0893283,1.0268579,0.96829176,0.9058213,0.8472553,0.78868926,0.698888,0.60908675,0.5192855,0.42557985,0.3357786,0.45291066,0.5661383,0.6832704,0.79649806,0.9136301,0.78868926,0.6676528,0.5466163,0.42167544,0.30063897,0.29673457,0.28892577,0.28502136,0.28111696,0.27330816,0.28111696,0.28502136,0.28892577,0.29673457,0.30063897,0.26159495,0.22645533,0.18741131,0.14836729,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.042948425,0.08589685,0.12884527,0.1717937,0.21083772,0.3318742,0.44900626,0.5661383,0.6832704,0.80040246,1.175225,1.5500476,1.9248703,2.2996929,2.6745155,2.8385005,3.0063896,3.1703746,3.3343596,3.4983444,3.5100577,3.521771,3.5295796,3.541293,3.5491016,3.408543,3.2640803,3.1235218,2.979059,2.8385005,2.8463092,2.8580225,2.8658314,2.8775444,2.8892577,3.2679846,3.6467118,4.029343,4.40807,4.786797,5.0210614,5.251421,5.4856853,5.716045,5.950309,6.8405128,7.7307167,8.62092,9.511124,10.401327,9.01136,7.621393,6.2314262,4.841459,3.4514916,3.1391394,2.8306916,2.5183394,2.2098918,1.901444,1.5734742,1.2455044,0.91753453,0.58956474,0.26159495,0.22645533,0.18741131,0.14836729,0.113227665,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.093705654,0.14055848,0.1835069,0.23035973,0.27330816,0.3553006,0.43338865,0.5153811,0.59346914,0.6754616,1.3118792,1.9443923,2.5808098,3.213323,3.8497405,4.2011366,4.5564375,4.9078336,5.2592297,5.610626,5.563773,5.5130157,5.462259,5.4115014,5.3607445,5.278752,5.196759,5.114767,5.0327744,4.950782,4.786797,4.6267166,4.462732,4.298747,4.138666,4.478349,4.8219366,5.165524,5.5091114,5.8487945,5.8566036,5.8644123,5.872221,5.8800297,5.8878384,5.833177,5.7824197,5.7316628,5.677001,5.6262436,5.6379566,5.64967,5.661383,5.6730967,5.688714,6.036206,6.3836975,6.7311897,7.0786815,7.426173,8.062591,8.699008,9.339331,9.975748,10.612165,10.889378,11.166591,11.443803,11.721016,11.998228,12.763491,13.524849,14.286208,15.051471,15.812829,16.863113,17.917301,18.97149,20.021774,21.075964,21.263374,21.450787,21.638197,21.82561,22.01302,22.903223,23.79733,24.69144,25.581644,26.475752,28.51385,30.548042,32.58614,34.62424,36.66234,36.9825,37.302658,37.62282,37.94298,38.26314,37.216763,36.166477,35.1201,34.07372,33.023434,31.297688,29.568039,27.842293,26.116547,24.386896,23.504501,22.622107,21.739712,20.857317,19.974922,19.604004,19.229181,18.858263,18.48344,18.112522,18.768461,19.420496,20.076437,20.732376,21.388315,20.252134,19.115953,17.983677,16.847496,15.711315,15.21936,14.727406,14.235451,13.743496,13.251541,12.408191,11.568744,10.729298,9.889851,9.050405,8.894228,8.741957,8.58578,8.429605,8.273428,8.261715,8.250002,8.238289,8.226576,8.210958,8.55845,8.905942,9.253433,9.600925,9.948417,10.737106,11.525795,12.31058,13.09927,13.887959,14.633699,15.375536,16.121277,16.867018,17.612759,17.628376,17.647898,17.663515,17.683039,17.698656,18.272602,18.84655,19.416592,19.99054,20.560583,20.927597,21.290705,21.657719,22.020828,22.387842,23.289759,24.191677,25.093594,25.999414,26.90133,27.014559,27.131691,27.244919,27.358147,27.475279,26.436708,25.398136,24.36347,23.3249,22.286327,20.049105,17.80798,15.566852,13.325725,11.088503,9.917182,8.745861,7.578445,6.407124,5.2358036,5.743376,6.250948,6.75852,7.266093,7.773665,7.918128,8.058686,8.203149,8.343708,8.488171,7.8556576,7.2270484,6.5984397,5.9659266,5.337318,5.2943697,5.251421,5.2084727,5.169429,5.12648,5.5286336,5.9346914,6.3407493,6.746807,7.1489606,7.164578,7.180196,7.195813,7.211431,7.223144,7.5433054,7.859562,8.175818,8.495979,8.812236,9.784432,10.752724,11.721016,12.693212,13.661504,14.130032,14.59856,15.063184,15.531713,16.00024,14.356487,12.716639,11.072885,9.4291315,7.7892823,7.914223,8.043069,8.171914,8.296855,8.4257,8.827853,9.230007,9.63216,10.034314,10.436467,9.600925,8.761478,7.9259367,7.08649,6.250948,6.036206,5.8214636,5.606722,5.388075,5.173333,5.270943,5.364649,5.4583545,5.5559645,5.64967,5.3295093,5.009348,4.689187,4.369026,4.0488653,4.3065557,4.564246,4.8219366,5.0796275,5.337318,4.728231,4.123049,3.513962,2.9087796,2.2996929,3.4710135,4.646239,5.8175592,6.98888,8.164105,7.5862536,7.008402,6.4305506,5.852699,5.2748475,5.12648,4.9742084,4.825841,4.6735697,4.5252023,4.716518,4.911738,5.1030536,5.2943697,5.4856853,5.6418614,5.7980375,5.9542136,6.1064854,6.262661,6.083059,5.9073606,5.7316628,5.55206,5.376362,5.196759,5.0210614,4.841459,4.6657605,4.4861584,5.3021784,6.1181984,6.9342184,7.746334,8.562354,8.175818,7.7892823,7.3988423,7.012306,6.6257706,7.676055,8.730244,9.784432,10.834716,11.888905,12.548749,13.212498,13.8762455,14.53609,15.199838,15.598087,15.996336,16.39068,16.788929,17.18718,17.230127,17.273075,17.316025,17.358973,17.40192,15.754263,14.106606,12.458947,10.81129,9.163632,9.183154,9.202676,9.2221985,9.24172,9.261242,9.850807,10.436467,11.0260315,11.611692,12.201257,12.056794,11.916236,11.771772,11.631214,11.486752,11.8303385,12.173926,12.513609,12.857197,13.200784,12.435521,11.674163,10.912805,10.151445,9.386183,8.78881,8.191436,7.5940623,6.996689,6.3993154,7.1880045,7.9766936,8.761478,9.550168,10.338858,9.757101,9.17925,8.597494,8.015738,7.437886,7.656533,7.871275,8.089922,8.308568,8.52331,7.9337454,7.3441806,6.754616,6.165051,5.575486,6.348558,7.1216297,7.890797,8.663869,9.43694,9.682918,9.928895,10.170968,10.416945,10.662923,9.741484,8.823949,7.90251,6.9810715,6.0635366,5.64967,5.2358036,4.825841,4.4119744,3.998108,4.0918136,4.185519,4.279225,4.369026,4.462732,4.454923,4.447114,4.4393053,4.4314966,4.423688,4.575959,4.728231,4.884407,5.036679,5.1889505,5.0796275,4.9742084,4.8648853,4.755562,4.650143,4.661856,4.6735697,4.689187,4.7009,4.7126136,4.9468775,5.1772375,5.4115014,5.6418614,5.8761253,5.282656,4.689187,4.095718,3.506153,2.912684,2.8892577,2.8658314,2.8463092,2.822883,2.7994564,2.612045,2.4246337,2.2372224,2.0498111,1.8623998,1.717937,1.5734742,1.4290112,1.2806439,1.1361811,1.0307622,0.92924774,0.8238289,0.71841,0.61299115,0.7066968,0.79649806,0.8902037,0.98390937,1.0737107,0.91753453,0.76135844,0.60127795,0.44510186,0.28892577,0.3279698,0.3670138,0.40605783,0.44900626,0.48805028,0.5114767,0.5309987,0.5544251,0.57785153,0.60127795,0.5231899,0.44900626,0.37482262,0.30063897,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.06637484,0.09761006,0.12884527,0.1639849,0.26940376,0.37872702,0.48414588,0.59346914,0.698888,1.0737107,1.4485333,1.8233559,2.1981785,2.5769055,2.7213683,2.8697357,3.018103,3.1664703,3.310933,3.3265507,3.3421683,3.357786,3.3734035,3.3890212,3.2172275,3.049338,2.8775444,2.7057507,2.5378613,2.541766,2.541766,2.5456703,2.5456703,2.5495746,3.057147,3.5647192,4.0722914,4.579864,5.087436,5.181142,5.270943,5.364649,5.4583545,5.548156,6.3993154,7.2465706,8.093826,8.941081,9.788337,8.6131115,7.4417906,6.27047,5.099149,3.9239242,3.5842414,3.2445583,2.9048753,2.5651922,2.2255092,1.815547,1.4055848,0.9956226,0.58566034,0.1756981,0.14836729,0.12494087,0.10151446,0.07418364,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.11713207,0.16008049,0.20302892,0.24597734,0.28892577,0.359205,0.42557985,0.4958591,0.5661383,0.63641757,1.33921,2.0420024,2.7447948,3.4475873,4.1503797,4.2362766,4.318269,4.4041657,4.4900627,4.575959,4.5369153,4.5017757,4.462732,4.423688,4.388548,4.380739,4.376835,4.3729305,4.369026,4.3612175,4.2753205,4.1894236,4.0996222,4.0137253,3.9239242,4.2557983,4.591577,4.9234514,5.2553253,5.5871997,5.481781,5.3724575,5.263134,5.1577153,5.0483923,4.939069,4.829746,4.7204223,4.6110992,4.5017757,4.5017757,4.5017757,4.5017757,4.5017757,4.5017757,4.677474,4.853172,5.0327744,5.2084727,5.388075,6.126007,6.8639393,7.601871,8.335898,9.073831,9.522837,9.971844,10.416945,10.865952,11.311053,11.900618,12.486279,13.075843,13.661504,14.251068,15.223265,16.195461,17.167656,18.139853,19.11205,19.713327,20.310701,20.911978,21.513256,22.11063,23.344421,24.578213,25.812004,27.04189,28.27568,30.149794,32.023907,33.901924,35.77604,37.65015,38.329517,39.008884,39.688248,40.37152,41.050884,40.258293,39.4696,38.680912,37.88832,37.09963,35.25285,33.406067,31.559284,29.708597,27.861814,27.330816,26.803722,26.272722,25.741724,25.210726,24.574308,23.933987,23.293663,22.653341,22.01302,22.782187,23.551353,24.324427,25.093594,25.86276,24.16044,22.458122,20.755802,19.053482,17.351164,16.46877,15.586374,14.703979,13.821584,12.939189,12.154405,11.365715,10.58093,9.796145,9.01136,8.792714,8.574067,8.351517,8.13287,7.914223,7.9259367,7.9376497,7.9493628,7.9610763,7.9766936,8.339804,8.706817,9.069926,9.43694,9.80005,10.662923,11.525795,12.388668,13.251541,14.114414,14.918721,15.723028,16.527334,17.331642,18.135948,17.96806,17.804073,17.636185,17.468296,17.300406,17.913397,18.530293,19.143284,19.76018,20.37317,20.548868,20.720663,20.892456,21.06425,21.236044,22.071587,22.907127,23.74267,24.578213,25.413754,25.87057,26.33129,26.792007,27.252728,27.713448,26.760773,25.812004,24.863234,23.910559,22.96179,20.716759,18.467823,16.218887,13.973856,11.72492,10.545791,9.366661,8.183627,7.0044975,5.825368,6.266566,6.7116675,7.152865,7.5940623,8.039165,8.121157,8.203149,8.285142,8.367134,8.449126,7.8049,7.1606736,6.5164475,5.8683167,5.22409,5.2045684,5.185046,5.165524,5.1460023,5.12648,5.5091114,5.891743,6.2743745,6.6531014,7.0357327,7.1099167,7.1841,7.2543793,7.328563,7.3988423,7.558923,7.715099,7.871275,8.031356,8.187531,9.17925,10.170968,11.166591,12.158309,13.150026,13.884054,14.614178,15.348206,16.07833,16.812357,15.067088,13.32182,11.576552,9.8312845,8.086017,8.347612,8.609207,8.866898,9.128492,9.386183,10.124115,10.858143,11.592171,12.326198,13.06413,11.912332,10.764437,9.612638,8.460839,7.3129454,6.8639393,6.4188375,5.969831,5.520825,5.0757227,5.040583,5.009348,4.9781127,4.9468775,4.911738,4.5447245,4.1777105,3.8106966,3.4436827,3.076669,3.193801,3.310933,3.4280653,3.5451972,3.6623292,3.4710135,3.2757936,3.084478,2.893162,2.7018464,3.4007344,4.1035266,4.806319,5.5091114,6.211904,6.028397,5.840986,5.657479,5.473972,5.2865605,5.2006636,5.1108627,5.024966,4.939069,4.8492675,5.0718184,5.290465,5.5091114,5.7316628,5.950309,6.2197127,6.4891167,6.75852,7.0318284,7.3012323,7.0903945,6.8795567,6.6687193,6.461786,6.250948,6.126007,6.0049706,5.883934,5.758993,5.6379566,6.211904,6.7819467,7.355894,7.9259367,8.499884,8.250002,8.00012,7.7502384,7.5003567,7.250475,8.160201,9.069926,9.979652,10.889378,11.799104,12.162213,12.525322,12.888432,13.251541,13.610746,14.079274,14.543899,15.008522,15.473146,15.93777,15.918248,15.902631,15.883108,15.867491,15.851873,14.4853325,13.118792,11.756155,10.389614,9.023073,9.105066,9.183154,9.265146,9.343235,9.425227,10.124115,10.826907,11.525795,12.224684,12.923572,12.654168,12.384764,12.11536,11.845957,11.576552,11.92014,12.263727,12.611219,12.954806,13.298394,12.564366,11.826434,11.088503,10.350571,9.612638,9.159728,8.706817,8.253906,7.800996,7.348085,8.062591,8.773191,9.487698,10.198298,10.912805,10.541886,10.170968,9.803954,9.433036,9.062118,8.944985,8.827853,8.710721,8.59359,8.476458,7.6526284,6.8287997,6.008875,5.185046,4.3612175,4.841459,5.3177958,5.794133,6.27047,6.7507114,6.89127,7.0357327,7.1762915,7.320754,7.461313,7.082586,6.703859,6.321227,5.9425,5.563773,5.423215,5.2865605,5.1499066,5.0132523,4.8765984,4.9820175,5.0913405,5.196759,5.3060827,5.4115014,5.481781,5.55206,5.6223392,5.6926184,5.7628975,5.872221,5.9815445,6.0908675,6.2040954,6.3134184,6.094772,5.8761253,5.661383,5.4427366,5.22409,5.3997884,5.575486,5.7511845,5.9268827,6.098676,6.3173227,6.5359693,6.7507114,6.969358,7.1880045,6.5281606,5.872221,5.2162814,4.5564375,3.900498,3.7833657,3.6701381,3.5569105,3.4397783,3.3265507,3.1859922,3.049338,2.912684,2.77603,2.639376,2.4090161,2.1786566,1.9482968,1.717937,1.4875772,1.3665408,1.2494087,1.1283722,1.0073358,0.8862993,0.95657855,1.0268579,1.097137,1.1674163,1.2376955,1.0463798,0.8511597,0.659844,0.46852827,0.27330816,0.359205,0.44510186,0.5309987,0.61689556,0.698888,0.7418364,0.78088045,0.8199245,0.8589685,0.9019169,0.78868926,0.6754616,0.5622339,0.44900626,0.3357786,0.26940376,0.20302892,0.13665408,0.06637484,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.21083772,0.30844778,0.40605783,0.5036679,0.60127795,0.97610056,1.3509232,1.7257458,2.1005683,2.475391,2.6042364,2.7330816,2.8658314,2.9946766,3.1235218,3.1469483,3.1664703,3.1859922,3.2055142,3.2250361,3.0259118,2.8306916,2.631567,2.436347,2.2372224,2.233318,2.2294137,2.2216048,2.2177005,2.2137961,2.8463092,3.4827268,4.1191444,4.7516575,5.388075,5.3412223,5.2943697,5.2436123,5.196759,5.1499066,5.9542136,6.75852,7.5667315,8.371038,9.175345,8.218767,7.266093,6.309514,5.35684,4.4002614,4.029343,3.6584249,3.2914112,2.920493,2.5495746,2.05762,1.5656652,1.0737107,0.58175594,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.14055848,0.1796025,0.21864653,0.26159495,0.30063897,0.359205,0.42167544,0.48024148,0.5388075,0.60127795,1.3704453,2.1396124,2.9087796,3.6818514,4.4510183,4.267512,4.084005,3.9044023,3.7208953,3.5373883,3.513962,3.4866312,3.4632049,3.435874,3.4124475,3.4866312,3.5569105,3.631094,3.7013733,3.775557,3.7638438,3.7482262,3.736513,3.7247996,3.7130866,4.0332475,4.357313,4.6813784,5.001539,5.3256044,5.1030536,4.8805027,4.657952,4.435401,4.21285,4.044961,3.8770714,3.7091823,3.541293,3.3734035,3.3616903,3.349977,3.338264,3.3265507,3.310933,3.3187418,3.3265507,3.3343596,3.3421683,3.349977,4.185519,5.024966,5.8644123,6.699954,7.5394006,8.156297,8.773191,9.390087,10.006983,10.6238785,11.037745,11.4516115,11.861574,12.27544,12.689307,13.579511,14.473619,15.363823,16.25793,17.148134,18.163279,19.174519,20.18576,21.200905,22.212145,23.785618,25.359093,26.928663,28.502136,30.075611,31.785738,33.49977,35.213802,36.92393,38.637966,39.676537,40.71901,41.757584,42.796154,43.838627,43.303726,42.772728,42.24173,41.706825,41.175827,39.208008,37.24019,35.27237,33.30455,31.336733,31.161034,30.981432,30.805735,30.626131,30.450434,29.540707,28.634886,27.729065,26.81934,25.913517,26.795912,27.682213,28.568512,29.450907,30.337206,28.068748,25.796385,23.527927,21.255566,18.987108,17.714273,16.441439,15.168603,13.895767,12.626837,11.896713,11.166591,10.436467,9.706344,8.976221,8.691199,8.406178,8.121157,7.8361354,7.551114,7.5862536,7.6252975,7.6643414,7.699481,7.7385254,8.121157,8.503788,8.886419,9.269051,9.651682,10.588739,11.525795,12.4628525,13.399908,14.336966,15.203742,16.066616,16.933393,17.796265,18.663042,18.311647,17.956347,17.60495,17.253553,16.898252,17.558098,18.214037,18.87388,19.52982,20.18576,20.166237,20.146715,20.127193,20.107672,20.08815,20.853413,21.62258,22.391747,23.15701,23.926178,24.730484,25.53479,26.339098,27.143404,27.951616,27.088743,26.22587,25.362997,24.500124,23.63725,21.380507,19.127666,16.870922,14.618082,12.361338,11.170495,9.983557,8.792714,7.601871,6.4110284,6.7897553,7.168483,7.5433054,7.9220324,8.300759,8.324185,8.343708,8.367134,8.39056,8.413987,7.7541428,7.094299,6.4305506,5.7707067,5.1108627,5.114767,5.1186714,5.1186714,5.1225758,5.12648,5.4856853,5.84489,6.2040954,6.5633,6.9264097,7.055255,7.1841,7.3168497,7.445695,7.57454,7.570636,7.570636,7.5667315,7.5667315,7.562827,8.577971,9.593117,10.608261,11.623405,12.63855,13.634172,14.633699,15.629322,16.628849,17.624472,15.77769,13.930907,12.084125,10.2334385,8.386656,8.781001,9.171441,9.565785,9.956225,10.350571,11.416472,12.486279,13.55218,14.621986,15.687888,14.223738,12.763491,11.29934,9.839094,8.374943,7.6955767,7.016211,6.336845,5.6535745,4.9742084,4.814128,4.6540475,4.493967,4.3338866,4.173806,3.7599394,3.3460727,2.9283018,2.514435,2.1005683,2.077142,2.0537157,2.0341935,2.0107672,1.9873407,2.2098918,2.4324427,2.6549935,2.8775444,3.1000953,3.3343596,3.5647192,3.7989833,4.029343,4.263607,4.4705405,4.677474,4.884407,5.0913405,5.298274,5.2748475,5.251421,5.22409,5.2006636,5.173333,5.423215,5.6691923,5.919074,6.165051,6.4110284,6.7975645,7.1841,7.5667315,7.9532676,8.335898,8.093826,7.8517528,7.60968,7.367607,7.125534,7.0591593,6.98888,6.9225054,6.8561306,6.785851,7.1177254,7.445695,7.7775693,8.109444,8.437413,8.324185,8.210958,8.101635,7.988407,7.8751793,8.644346,9.40961,10.178777,10.944039,11.713207,11.775677,11.838148,11.900618,11.963089,12.025558,12.556558,13.091461,13.622459,14.153459,14.688361,14.610273,14.532186,14.454097,14.376009,14.301826,13.216402,12.134882,11.053363,9.971844,8.886419,9.026978,9.167537,9.308095,9.448653,9.589212,10.401327,11.213444,12.025558,12.837675,13.64979,13.251541,12.853292,12.458947,12.0606985,11.66245,12.009941,12.357433,12.704925,13.052417,13.399908,12.689307,11.974802,11.2642,10.549695,9.839094,9.530646,9.2221985,8.913751,8.609207,8.300759,8.937177,9.573594,10.213917,10.850334,11.486752,11.326671,11.166591,11.00651,10.84643,10.686349,10.2334385,9.784432,9.331521,8.878611,8.4257,7.3715115,6.3134184,5.2592297,4.2050414,3.1508527,3.3343596,3.513962,3.697469,3.8809757,4.0605783,4.1035266,4.142571,4.181615,4.220659,4.263607,4.423688,4.5837684,4.743849,4.903929,5.0640097,5.2006636,5.337318,5.473972,5.610626,5.7511845,5.872221,5.9932575,6.1181984,6.239235,6.364176,6.5086384,6.657006,6.805373,6.9537406,7.098203,7.168483,7.2348576,7.3012323,7.3715115,7.437886,7.1099167,6.7819467,6.453977,6.126007,5.801942,6.13772,6.473499,6.813182,7.1489606,7.4886436,7.6916723,7.890797,8.093826,8.296855,8.499884,7.7775693,7.055255,6.3329406,5.610626,4.8883114,4.6813784,4.4705405,4.263607,4.056674,3.8497405,3.7638438,3.6740425,3.5881457,3.4983444,3.4124475,3.096191,2.7838387,2.4675822,2.1513257,1.8389735,1.7023194,1.5656652,1.4329157,1.2962615,1.1635119,1.2103647,1.2572175,1.3040704,1.3509232,1.4016805,1.1713207,0.94486535,0.71841,0.49195468,0.26159495,0.39434463,0.5231899,0.6520352,0.78088045,0.9136301,0.96829176,1.0268579,1.0854238,1.1439898,1.1986516,1.0502841,0.9019169,0.74964523,0.60127795,0.44900626,0.359205,0.26940376,0.1796025,0.08980125,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.14836729,0.23816854,0.3240654,0.41386664,0.4997635,0.8745861,1.2494087,1.6242313,1.999054,2.3738766,2.4871042,2.6003318,2.7135596,2.8267872,2.9361105,2.9634414,2.9868677,3.0141985,3.0376248,3.0610514,2.8385005,2.612045,2.3855898,2.1630387,1.9365835,1.9248703,1.9131571,1.901444,1.8858263,1.8741131,2.639376,3.4007344,4.1620927,4.9234514,5.688714,5.5013027,5.3138914,5.12648,4.939069,4.7516575,5.5130157,6.2743745,7.0357327,7.800996,8.562354,7.824422,7.08649,6.348558,5.610626,4.8765984,4.474445,4.0761957,3.6740425,3.2757936,2.87364,2.2996929,1.7257458,1.1517987,0.57394713,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.1639849,0.19912452,0.23816854,0.27330816,0.31235218,0.3631094,0.41386664,0.46071947,0.5114767,0.5622339,1.4016805,2.2372224,3.076669,3.912211,4.7516575,4.298747,3.8497405,3.4007344,2.951728,2.4988174,2.4871042,2.475391,2.463678,2.4480603,2.436347,2.5886188,2.736986,2.8892577,3.0376248,3.1859922,3.2484627,3.310933,3.3734035,3.435874,3.4983444,3.8106966,4.123049,4.4393053,4.7516575,5.0640097,4.7243266,4.388548,4.0488653,3.7130866,3.3734035,3.1508527,2.9243972,2.7018464,2.475391,2.2489357,2.2255092,2.1981785,2.174752,2.1513257,2.1239948,1.9639144,1.7999294,1.6359446,1.475864,1.3118792,2.2489357,3.1859922,4.126953,5.0640097,6.001066,6.785851,7.57454,8.36323,9.151918,9.936704,10.174872,10.413041,10.651209,10.889378,11.123642,11.935758,12.751778,13.563893,14.376009,15.188125,16.613232,18.038338,19.463446,20.888552,22.31366,24.226816,26.136068,28.049225,29.962383,31.87554,33.425587,34.975636,36.525684,38.07573,39.62578,41.023556,42.425236,43.826916,45.22469,46.626373,46.34916,46.07585,45.798637,45.52533,45.24812,43.163166,41.07431,38.98936,36.900505,34.81165,34.98735,35.163048,35.338745,35.514442,35.686237,34.511013,33.335785,32.16056,30.98924,29.814016,30.813543,31.81307,32.812595,33.812122,34.81165,31.97315,29.138554,26.300053,23.461554,20.623053,18.963682,17.300406,15.637131,13.973856,12.31058,11.639023,10.963562,10.2881,9.612638,8.937177,8.58578,8.238289,7.8868923,7.5394006,7.1880045,7.250475,7.3129454,7.375416,7.437886,7.5003567,7.898606,8.300759,8.699008,9.101162,9.499411,10.510651,11.525795,12.537036,13.548276,14.56342,15.488764,16.414106,17.33945,18.26089,19.186234,18.651329,18.112522,17.573715,17.03881,16.500004,17.198893,17.901684,18.600573,19.29946,19.998348,19.78751,19.576674,19.36193,19.151093,18.936352,19.639143,20.338032,21.036919,21.735807,22.4386,23.586494,24.738293,25.886187,27.037985,28.18588,27.412807,26.635832,25.86276,25.085785,24.312714,22.048159,19.78751,17.526861,15.262308,13.001659,11.799104,10.600452,9.4018,8.1992445,7.000593,7.3129454,7.6252975,7.9376497,8.250002,8.562354,8.52331,8.488171,8.449126,8.413987,8.374943,7.699481,7.0240197,6.348558,5.6730967,5.001539,5.024966,5.0483923,5.0757227,5.099149,5.12648,5.462259,5.801942,6.13772,6.473499,6.813182,7.000593,7.1880045,7.375416,7.562827,7.7502384,7.5862536,7.426173,7.262188,7.098203,6.9381227,7.9766936,9.01136,10.049932,11.088503,12.123169,13.388195,14.649317,15.914344,17.175465,18.436588,16.48829,14.53609,12.587793,10.6355915,8.687295,9.21439,9.737579,10.260769,10.787864,11.311053,12.712734,14.11051,15.51219,16.91387,18.311647,16.539047,14.762545,12.986042,11.213444,9.43694,8.52331,7.6135845,6.699954,5.786324,4.8765984,4.5876727,4.298747,4.0137253,3.7247996,3.435874,2.9751544,2.514435,2.0498111,1.5890918,1.1244678,0.96438736,0.80040246,0.63641757,0.47633708,0.31235218,0.94876975,1.5890918,2.2255092,2.8619268,3.4983444,3.2640803,3.0259118,2.787743,2.5495746,2.3114061,2.912684,3.513962,4.1113358,4.7126136,5.3138914,5.349031,5.388075,5.423215,5.462259,5.5013027,5.774611,6.0518236,6.3251314,6.5984397,6.8756523,7.375416,7.8751793,8.374943,8.874706,9.37447,9.101162,8.823949,8.550641,8.273428,8.00012,7.988407,7.9766936,7.9610763,7.9493628,7.9376497,8.023546,8.113348,8.1992445,8.289046,8.374943,8.398369,8.4257,8.449126,8.476458,8.499884,9.124588,9.749292,10.373997,10.998701,11.623405,11.389141,11.150972,10.912805,10.674636,10.436467,11.037745,11.639023,12.236397,12.837675,13.438952,13.298394,13.16174,13.025085,12.888432,12.751778,11.951375,11.150972,10.350571,9.550168,8.749765,8.94889,9.151918,9.351044,9.550168,9.749292,10.674636,11.599979,12.525322,13.450665,14.376009,13.848915,13.325725,12.798631,12.27544,11.748346,12.099743,12.4511385,12.798631,13.150026,13.501423,12.814248,12.123169,11.435994,10.748819,10.061645,9.901564,9.737579,9.573594,9.413514,9.249529,9.811763,10.373997,10.936231,11.498465,12.0606985,12.111456,12.162213,12.212971,12.263727,12.31058,11.525795,10.737106,9.948417,9.163632,8.374943,7.08649,5.801942,4.513489,3.2250361,1.9365835,1.8233559,1.7140326,1.6008049,1.4875772,1.3743496,1.3118792,1.2494087,1.1869383,1.1244678,1.0619974,1.7608855,2.463678,3.1625657,3.8614538,4.564246,4.9742084,5.388075,5.801942,6.211904,6.6257706,6.7624245,6.899079,7.0357327,7.1762915,7.3129454,7.5394006,7.7619514,7.988407,8.210958,8.437413,8.460839,8.488171,8.511597,8.538928,8.562354,8.125061,7.687768,7.250475,6.813182,6.375889,6.8756523,7.375416,7.8751793,8.374943,8.874706,9.062118,9.249529,9.43694,9.6243515,9.811763,9.023073,8.238289,7.4495993,6.66091,5.8761253,5.575486,5.2748475,4.9742084,4.6735697,4.376835,4.337791,4.298747,4.263607,4.224563,4.1894236,3.78727,3.3890212,2.9868677,2.5886188,2.1864653,2.0380979,1.8858263,1.737459,1.5890918,1.43682,1.4641509,1.4875772,1.5110037,1.5383345,1.5617609,1.3001659,1.038571,0.77307165,0.5114767,0.24988174,0.42557985,0.60127795,0.77307165,0.94876975,1.1244678,1.1986516,1.2767396,1.3509232,1.4251068,1.4992905,1.3118792,1.1244678,0.93705654,0.74964523,0.5622339,0.44900626,0.3357786,0.22645533,0.113227665,0.0,0.039044023,0.07418364,0.113227665,0.14836729,0.18741131,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.1756981,0.25378615,0.3318742,0.40996224,0.48805028,0.39824903,0.30844778,0.21864653,0.12884527,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.14055848,0.22255093,0.30063897,0.38263142,0.46071947,0.77307165,1.0815194,1.3938715,1.7023194,2.0107672,2.1396124,2.2684577,2.3933985,2.522244,2.6510892,2.6588979,2.6706111,2.67842,2.690133,2.7018464,2.514435,2.330928,2.1435168,1.9600099,1.7765031,1.7608855,1.7452679,1.7296503,1.7140326,1.698415,2.4480603,3.2016098,3.951255,4.7009,5.4505453,5.4310236,5.4115014,5.388075,5.368553,5.349031,5.9151692,6.481308,7.043542,7.60968,8.175818,7.504261,6.8366084,6.165051,5.493494,4.825841,4.4041657,3.9863946,3.5647192,3.1430438,2.7252727,2.1786566,1.6359446,1.0893283,0.5466163,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.07418364,0.062470436,0.05075723,0.039044023,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.14836729,0.19522011,0.24207294,0.28892577,0.3357786,0.43729305,0.5388075,0.63641757,0.737932,0.8394465,1.5734742,2.3075018,3.0415294,3.775557,4.513489,4.0644827,3.619381,3.1703746,2.7213683,2.2762666,2.2137961,2.15523,2.096664,2.0341935,1.9756275,2.1122816,2.2489357,2.3855898,2.5261483,2.6628022,2.7291772,2.795552,2.8658314,2.9322062,2.998581,3.2367494,3.474918,3.7130866,3.951255,4.185519,3.9044023,3.6232853,3.338264,3.057147,2.77603,2.5847144,2.3933985,2.2059872,2.0146716,1.8233559,1.7999294,1.7765031,1.7491722,1.7257458,1.698415,1.5734742,1.4485333,1.3235924,1.1986516,1.0737107,1.8780174,2.67842,3.4827268,4.283129,5.087436,5.825368,6.5633,7.3012323,8.039165,8.773191,9.066022,9.354948,9.643873,9.936704,10.22563,10.998701,11.775677,12.548749,13.325725,14.098797,15.35211,16.605423,17.858736,19.108145,20.361458,22.024733,23.68801,25.351284,27.010654,28.673931,29.876486,31.075138,32.27379,33.476345,34.674995,35.72528,36.77947,37.833656,38.88394,39.93813,39.633587,39.332947,39.028404,38.727764,38.42322,36.740425,35.06153,33.378735,31.695938,30.01314,30.286448,30.555853,30.82916,31.102468,31.375776,30.680794,29.989714,29.298634,28.603651,27.91257,28.693453,29.470428,30.251308,31.032188,31.81307,29.634413,27.455757,25.281004,23.102348,20.92369,19.666473,18.409256,17.152039,15.894821,14.637604,14.258877,13.884054,13.505327,13.1266,12.751778,12.400381,12.0489855,11.701493,11.350098,10.998701,10.920613,10.838621,10.760532,10.67854,10.600452,10.924518,11.2446785,11.568744,11.888905,12.212971,12.989946,13.766922,14.543899,15.320874,16.101755,16.820166,17.538574,18.26089,18.9793,19.701614,19.34241,18.983204,18.627903,18.268698,17.913397,18.526388,19.143284,19.756275,20.37317,20.986162,20.92369,20.861221,20.79875,20.73628,20.67381,21.325846,21.973976,22.62601,23.274141,23.926178,25.273195,26.620214,27.967234,29.314253,30.66127,29.610987,28.556799,27.506514,26.452326,25.398136,23.055496,20.716759,18.374117,16.031475,13.688834,12.486279,11.287627,10.088976,8.886419,7.687768,7.7541428,7.824422,7.890797,7.957172,8.023546,7.941554,7.859562,7.7775693,7.6955767,7.6135845,7.043542,6.473499,5.903456,5.3334136,4.7633705,4.7789884,4.7907014,4.806319,4.8219366,4.8375545,5.1616197,5.4856853,5.813655,6.13772,6.461786,6.7116675,6.9615493,7.211431,7.461313,7.7111945,7.6409154,7.570636,7.504261,7.433982,7.363703,8.4178915,9.47208,10.526268,11.584361,12.63855,13.72007,14.801589,15.883108,16.968533,18.05005,16.402393,14.754736,13.107079,11.45942,9.811763,10.194394,10.573121,10.951848,11.334479,11.713207,12.63855,13.567798,14.493141,15.422389,16.351637,14.875772,13.403813,11.931853,10.459893,8.987934,8.140678,7.2934237,6.446168,5.5989127,4.7516575,4.478349,4.2089458,3.9395418,3.6701381,3.4007344,2.9829633,2.5651922,2.1474214,1.7296503,1.3118792,1.2259823,1.1439898,1.0580931,0.97219616,0.8862993,1.3118792,1.737459,2.1630387,2.5886188,3.0141985,2.8267872,2.6432803,2.455869,2.2723622,2.0888553,2.6081407,3.1313305,3.6545205,4.1777105,4.7009,4.6813784,4.6657605,4.646239,4.630621,4.6110992,4.8492675,5.087436,5.3256044,5.563773,5.7980375,6.2197127,6.6413884,7.0591593,7.480835,7.898606,7.6799593,7.461313,7.238762,7.0201154,6.801469,6.7975645,6.79366,6.79366,6.7897553,6.785851,6.8756523,6.9615493,7.0513506,7.137247,7.223144,7.2582836,7.2934237,7.328563,7.363703,7.3988423,7.8947015,8.39056,8.886419,9.378374,9.874233,9.671205,9.464272,9.261242,9.054309,8.85128,9.405705,9.96013,10.514555,11.06898,11.623405,11.666354,11.705398,11.744442,11.783486,11.826434,11.158782,10.495033,9.8312845,9.163632,8.499884,8.769287,9.0386915,9.308095,9.581403,9.850807,10.584834,11.318862,12.056794,12.790822,13.524849,13.134409,12.743969,12.353529,11.963089,11.576552,11.709302,11.838148,11.970898,12.103647,12.236397,11.756155,11.272009,10.791768,10.307622,9.823476,9.893755,9.964035,10.034314,10.104593,10.174872,10.557504,10.940135,11.322766,11.705398,12.08803,12.326198,12.564366,12.798631,13.036799,13.274967,12.67369,12.068507,11.46723,10.865952,10.260769,9.269051,8.273428,7.277806,6.282183,5.2865605,5.181142,5.0796275,4.9742084,4.8687897,4.7633705,4.806319,4.8492675,4.8883114,4.93126,4.9742084,5.520825,6.0713453,6.617962,7.164578,7.7111945,7.898606,8.082112,8.269524,8.453031,8.636538,8.734148,8.831758,8.929368,9.026978,9.124588,9.37447,9.620447,9.866425,10.116306,10.362284,10.4637985,10.569217,10.670732,10.772245,10.87376,10.61607,10.358379,10.104593,9.846903,9.589212,9.956225,10.327144,10.698062,11.06898,11.435994,11.49456,11.549222,11.603884,11.6585455,11.713207,10.924518,10.135828,9.351044,8.562354,7.773665,7.4027467,7.0318284,6.657006,6.2860875,5.911265,5.7121406,5.5130157,5.3138914,5.1108627,4.911738,4.482254,4.0527697,3.6232853,3.193801,2.7643168,2.6588979,2.5573835,2.455869,2.3543546,2.2489357,2.2762666,2.2996929,2.3231194,2.35045,2.3738766,2.174752,1.9756275,1.7765031,1.5734742,1.3743496,1.43682,1.4992905,1.5617609,1.6242313,1.6867018,1.6710842,1.6515622,1.6359446,1.6164225,1.6008049,1.5110037,1.4251068,1.33921,1.2494087,1.1635119,0.97219616,0.78088045,0.59346914,0.40215343,0.21083772,0.28111696,0.3513962,0.42167544,0.49195468,0.5622339,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.3553006,0.5114767,0.6637484,0.8199245,0.97610056,0.79649806,0.61689556,0.43338865,0.25378615,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.13665408,0.20693332,0.28111696,0.3513962,0.42557985,0.6715572,0.9136301,1.1596074,1.4055848,1.6515622,1.7921207,1.9365835,2.077142,2.2216048,2.3621633,2.358259,2.3543546,2.3465457,2.3426414,2.338737,2.194274,2.0459068,1.901444,1.756981,1.6125181,1.5969005,1.5773785,1.5617609,1.542239,1.5266213,2.260649,2.998581,3.736513,4.474445,5.212377,5.3607445,5.5091114,5.6535745,5.801942,5.950309,6.3173227,6.6843367,7.0513506,7.4183645,7.7892823,7.1841,6.5828223,5.9815445,5.376362,4.775084,4.3338866,3.8965936,3.455396,3.0141985,2.5769055,2.0615244,1.5461433,1.0307622,0.5153811,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.1756981,0.14836729,0.12494087,0.10151446,0.07418364,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.13274968,0.19131571,0.24597734,0.30454338,0.3631094,0.5114767,0.6637484,0.81211567,0.96438736,1.1127546,1.7452679,2.377781,3.0102942,3.6428072,4.2753205,3.8302186,3.3851168,2.9400148,2.494913,2.0498111,1.9443923,1.8350691,1.7257458,1.620327,1.5110037,1.6359446,1.7608855,1.8858263,2.0107672,2.135708,2.2098918,2.2840753,2.3543546,2.4285383,2.4988174,2.6628022,2.8267872,2.9868677,3.1508527,3.310933,3.084478,2.8580225,2.631567,2.4012074,2.174752,2.018576,1.8663043,1.7101282,1.5539521,1.4016805,1.3743496,1.3509232,1.3235924,1.3001659,1.2767396,1.1869383,1.1010414,1.0112402,0.92534333,0.8394465,1.5031948,2.1708477,2.8385005,3.506153,4.173806,4.860981,5.548156,6.239235,6.9264097,7.6135845,7.9532676,8.296855,8.640442,8.98403,9.323712,10.061645,10.799577,11.537509,12.27544,13.013372,14.090988,15.172507,16.254026,17.331642,18.41316,19.826555,21.236044,22.649437,24.062832,25.476225,26.32348,27.17464,28.025799,28.876959,29.724215,30.430912,31.133703,31.8404,32.547096,33.24989,32.92192,32.590046,32.262077,31.930202,31.598328,30.321589,29.044847,27.768108,26.49137,25.210726,25.581644,25.952562,26.32348,26.694399,27.061413,26.854479,26.64364,26.432804,26.221966,26.011127,26.573362,27.131691,27.693926,28.252254,28.81449,27.295675,25.776863,24.25805,22.743143,21.22433,20.37317,19.518106,18.666946,17.815788,16.960724,16.882635,16.800642,16.722555,16.640562,16.562475,16.211079,15.863586,15.51219,15.160794,14.813302,14.590752,14.3682,14.145649,13.923099,13.700547,13.946525,14.188598,14.434575,14.6805525,14.92653,15.469242,16.008049,16.55076,17.093473,17.636185,18.151566,18.666946,19.18233,19.69771,20.21309,20.033487,19.85779,19.678188,19.50249,19.326792,19.853886,20.384884,20.915882,21.446882,21.973976,22.063778,22.149673,22.23557,22.325373,22.411268,23.012547,23.613825,24.211199,24.812477,25.413754,26.955994,28.502136,30.048279,31.590519,33.13666,31.809166,30.477764,29.146362,27.818867,26.487465,24.066736,21.642101,19.221373,16.796738,14.376009,13.173453,11.974802,10.77615,9.573594,8.374943,8.1992445,8.019642,7.843944,7.6643414,7.4886436,7.3597984,7.230953,7.1060123,6.9771667,6.8483214,6.3836975,5.919074,5.45445,4.989826,4.5252023,4.5291066,4.5369153,4.5408196,4.5447245,4.548629,4.860981,5.173333,5.4856853,5.801942,6.114294,6.426646,6.7389984,7.0513506,7.363703,7.676055,7.6955767,7.719003,7.7424297,7.7658563,7.7892823,8.859089,9.932799,11.00651,12.076316,13.150026,14.051944,14.95386,15.855778,16.761599,17.663515,16.316498,14.973383,13.626364,12.28325,10.936231,11.174399,11.408664,11.642927,11.877192,12.111456,12.568271,13.021181,13.477997,13.930907,14.387722,13.216402,12.0489855,10.877665,9.706344,8.538928,7.7541428,6.9732623,6.1884775,5.407597,4.6267166,4.3729305,4.1191444,3.8692627,3.6154766,3.3616903,2.9907722,2.6159496,2.2450314,1.8741131,1.4992905,1.4914817,1.4836729,1.475864,1.4680552,1.4641509,1.6749885,1.8858263,2.1005683,2.3114061,2.5261483,2.3933985,2.260649,2.1278992,1.9951496,1.8623998,2.3075018,2.7526035,3.1977055,3.6428072,4.087909,4.0137253,3.9434462,3.8692627,3.7989833,3.7247996,3.9239242,4.126953,4.3260775,4.5252023,4.7243266,5.0640097,5.4036927,5.743376,6.086963,6.426646,6.2587566,6.094772,5.930787,5.7668023,5.5989127,5.606722,5.6145306,5.6223392,5.630148,5.6379566,5.7238536,5.813655,5.899552,5.989353,6.0752497,6.1181984,6.165051,6.211904,6.2548523,6.3017054,6.6648145,7.0318284,7.394938,7.7619514,8.125061,7.9532676,7.7814736,7.605776,7.433982,7.262188,7.773665,8.281238,8.792714,9.304191,9.811763,10.03041,10.249056,10.4637985,10.682445,10.901091,10.370092,9.839094,9.308095,8.781001,8.250002,8.589685,8.929368,9.269051,9.608734,9.948417,10.495033,11.04165,11.584361,12.130978,12.67369,12.419904,12.166118,11.908427,11.654641,11.400854,11.314958,11.229061,11.143164,11.061172,10.975275,10.698062,10.42085,10.143637,9.866425,9.589212,9.889851,10.194394,10.495033,10.795672,11.100216,11.303245,11.506273,11.709302,11.908427,12.111456,12.537036,12.962616,13.388195,13.813775,14.239355,13.821584,13.403813,12.986042,12.568271,12.150499,11.447707,10.744915,10.042123,9.339331,8.636538,8.538928,8.441318,8.343708,8.246098,8.148487,8.296855,8.445222,8.59359,8.738052,8.886419,9.280765,9.679013,10.073358,10.467703,10.862047,10.819098,10.77615,10.733202,10.694158,10.651209,10.705871,10.764437,10.823003,10.881569,10.936231,11.205634,11.478943,11.748346,12.01775,12.287154,12.466757,12.6463585,12.825961,13.005564,13.189071,13.110983,13.032895,12.954806,12.8767185,12.798631,13.040704,13.2788725,13.520945,13.759113,14.001186,13.923099,13.845011,13.766922,13.688834,13.610746,12.825961,12.037272,11.248583,10.4637985,9.675109,9.230007,8.784905,8.339804,7.8947015,7.4495993,7.08649,6.7233806,6.364176,6.001066,5.6379566,5.1772375,4.716518,4.2557983,3.7989833,3.338264,3.2836022,3.2289407,3.174279,3.1157131,3.0610514,3.0883822,3.1118085,3.1391394,3.1625657,3.1859922,3.049338,2.912684,2.77603,2.639376,2.4988174,2.4480603,2.4012074,2.35045,2.2996929,2.2489357,2.1396124,2.0302892,1.9209659,1.8116426,1.698415,1.7140326,1.7257458,1.737459,1.7491722,1.7608855,1.4953861,1.2259823,0.96048295,0.6910792,0.42557985,0.5270943,0.62860876,0.7340276,0.8355421,0.93705654,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.5309987,0.76526284,0.9956226,1.2298868,1.4641509,1.1908426,0.92143893,0.6520352,0.38263142,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.12884527,0.19131571,0.25769055,0.3240654,0.38653582,0.5661383,0.74574083,0.92924774,1.1088502,1.2884527,1.4446288,1.6008049,1.7608855,1.9170616,2.0732377,2.0537157,2.0341935,2.0146716,1.9951496,1.9756275,1.8702087,1.7647898,1.6593709,1.5539521,1.4485333,1.4290112,1.4094892,1.3899672,1.3704453,1.3509232,2.0732377,2.7994564,3.5256753,4.251894,4.9742084,5.290465,5.606722,5.919074,6.2353306,6.551587,6.719476,6.89127,7.0591593,7.230953,7.3988423,6.8639393,6.329036,5.794133,5.2592297,4.7243266,4.263607,3.8067923,3.3460727,2.8853533,2.4246337,1.9404879,1.456342,0.96829176,0.48414588,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.113227665,0.14836729,0.18741131,0.22645533,0.26159495,0.22645533,0.18741131,0.14836729,0.113227665,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.11713207,0.1835069,0.25378615,0.32016098,0.38653582,0.58566034,0.78868926,0.9878138,1.1869383,1.3860629,1.9170616,2.4480603,2.979059,3.506153,4.037152,3.5959544,3.1508527,2.7096553,2.2684577,1.8233559,1.6710842,1.5149081,1.358732,1.2064602,1.0502841,1.1635119,1.2767396,1.3860629,1.4992905,1.6125181,1.6906061,1.7686942,1.8467822,1.9209659,1.999054,2.0888553,2.174752,2.260649,2.35045,2.436347,2.2645533,2.0927596,1.9209659,1.7491722,1.5734742,1.456342,1.3353056,1.2142692,1.0932326,0.97610056,0.94876975,0.92534333,0.9019169,0.8745861,0.8511597,0.80040246,0.74964523,0.698888,0.6481308,0.60127795,1.1322767,1.6632754,2.1981785,2.7291772,3.2640803,3.900498,4.5369153,5.173333,5.813655,6.4500723,6.844417,7.238762,7.633106,8.031356,8.4257,9.124588,9.823476,10.526268,11.225157,11.924045,12.83377,13.739592,14.649317,15.555139,16.46096,17.624472,18.787983,19.951496,21.111103,22.274614,22.774378,23.274141,23.773905,24.273668,24.773432,25.132637,25.487938,25.847143,26.206348,26.56165,26.206348,25.847143,25.487938,25.132637,24.773432,23.90275,23.028164,22.157482,21.282896,20.412214,20.880743,21.349272,21.813896,22.282423,22.750952,23.02426,23.293663,23.566973,23.84028,24.113588,24.453272,24.792953,25.132637,25.47232,25.812004,24.953035,24.097971,23.239002,22.383938,21.52497,21.075964,20.630861,20.181856,19.736753,19.287746,19.506393,19.721136,19.939783,20.158428,20.37317,20.025679,19.674282,19.326792,18.975395,18.623999,18.26089,17.893875,17.530766,17.163752,16.800642,16.968533,17.136421,17.30431,17.468296,17.636185,17.944633,18.25308,18.56153,18.866072,19.174519,19.486872,19.795319,20.103767,20.416119,20.724567,20.728472,20.728472,20.732376,20.73628,20.73628,21.181383,21.626484,22.071587,22.516687,22.96179,23.199959,23.438128,23.676296,23.914463,24.148727,24.69925,25.24977,25.80029,26.350811,26.90133,28.642694,30.384058,32.129326,33.87069,35.612053,34.00344,32.39873,30.790115,29.181503,27.576794,25.074072,22.57135,20.068628,17.565907,15.063184,13.860628,12.661977,11.4633255,10.260769,9.062118,8.640442,8.218767,7.793187,7.3715115,6.949836,6.7780423,6.606249,6.4305506,6.2587566,6.086963,5.727758,5.368553,5.009348,4.646239,4.2870336,4.283129,4.279225,4.271416,4.267512,4.263607,4.564246,4.860981,5.1616197,5.462259,5.7628975,6.13772,6.5125427,6.8873653,7.262188,7.6370106,7.7541428,7.8673706,7.9805984,8.097731,8.210958,9.304191,10.393518,11.482847,12.572175,13.661504,14.383818,15.1061325,15.828446,16.55076,17.273075,16.2306,15.188125,14.145649,13.103174,12.0606985,12.154405,12.244205,12.334006,12.423808,12.513609,12.494087,12.47847,12.458947,12.44333,12.423808,11.557031,10.690253,9.823476,8.956698,8.086017,7.3715115,6.6531014,5.9346914,5.2162814,4.5017757,4.263607,4.029343,3.795079,3.5608149,3.3265507,2.998581,2.6706111,2.3426414,2.0146716,1.6867018,1.756981,1.8272603,1.8975395,1.9678187,2.0380979,2.0380979,2.0380979,2.0380979,2.0380979,2.0380979,1.9561055,1.8780174,1.796025,1.717937,1.6359446,2.0068626,2.3738766,2.7408905,3.1079042,3.474918,3.3460727,3.2211318,3.0922866,2.9634414,2.8385005,2.998581,3.1625657,3.3265507,3.4866312,3.6506162,3.9083066,4.169902,4.4314966,4.689187,4.950782,4.841459,4.728231,4.618908,4.5095844,4.4002614,4.415879,4.435401,4.4510183,4.4705405,4.4861584,4.575959,4.661856,4.7516575,4.8375545,4.9234514,4.9781127,5.036679,5.0913405,5.1460023,5.2006636,5.434928,5.6691923,5.903456,6.141625,6.375889,6.2353306,6.094772,5.9542136,5.813655,5.6730967,6.141625,6.606249,7.0708723,7.535496,8.00012,8.3944645,8.78881,9.183154,9.581403,9.975748,9.581403,9.183154,8.78881,8.3944645,8.00012,8.410083,8.8200445,9.230007,9.639969,10.049932,10.405232,10.760532,11.115833,11.471134,11.826434,11.705398,11.584361,11.4633255,11.346193,11.225157,10.920613,10.619974,10.319335,10.0147915,9.714153,9.639969,9.565785,9.495506,9.421323,9.351044,9.885946,10.42085,10.955752,11.490656,12.025558,12.0489855,12.068507,12.091934,12.11536,12.138786,12.751778,13.360865,13.973856,14.586847,15.199838,14.965574,14.735214,14.50095,14.27059,14.036326,13.626364,13.216402,12.806439,12.396477,11.986515,11.896713,11.806912,11.717112,11.62731,11.537509,11.791295,12.041177,12.294963,12.548749,12.798631,13.040704,13.286681,13.528754,13.770826,14.012899,13.743496,13.4740925,13.200784,12.93138,12.661977,12.681499,12.697116,12.716639,12.732256,12.751778,13.040704,13.333533,13.626364,13.919194,14.212025,14.469715,14.727406,14.985096,15.242786,15.500477,15.601992,15.7035055,15.808925,15.9104395,16.011953,16.121277,16.234505,16.343828,16.453152,16.562475,16.351637,16.140799,15.933866,15.723028,15.51219,14.723501,13.938716,13.150026,12.361338,11.576552,11.057267,10.541886,10.0226,9.503315,8.987934,8.460839,7.9376497,7.4144597,6.8873653,6.364176,5.872221,5.3841705,4.892216,4.4041657,3.912211,3.9044023,3.8965936,3.8887846,3.8809757,3.873167,3.900498,3.9239242,3.951255,3.9746814,3.998108,3.9239242,3.8497405,3.775557,3.7013733,3.6232853,3.4632049,3.2992198,3.1391394,2.9751544,2.8111696,2.6081407,2.4090161,2.2059872,2.0029583,1.7999294,1.9131571,2.0263848,2.135708,2.2489357,2.3621633,2.018576,1.6710842,1.3274968,0.98390937,0.63641757,0.77307165,0.9058213,1.0424755,1.1791295,1.3118792,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,0.7106012,1.0190489,1.3314011,1.639849,1.9482968,1.5890918,1.2298868,0.8706817,0.5114767,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.12103647,0.1756981,0.23426414,0.29283017,0.3513962,0.46462387,0.58175594,0.6949836,0.80821127,0.92534333,1.097137,1.2689307,1.4407244,1.6164225,1.7882162,1.7530766,1.717937,1.6827974,1.6476578,1.6125181,1.5461433,1.4836729,1.4172981,1.3509232,1.2884527,1.2650263,1.2415999,1.2181735,1.1986516,1.175225,1.8858263,2.6003318,3.310933,4.025439,4.73604,5.2201858,5.704332,6.184573,6.6687193,7.1489606,7.1216297,7.094299,7.066968,7.039637,7.012306,6.5437784,6.0791545,5.610626,5.142098,4.6735697,4.193328,3.7130866,3.2367494,2.7565079,2.2762666,1.8194515,1.3665408,0.9097257,0.45681506,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.14836729,0.19912452,0.24988174,0.30063897,0.3513962,0.30063897,0.24988174,0.19912452,0.14836729,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.10151446,0.1796025,0.25769055,0.3357786,0.41386664,0.6637484,0.9136301,1.1635119,1.4133936,1.6632754,2.0888553,2.5183394,2.9439192,3.3734035,3.7989833,3.3616903,2.920493,2.4792955,2.0380979,1.6008049,1.397776,1.1947471,0.9917182,0.78868926,0.58566034,0.6871748,0.78868926,0.8862993,0.9878138,1.0893283,1.1713207,1.2533131,1.3353056,1.4172981,1.4992905,1.5110037,1.5266213,1.5383345,1.5500476,1.5617609,1.4446288,1.3274968,1.2103647,1.0932326,0.97610056,0.8902037,0.80430686,0.71841,0.63641757,0.5505207,0.5231899,0.4997635,0.47633708,0.44900626,0.42557985,0.41386664,0.39824903,0.38653582,0.37482262,0.3631094,0.76135844,1.1557031,1.5539521,1.9522011,2.35045,2.9361105,3.5256753,4.1113358,4.7009,5.2865605,5.735567,6.180669,6.629675,7.0786815,7.523783,8.187531,8.85128,9.511124,10.174872,10.838621,11.572648,12.306676,13.040704,13.778636,14.512663,15.426293,16.33602,17.24965,18.163279,19.073006,19.225277,19.373644,19.525915,19.674282,19.826555,19.834364,19.846077,19.853886,19.865599,19.873407,19.490776,19.10424,18.72161,18.335073,17.948538,17.483913,17.015385,16.546856,16.07833,15.613705,16.175938,16.742077,17.308216,17.874353,18.436588,19.194042,19.947592,20.701141,21.458595,22.212145,22.333181,22.454218,22.57135,22.692387,22.813423,22.614298,22.419077,22.219954,22.020828,21.82561,21.78266,21.739712,21.696764,21.653814,21.610867,22.126247,22.641628,23.15701,23.67239,24.187773,23.836376,23.488884,23.137487,22.78609,22.4386,21.931028,21.423454,20.915882,20.40831,19.900738,19.99054,20.080341,20.170141,20.259943,20.349745,20.423927,20.494207,20.568392,20.63867,20.712854,20.818274,20.92369,21.02911,21.130625,21.236044,21.41955,21.603058,21.786564,21.966167,22.149673,22.508879,22.868084,23.231194,23.590399,23.949604,24.33614,24.72658,25.113115,25.499651,25.886187,26.38595,26.885714,27.389381,27.889145,28.388908,30.329397,32.26598,34.206467,36.146957,38.087444,36.20162,34.315792,32.43387,30.548042,28.662216,26.081408,23.496693,20.915882,18.33117,15.750359,14.551707,13.349152,12.150499,10.951848,9.749292,9.081639,8.413987,7.746334,7.0786815,6.4110284,6.196286,5.9776397,5.758993,5.5442514,5.3256044,5.0718184,4.814128,4.560342,4.3065557,4.0488653,4.0332475,4.0215344,4.0059166,3.9902992,3.9746814,4.263607,4.548629,4.8375545,5.12648,5.4115014,5.8487945,6.2860875,6.7233806,7.1606736,7.601871,7.8088045,8.015738,8.2226715,8.429605,8.636538,9.745388,10.8542385,11.959184,13.068034,14.176885,14.7156925,15.258404,15.801116,16.343828,16.88654,16.148607,15.406772,14.668839,13.927003,13.189071,13.134409,13.075843,13.021181,12.96652,12.911859,12.423808,11.931853,11.443803,10.951848,10.4637985,9.897659,9.331521,8.769287,8.203149,7.6370106,6.984976,6.3329406,5.6809053,5.02887,4.376835,4.1581883,3.9395418,3.7208953,3.506153,3.2875066,3.0063896,2.7213683,2.4402514,2.1591344,1.8741131,2.0224805,2.1708477,2.3192148,2.463678,2.612045,2.4012074,2.1864653,1.9756275,1.7608855,1.5500476,1.5227169,1.4953861,1.4680552,1.4407244,1.4133936,1.7023194,1.9912452,2.2840753,2.5730011,2.8619268,2.67842,2.4988174,2.3153105,2.1318035,1.9482968,2.0732377,2.1981785,2.3231194,2.4480603,2.5769055,2.7565079,2.9361105,3.1157131,3.2953155,3.474918,3.4202564,3.3655949,3.310933,3.2562714,3.2016098,3.2289407,3.2562714,3.2836022,3.310933,3.338264,3.4241607,3.513962,3.5998588,3.6857557,3.775557,3.8419318,3.9044023,3.970777,4.0332475,4.0996222,4.2050414,4.31046,4.415879,4.521298,4.6267166,4.5173936,4.40807,4.3026514,4.193328,4.087909,4.50568,4.927356,5.349031,5.7668023,6.1884775,6.75852,7.3324676,7.9064145,8.476458,9.050405,8.78881,8.531119,8.269524,8.011833,7.7502384,8.23048,8.710721,9.190963,9.671205,10.151445,10.315431,10.479416,10.6434,10.81129,10.975275,10.990892,11.00651,11.018223,11.033841,11.0494585,10.530173,10.010887,9.491602,8.968412,8.449126,8.581876,8.714626,8.847376,8.980125,9.112875,9.878138,10.647305,11.416472,12.181735,12.950902,12.790822,12.634645,12.47847,12.318389,12.162213,12.962616,13.763018,14.56342,15.363823,16.164225,16.113468,16.066616,16.019762,15.97291,15.926057,15.808925,15.6917925,15.570756,15.453624,15.336493,15.254499,15.172507,15.090515,15.008522,14.92653,15.281831,15.641035,15.996336,16.355541,16.710842,16.800642,16.894348,16.98415,17.073952,17.163752,16.663988,16.168129,15.668366,15.172507,14.676648,14.653222,14.629795,14.606369,14.586847,14.56342,14.875772,15.192029,15.5082855,15.820638,16.136894,16.472673,16.808453,17.14423,17.476105,17.811884,18.096905,18.378021,18.659138,18.94416,19.225277,19.205755,19.186234,19.16671,19.143284,19.123762,18.784079,18.440493,18.096905,17.753317,17.413633,16.624945,15.836256,15.051471,14.262781,13.4740925,12.884527,12.294963,11.705398,11.115833,10.526268,9.839094,9.148014,8.460839,7.773665,7.08649,6.5672045,6.0479193,5.5286336,5.009348,4.4861584,4.5291066,4.5681505,4.607195,4.646239,4.689187,4.7126136,4.73604,4.7633705,4.786797,4.814128,4.7985106,4.786797,4.775084,4.7633705,4.7516575,4.474445,4.2011366,3.9239242,3.6506162,3.3734035,3.0805733,2.7838387,2.4910088,2.194274,1.901444,2.1122816,2.3231194,2.5378613,2.7486992,2.9634414,2.541766,2.1161861,1.6945106,1.2728351,0.8511597,1.0190489,1.1869383,1.3509232,1.5188124,1.6867018,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.8862993,1.2767396,1.6632754,2.0498111,2.436347,1.9873407,1.5383345,1.0893283,0.63641757,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.113227665,0.1639849,0.21083772,0.26159495,0.31235218,0.3631094,0.41386664,0.46071947,0.5114767,0.5622339,0.74964523,0.93705654,1.1244678,1.3118792,1.4992905,1.4485333,1.4016805,1.3509232,1.3001659,1.2494087,1.2259823,1.1986516,1.175225,1.1517987,1.1244678,1.1010414,1.0737107,1.0502841,1.0268579,0.999527,1.698415,2.4012074,3.1000953,3.7989833,4.5017757,5.1499066,5.7980375,6.4500723,7.098203,7.7502384,7.523783,7.3012323,7.0747766,6.8483214,6.6257706,6.223617,5.825368,5.423215,5.024966,4.6267166,4.126953,3.6232853,3.1235218,2.6237583,2.1239948,1.698415,1.2767396,0.8511597,0.42557985,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.18741131,0.24988174,0.31235218,0.37482262,0.43729305,0.37482262,0.31235218,0.24988174,0.18741131,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08589685,0.1756981,0.26159495,0.3513962,0.43729305,0.737932,1.038571,1.33921,1.6359446,1.9365835,2.260649,2.5886188,2.912684,3.2367494,3.5608149,3.1235218,2.6862288,2.2489357,1.8116426,1.3743496,1.1244678,0.8745861,0.62470436,0.37482262,0.12494087,0.21083772,0.30063897,0.38653582,0.47633708,0.5622339,0.6481308,0.737932,0.8238289,0.9136301,0.999527,0.93705654,0.8745861,0.81211567,0.74964523,0.6871748,0.62470436,0.5622339,0.4997635,0.43729305,0.37482262,0.3240654,0.27330816,0.22645533,0.1756981,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.38653582,0.6481308,0.9136301,1.175225,1.43682,1.9756275,2.514435,3.049338,3.5881457,4.123049,4.6267166,5.12648,5.6262436,6.126007,6.6257706,7.250475,7.8751793,8.499884,9.124588,9.749292,10.311526,10.87376,11.435994,11.998228,12.564366,13.224211,13.887959,14.551707,15.211552,15.875299,15.676175,15.473146,15.274021,15.074897,14.875772,14.53609,14.200311,13.860628,13.524849,13.189071,12.775204,12.361338,11.951375,11.537509,11.123642,11.061172,10.998701,10.936231,10.87376,10.81129,11.475039,12.138786,12.798631,13.462379,14.126127,15.363823,16.601519,17.839214,19.07691,20.310701,20.21309,20.111576,20.013966,19.91245,19.810938,20.27556,20.73628,21.200905,21.661623,22.126247,22.489357,22.848562,23.211672,23.574781,23.937891,24.750006,25.562122,26.374237,27.186354,27.998468,27.650976,27.29958,26.948185,26.600693,26.249296,25.601166,24.949131,24.300999,23.648964,23.000834,23.012547,23.02426,23.035973,23.05159,23.063305,22.899319,22.739239,22.575254,22.411268,22.251188,22.149673,22.048159,21.95055,21.849035,21.751425,22.11063,22.47374,22.83685,23.199959,23.563068,23.836376,24.113588,24.386896,24.664108,24.937418,25.476225,26.011127,26.549934,27.088743,27.623646,28.076557,28.525562,28.97457,29.423576,29.876486,32.012196,34.151806,36.287514,38.42322,40.562836,38.399796,36.23676,34.07372,31.910679,29.751545,27.088743,24.425941,21.763138,19.100336,16.437534,15.238882,14.036326,12.837675,11.639023,10.436467,9.526741,8.6131115,7.699481,6.785851,5.8761253,5.610626,5.349031,5.087436,4.825841,4.564246,4.4119744,4.263607,4.1113358,3.9629683,3.8106966,3.78727,3.7638438,3.736513,3.7130866,3.6857557,3.9629683,4.2362766,4.513489,4.786797,5.0640097,5.563773,6.0635366,6.5633,7.0630636,7.562827,7.8634663,8.164105,8.460839,8.761478,9.062118,10.186585,11.311053,12.439425,13.563893,14.688361,15.051471,15.410676,15.773785,16.136894,16.500004,16.062712,15.625418,15.188125,14.750832,14.313539,14.114414,13.911386,13.712261,13.513136,13.314012,12.349625,11.389141,10.424754,9.464272,8.499884,8.238289,7.9766936,7.7111945,7.4495993,7.1880045,6.5984397,6.012779,5.423215,4.8375545,4.251894,4.0488653,3.8497405,3.6506162,3.4514916,3.2484627,3.0141985,2.77603,2.5378613,2.2996929,2.0615244,2.2879796,2.514435,2.736986,2.9634414,3.1859922,2.7643168,2.338737,1.9131571,1.4875772,1.0619974,1.0893283,1.1127546,1.1361811,1.1635119,1.1869383,1.4016805,1.6125181,1.8233559,2.0380979,2.2489357,2.0107672,1.7765031,1.5383345,1.3001659,1.0619974,1.1517987,1.2376955,1.3235924,1.4133936,1.4992905,1.6008049,1.698415,1.7999294,1.901444,1.999054,1.999054,1.999054,1.999054,1.999054,1.999054,2.0380979,2.0732377,2.1122816,2.1513257,2.1864653,2.2762666,2.3621633,2.4480603,2.5378613,2.6237583,2.7018464,2.77603,2.8502135,2.9243972,2.998581,2.9751544,2.951728,2.9243972,2.900971,2.87364,2.7994564,2.7252727,2.6510892,2.5769055,2.4988174,2.87364,3.2484627,3.6232853,3.998108,4.376835,5.12648,5.8761253,6.6257706,7.375416,8.125061,8.00012,7.8751793,7.7502384,7.6252975,7.5003567,8.050878,8.601398,9.151918,9.698535,10.249056,10.22563,10.198298,10.174872,10.151445,10.124115,10.276386,10.424754,10.573121,10.725393,10.87376,10.135828,9.4018,8.663869,7.9259367,7.1880045,7.523783,7.8634663,8.1992445,8.538928,8.874706,9.874233,10.87376,11.873287,12.8767185,13.8762455,13.536563,13.200784,12.861101,12.525322,12.185639,13.173453,14.161267,15.14908,16.136894,17.124708,17.261362,17.40192,17.538574,17.675228,17.811884,17.987581,18.163279,18.338978,18.51077,18.68647,18.612286,18.538101,18.463919,18.38583,18.311647,18.77627,19.23699,19.701614,20.162333,20.623053,20.560583,20.498112,20.435642,20.37317,20.310701,19.588387,18.862167,18.135948,17.413633,16.687416,16.624945,16.562475,16.500004,16.437534,16.375063,16.710842,17.050524,17.386303,17.725986,18.061766,18.475632,18.885593,19.29946,19.713327,20.12329,20.587914,21.048632,21.513256,21.973976,22.4386,22.286327,22.13796,21.98569,21.837322,21.688955,21.212618,20.73628,20.263847,19.78751,19.311174,18.526388,17.7377,16.94901,16.164225,15.375536,14.711788,14.048039,13.388195,12.724447,12.0606985,11.213444,10.362284,9.511124,8.663869,7.812709,7.262188,6.7116675,6.1611466,5.610626,5.0640097,5.1499066,5.2358036,5.3256044,5.4115014,5.5013027,5.5247293,5.548156,5.575486,5.5989127,5.6262436,5.6730967,5.7238536,5.774611,5.825368,5.8761253,5.4856853,5.099149,4.7126136,4.3260775,3.9356375,3.5491016,3.1625657,2.77603,2.3855898,1.999054,2.3114061,2.6237583,2.9361105,3.2484627,3.5608149,3.0610514,2.5612879,2.0615244,1.5617609,1.0619974,1.261122,1.4641509,1.6632754,1.8623998,2.0615244,0.5622339,0.62470436,0.6871748,0.74964523,0.81211567,0.8745861,1.1400855,1.4055848,1.6710842,1.9365835,2.1981785,1.7921207,1.3860629,0.97610056,0.5700427,0.1639849,0.12884527,0.09761006,0.06637484,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.10932326,0.15227169,0.19912452,0.24207294,0.28892577,0.3318742,0.3709182,0.41386664,0.45681506,0.4997635,0.6559396,0.80821127,0.96438736,1.1205635,1.2767396,1.2376955,1.1986516,1.1635119,1.1244678,1.0893283,1.0737107,1.0619974,1.0502841,1.038571,1.0268579,1.0112402,0.999527,0.9878138,0.97610056,0.96438736,1.6008049,2.2372224,2.87364,3.513962,4.1503797,4.7789884,5.4036927,6.0323014,6.66091,7.2856145,7.008402,6.7311897,6.453977,6.1767645,5.899552,5.5559645,5.2084727,4.8648853,4.521298,4.173806,3.7521305,3.330455,2.9087796,2.4831998,2.0615244,1.6515622,1.2415999,0.8316377,0.42167544,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.16008049,0.21864653,0.28111696,0.339683,0.39824903,0.3553006,0.30844778,0.26549935,0.21864653,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08199245,0.1639849,0.24597734,0.3318742,0.41386664,0.7106012,1.0112402,1.3118792,1.6125181,1.9131571,2.1786566,2.4480603,2.7135596,2.9829633,3.2484627,2.8306916,2.4090161,1.9912452,1.5695697,1.1517987,0.94096094,0.7301232,0.5192855,0.30844778,0.10151446,0.1717937,0.23816854,0.30844778,0.37872702,0.44900626,0.5231899,0.59346914,0.6676528,0.7418364,0.81211567,0.77307165,0.7340276,0.6910792,0.6520352,0.61299115,0.5544251,0.4958591,0.44119745,0.38263142,0.3240654,0.28111696,0.23426414,0.19131571,0.14446288,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.30844778,0.5192855,0.7301232,0.94096094,1.1517987,1.6008049,2.0498111,2.4988174,2.951728,3.4007344,3.8692627,4.3338866,4.802415,5.270943,5.735567,6.289992,6.8405128,7.394938,7.9493628,8.499884,9.0465,9.593117,10.143637,10.690253,11.23687,11.834243,12.431617,13.028991,13.626364,14.223738,14.079274,13.934812,13.790349,13.645885,13.501423,13.282777,13.06413,12.845484,12.630741,12.412095,12.056794,11.697589,11.338385,10.983084,10.6238785,10.510651,10.401327,10.2881,10.174872,10.061645,10.48332,10.901091,11.322766,11.740538,12.162213,13.079747,13.997282,14.914817,15.832351,16.749886,16.679607,16.609327,16.539047,16.46877,16.398489,16.777216,17.155943,17.530766,17.909492,18.28822,18.64352,19.002726,19.358027,19.717232,20.076437,20.884647,21.69286,22.504974,23.313187,24.125301,24.043308,23.965221,23.883228,23.805141,23.723148,23.445936,23.164818,22.883701,22.60649,22.325373,22.4386,22.551826,22.66115,22.774378,22.887606,22.821232,22.75876,22.692387,22.62601,22.563541,22.493261,22.426888,22.360512,22.294136,22.223858,22.665054,23.106253,23.543545,23.984743,24.425941,24.835903,25.24977,25.663635,26.073599,26.487465,26.971611,27.455757,27.943808,28.427954,28.912098,29.263494,29.618795,29.970192,30.321589,30.67689,32.226936,33.77308,35.323128,36.873177,38.42322,36.61158,34.79994,32.988297,31.176653,29.361105,26.600693,23.836376,21.075964,18.311647,15.551234,14.383818,13.220306,12.056794,10.889378,9.725866,8.913751,8.105539,7.2934237,6.4852123,5.6730967,5.462259,5.251421,5.036679,4.825841,4.6110992,4.50568,4.4041657,4.298747,4.193328,4.087909,4.1113358,4.1308575,4.154284,4.1777105,4.2011366,4.474445,4.743849,5.017157,5.290465,5.563773,5.9542136,6.3407493,6.7311897,7.1216297,7.5120697,7.8751793,8.238289,8.601398,8.960603,9.323712,10.471607,11.615597,12.759586,13.903577,15.051471,15.605896,16.16032,16.714746,17.26917,17.823597,17.308216,16.796738,16.281357,15.765976,15.250595,15.098324,14.946052,14.79378,14.641508,14.489237,13.4740925,12.458947,11.443803,10.4286585,9.413514,9.093353,8.773191,8.453031,8.13287,7.812709,7.2036223,6.5984397,5.989353,5.3841705,4.775084,4.6813784,4.591577,4.4978714,4.4041657,4.3143644,4.462732,4.6110992,4.7633705,4.911738,5.0640097,5.3295093,5.591104,5.8566036,6.1221027,6.387602,5.661383,4.93126,4.2050414,3.4788225,2.7486992,2.822883,2.893162,2.9673457,3.0415294,3.1118085,3.1898966,3.2679846,3.3460727,3.4241607,3.4983444,3.252367,3.0063896,2.7565079,2.5105307,2.260649,2.2216048,2.182561,2.1435168,2.1044729,2.0615244,2.0498111,2.0380979,2.0263848,2.0107672,1.999054,1.9600099,1.9209659,1.8819219,1.8389735,1.7999294,1.8389735,1.8819219,1.9209659,1.9600099,1.999054,2.084951,2.1708477,2.2567444,2.338737,2.4246337,2.455869,2.4831998,2.514435,2.5456703,2.5769055,2.5769055,2.5769055,2.5769055,2.5769055,2.5769055,2.522244,2.4714866,2.416825,2.366068,2.3114061,2.6237583,2.9361105,3.2484627,3.5608149,3.873167,4.4861584,5.099149,5.7121406,6.3251314,6.9381227,6.89127,6.8405128,6.79366,6.746807,6.699954,7.1450562,7.590158,8.03526,8.480362,8.925464,8.925464,8.925464,8.925464,8.925464,8.925464,9.101162,9.280765,9.456462,9.636065,9.811763,9.323712,8.831758,8.343708,7.8517528,7.363703,7.6838636,8.007929,8.32809,8.652155,8.976221,9.86252,10.748819,11.639023,12.525322,13.411622,13.181262,12.950902,12.720543,12.494087,12.263727,13.075843,13.887959,14.700074,15.51219,16.324306,16.574188,16.82407,17.073952,17.323833,17.573715,17.749413,17.92511,18.10081,18.276506,18.448301,18.362404,18.276506,18.186707,18.10081,18.011007,18.381926,18.752844,19.123762,19.490776,19.861694,19.853886,19.842173,19.834364,19.82265,19.810938,19.229181,18.64352,18.057861,17.4722,16.88654,16.765503,16.640562,16.519526,16.398489,16.273548,16.59371,16.909966,17.226223,17.546383,17.86264,18.124235,18.38583,18.651329,18.912924,19.174519,19.416592,19.65476,19.896833,20.135002,20.37317,20.236517,20.095959,19.9554,19.814842,19.674282,19.190138,18.705992,18.217941,17.733795,17.24965,16.628849,16.008049,15.391153,14.770353,14.149553,13.477997,12.810344,12.138786,11.471134,10.799577,10.159255,9.515028,8.870802,8.23048,7.5862536,7.094299,6.5984397,6.1025805,5.606722,5.1108627,5.138193,5.169429,5.196759,5.22409,5.251421,5.2475166,5.2436123,5.2436123,5.239708,5.2358036,5.2045684,5.173333,5.138193,5.1069584,5.0757227,4.8765984,4.6735697,4.474445,4.2753205,4.0761957,3.7130866,3.349977,2.9868677,2.6237583,2.260649,2.4910088,2.7213683,2.951728,3.182088,3.4124475,3.0063896,2.6042364,2.1981785,1.7921207,1.3860629,1.5656652,1.7413634,1.9209659,2.096664,2.2762666,1.1244678,1.1517987,1.175225,1.1986516,1.2259823,1.2494087,1.3938715,1.53443,1.678893,1.8194515,1.9639144,1.5969005,1.2337911,0.8667773,0.5036679,0.13665408,0.10932326,0.08199245,0.05466163,0.027330816,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.10151446,0.14055848,0.1835069,0.22255093,0.26159495,0.29673457,0.3318742,0.3670138,0.40215343,0.43729305,0.5583295,0.6832704,0.80430686,0.92924774,1.0502841,1.0268579,0.999527,0.97610056,0.94876975,0.92534333,0.92534333,0.92534333,0.92534333,0.92534333,0.92534333,0.92534333,0.92534333,0.92534333,0.92534333,0.92534333,1.4992905,2.0732377,2.6510892,3.2250361,3.7989833,4.4041657,5.009348,5.6145306,6.2197127,6.824895,6.4969254,6.165051,5.833177,5.505207,5.173333,4.884407,4.5954814,4.3065557,4.0137253,3.7247996,3.3812122,3.0337205,2.690133,2.3465457,1.999054,1.6047094,1.2103647,0.8160201,0.42167544,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.13274968,0.19131571,0.24597734,0.30454338,0.3631094,0.3357786,0.30844778,0.28111696,0.25378615,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.078088045,0.15617609,0.23426414,0.30844778,0.38653582,0.6871748,0.9878138,1.2884527,1.5890918,1.8858263,2.096664,2.3075018,2.5183394,2.7291772,2.9361105,2.533957,2.1318035,1.7296503,1.3274968,0.92534333,0.75354964,0.58566034,0.41386664,0.24597734,0.07418364,0.12884527,0.1796025,0.23426414,0.28502136,0.3357786,0.39434463,0.45291066,0.5114767,0.5661383,0.62470436,0.60908675,0.58956474,0.57394713,0.5544251,0.5388075,0.48414588,0.43338865,0.37872702,0.3279698,0.27330816,0.23426414,0.19522011,0.15617609,0.113227665,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.015617609,0.031235218,0.046852827,0.058566034,0.07418364,0.23426414,0.39044023,0.5466163,0.7066968,0.8628729,1.2259823,1.5890918,1.9482968,2.3114061,2.6745155,3.1118085,3.5451972,3.978586,4.415879,4.8492675,5.3295093,5.8097506,6.289992,6.7702336,7.250475,7.7814736,8.316377,8.847376,9.378374,9.913278,10.444276,10.979179,11.510178,12.041177,12.576079,12.486279,12.396477,12.306676,12.216875,12.123169,12.029464,11.931853,11.834243,11.736633,11.639023,11.334479,11.033841,10.729298,10.4286585,10.124115,9.964035,9.80005,9.636065,9.475985,9.311999,9.491602,9.6673,9.846903,10.0226,10.198298,10.795672,11.39695,11.994324,12.591698,13.189071,13.146122,13.107079,13.068034,13.028991,12.986042,13.2788725,13.571702,13.864532,14.157363,14.450192,14.801589,15.15689,15.5082855,15.859682,16.211079,17.019289,17.827501,18.635712,19.443924,20.24823,20.439547,20.630861,20.818274,21.009588,21.200905,21.290705,21.380507,21.470308,21.56011,21.64991,21.860748,22.07549,22.286327,22.50107,22.711908,22.743143,22.778282,22.809519,22.840754,22.875893,22.840754,22.805614,22.770473,22.735334,22.700195,23.215576,23.734861,24.254147,24.769527,25.288813,25.839334,26.38595,26.936472,27.486992,28.037512,28.470901,28.90429,29.333775,29.767162,30.200552,30.454338,30.708124,30.965815,31.2196,31.473387,32.437775,33.39826,34.362644,35.323128,36.287514,34.823364,33.363117,31.898966,30.43872,28.97457,26.112642,23.250715,20.388788,17.526861,14.661031,13.532659,12.404286,11.272009,10.143637,9.01136,8.304664,7.5979667,6.89127,6.180669,5.473972,5.3138914,5.1499066,4.985922,4.825841,4.661856,4.60329,4.5408196,4.482254,4.423688,4.3612175,4.4314966,4.5017757,4.572055,4.6423345,4.7126136,4.9820175,5.251421,5.520825,5.794133,6.0635366,6.3407493,6.621866,6.902983,7.1841,7.461313,7.8868923,8.312472,8.738052,9.163632,9.589212,10.752724,11.916236,13.083652,14.247164,15.410676,16.16032,16.906061,17.655706,18.401447,19.151093,18.557625,17.964155,17.370686,16.78112,16.187653,16.082233,15.976814,15.871395,15.765976,15.660558,14.594656,13.528754,12.458947,11.393045,10.323239,9.948417,9.56969,9.190963,8.81614,8.437413,7.8088045,7.1841,6.5554914,5.9268827,5.298274,5.3138914,5.3295093,5.3451266,5.3607445,5.376362,5.911265,6.4500723,6.98888,7.523783,8.062591,8.367134,8.671678,8.976221,9.280765,9.589212,8.55845,7.5276875,6.4969254,5.466163,4.4393053,4.5564375,4.677474,4.7985106,4.9156423,5.036679,4.9781127,4.9234514,4.8648853,4.806319,4.7516575,4.493967,4.2362766,3.978586,3.7208953,3.4632049,3.2953155,3.1274261,2.959537,2.7916477,2.6237583,2.4988174,2.3738766,2.2489357,2.1239948,1.999054,1.9209659,1.8389735,1.7608855,1.678893,1.6008049,1.6437533,1.6867018,1.7257458,1.7686942,1.8116426,1.893635,1.9756275,2.0615244,2.1435168,2.2255092,2.2098918,2.194274,2.1786566,2.1669433,2.1513257,2.174752,2.1981785,2.2255092,2.2489357,2.2762666,2.2450314,2.2137961,2.1864653,2.15523,2.1239948,2.3738766,2.6237583,2.87364,3.1235218,3.3734035,3.8497405,4.3260775,4.7985106,5.2748475,5.7511845,5.7785153,5.8097506,5.840986,5.8683167,5.899552,6.239235,6.578918,6.918601,7.2582836,7.601871,7.6252975,7.648724,7.676055,7.699481,7.726812,7.929841,8.136774,8.339804,8.546737,8.749765,8.507692,8.265619,8.023546,7.7814736,7.5394006,7.843944,8.152391,8.460839,8.769287,9.073831,9.850807,10.6238785,11.400854,12.173926,12.950902,12.825961,12.704925,12.583888,12.458947,12.337912,12.974329,13.610746,14.251068,14.8874855,15.523903,15.8870125,16.250122,16.613232,16.976341,17.33945,17.511244,17.686943,17.86264,18.038338,18.214037,18.112522,18.011007,17.913397,17.811884,17.714273,17.991486,18.268698,18.54591,18.823124,19.100336,19.143284,19.186234,19.229181,19.268225,19.311174,18.866072,18.420969,17.975868,17.530766,17.085665,16.906061,16.722555,16.539047,16.359446,16.175938,16.472673,16.769407,17.066143,17.366781,17.663515,17.776743,17.886066,17.999294,18.112522,18.22575,18.241367,18.26089,18.276506,18.296028,18.311647,18.182802,18.053955,17.921206,17.79236,17.663515,17.167656,16.671797,16.175938,15.683984,15.188125,14.735214,14.282304,13.829392,13.376482,12.923572,12.24811,11.568744,10.893282,10.213917,9.538455,9.101162,8.667773,8.234385,7.7970915,7.363703,6.9225054,6.481308,6.044015,5.602817,5.1616197,5.1303844,5.099149,5.0640097,5.0327744,5.001539,4.970304,4.939069,4.911738,4.8805027,4.8492675,4.73604,4.618908,4.50568,4.388548,4.2753205,4.263607,4.251894,4.2362766,4.224563,4.21285,3.873167,3.5373883,3.2016098,2.8619268,2.5261483,2.6706111,2.8189783,2.9673457,3.1157131,3.2640803,2.951728,2.6432803,2.330928,2.0224805,1.7140326,1.8663043,2.0224805,2.1786566,2.330928,2.4871042,1.6867018,1.6749885,1.6632754,1.6515622,1.6359446,1.6242313,1.6437533,1.6632754,1.6867018,1.7062237,1.7257458,1.4016805,1.0815194,0.75745404,0.43338865,0.113227665,0.08980125,0.06637484,0.046852827,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.09761006,0.13274968,0.1678893,0.20302892,0.23816854,0.26549935,0.29283017,0.32016098,0.3474918,0.37482262,0.46462387,0.5544251,0.6442264,0.7340276,0.8238289,0.81211567,0.80040246,0.78868926,0.77307165,0.76135844,0.77307165,0.78868926,0.80040246,0.81211567,0.8238289,0.8394465,0.8511597,0.8628729,0.8745861,0.8862993,1.4016805,1.9131571,2.4246337,2.9361105,3.4514916,4.0332475,4.6150036,5.196759,5.7785153,6.364176,5.9815445,5.5989127,5.2162814,4.83365,4.4510183,4.2167544,3.978586,3.7443218,3.5100577,3.2757936,3.0063896,2.7408905,2.4714866,2.2059872,1.9365835,1.5578566,1.1791295,0.79649806,0.41777104,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.10541886,0.16008049,0.21474212,0.26940376,0.3240654,0.31625658,0.30454338,0.29673457,0.28502136,0.27330816,0.21864653,0.1639849,0.10932326,0.05466163,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07418364,0.14446288,0.21864653,0.28892577,0.3631094,0.6637484,0.96438736,1.261122,1.5617609,1.8623998,2.0146716,2.1669433,2.3192148,2.4714866,2.6237583,2.241127,1.8545911,1.4680552,1.0854238,0.698888,0.5700427,0.44119745,0.30844778,0.1796025,0.05075723,0.08589685,0.12103647,0.15617609,0.19131571,0.22645533,0.26940376,0.30844778,0.3513962,0.39434463,0.43729305,0.44119745,0.44900626,0.45291066,0.45681506,0.46071947,0.41386664,0.3670138,0.32016098,0.27330816,0.22645533,0.19131571,0.15617609,0.12103647,0.08589685,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.15617609,0.26159495,0.3631094,0.46852827,0.57394713,0.8511597,1.1244678,1.4016805,1.6749885,1.9482968,2.3543546,2.7565079,3.1586614,3.5608149,3.9629683,4.369026,4.7789884,5.185046,5.591104,6.001066,6.5164475,7.0357327,7.551114,8.070399,8.58578,9.054309,9.522837,9.991365,10.455989,10.924518,10.889378,10.8542385,10.819098,10.783959,10.748819,10.772245,10.795672,10.819098,10.838621,10.862047,10.61607,10.366188,10.120211,9.874233,9.6243515,9.413514,9.198771,8.987934,8.773191,8.562354,8.495979,8.433509,8.367134,8.300759,8.238289,8.515501,8.792714,9.069926,9.347139,9.6243515,9.616543,9.60483,9.593117,9.585307,9.573594,9.780528,9.991365,10.198298,10.405232,10.612165,10.959657,11.307149,11.654641,12.002132,12.349625,13.153932,13.958238,14.766449,15.570756,16.375063,16.835783,17.296501,17.753317,18.214037,18.674755,19.135475,19.596195,20.056915,20.51373,20.97445,21.2868,21.599154,21.911505,22.223858,22.53621,22.668959,22.797804,22.926651,23.0594,23.188246,23.184341,23.184341,23.180437,23.176533,23.176533,23.77,24.36347,24.960844,25.554314,26.151686,26.838861,27.526035,28.213211,28.900385,29.58756,29.966288,30.348919,30.727646,31.106373,31.489004,31.64518,31.801357,31.961437,32.117615,32.27379,32.648613,33.023434,33.39826,33.77308,34.151806,33.03905,31.926298,30.813543,29.700788,28.588034,25.624592,22.66115,19.701614,16.738173,13.774731,12.681499,11.584361,10.491129,9.393991,8.300759,7.6955767,7.0903945,6.4852123,5.8800297,5.2748475,5.1616197,5.0483923,4.939069,4.825841,4.7126136,4.6969957,4.6813784,4.6657605,4.6540475,4.6384296,4.755562,4.872694,4.989826,5.1069584,5.22409,5.493494,5.758993,6.028397,6.2938967,6.5633,6.7311897,6.902983,7.0708723,7.2426662,7.4105554,7.898606,8.386656,8.874706,9.362757,9.850807,11.033841,12.220779,13.403813,14.590752,15.773785,16.714746,17.655706,18.596668,19.533724,20.474686,19.803127,19.135475,18.463919,17.796265,17.124708,17.066143,17.01148,16.952915,16.894348,16.835783,15.719124,14.59856,13.477997,12.357433,11.23687,10.803481,10.366188,9.932799,9.499411,9.062118,8.413987,7.7658563,7.1216297,6.473499,5.825368,5.9464045,6.0713453,6.192382,6.3134184,6.4383593,7.363703,8.289046,9.21439,10.135828,11.061172,11.408664,11.752251,12.095839,12.44333,12.786918,11.455516,10.124115,8.78881,7.4574084,6.126007,6.2938967,6.461786,6.6257706,6.79366,6.9615493,6.7702336,6.578918,6.3836975,6.192382,6.001066,5.7316628,5.466163,5.196759,4.93126,4.661856,4.369026,4.0722914,3.7794614,3.4827268,3.1859922,2.951728,2.7135596,2.475391,2.2372224,1.999054,1.8819219,1.7608855,1.639849,1.5188124,1.4016805,1.4446288,1.4914817,1.53443,1.5812829,1.6242313,1.7062237,1.7843118,1.8663043,1.9443923,2.0263848,1.9639144,1.9053483,1.8467822,1.7843118,1.7257458,1.7765031,1.8233559,1.8741131,1.9248703,1.9756275,1.9678187,1.9600099,1.9522011,1.9443923,1.9365835,2.1239948,2.3114061,2.4988174,2.6862288,2.87364,3.213323,3.5491016,3.8887846,4.224563,4.564246,4.6696653,4.7789884,4.884407,4.9937305,5.099149,5.3334136,5.571582,5.805846,6.04011,6.2743745,6.3251314,6.375889,6.426646,6.473499,6.524256,6.75852,6.98888,7.223144,7.453504,7.687768,7.6916723,7.6955767,7.703386,7.70729,7.7111945,8.0040245,8.296855,8.589685,8.882515,9.175345,9.839094,10.498938,11.162686,11.826434,12.486279,12.470661,12.458947,12.44333,12.427712,12.412095,12.8767185,13.337439,13.798158,14.262781,14.723501,15.199838,15.676175,16.148607,16.624945,17.101282,17.273075,17.448774,17.624472,17.800169,17.975868,17.86264,17.749413,17.636185,17.526861,17.413633,17.597141,17.780647,17.96806,18.151566,18.338978,18.432684,18.526388,18.623999,18.717705,18.81141,18.506866,18.202324,17.89778,17.593237,17.288692,17.04662,16.800642,16.55857,16.316498,16.074425,16.351637,16.628849,16.906061,17.183275,17.464392,17.425346,17.386303,17.351164,17.31212,17.273075,17.070047,16.863113,16.660084,16.453152,16.250122,16.129086,16.008049,15.890917,15.76988,15.648844,15.145176,14.641508,14.133936,13.630268,13.1266,12.841579,12.556558,12.271536,11.986515,11.701493,11.014318,10.331048,9.643873,8.960603,8.273428,8.046973,7.8205175,7.5940623,7.363703,7.137247,6.7507114,6.36808,5.9815445,5.5989127,5.212377,5.1186714,5.02887,4.9351645,4.841459,4.7516575,4.6930914,4.6345253,4.575959,4.521298,4.462732,4.263607,4.068387,3.8692627,3.6740425,3.474918,3.6506162,3.8263142,3.998108,4.173806,4.349504,4.037152,3.7247996,3.4124475,3.1000953,2.787743,2.854118,2.9165885,2.9829633,3.049338,3.1118085,2.8970666,2.6823244,2.4675822,2.25284,2.0380979,2.1708477,2.3035975,2.436347,2.5690966,2.7018464,2.2489357,2.1981785,2.1513257,2.1005683,2.0498111,1.999054,1.8975395,1.796025,1.6906061,1.5890918,1.4875772,1.2064602,0.92924774,0.6481308,0.3670138,0.08589685,0.07027924,0.05075723,0.03513962,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.093705654,0.12103647,0.15227169,0.1835069,0.21083772,0.23426414,0.25378615,0.27330816,0.29283017,0.31235218,0.3709182,0.42557985,0.48414588,0.5427119,0.60127795,0.60127795,0.60127795,0.60127795,0.60127795,0.60127795,0.62470436,0.6481308,0.6754616,0.698888,0.7262188,0.74964523,0.77307165,0.80040246,0.8238289,0.8511597,1.3001659,1.7491722,2.1981785,2.6510892,3.1000953,3.6584249,4.220659,4.7789884,5.3412223,5.899552,5.466163,5.02887,4.5954814,4.1581883,3.7247996,3.5451972,3.3655949,3.1859922,3.0063896,2.8267872,2.6354716,2.4441557,2.2567444,2.0654287,1.8741131,1.5110037,1.1439898,0.78088045,0.41386664,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.078088045,0.12884527,0.1835069,0.23426414,0.28892577,0.29673457,0.30063897,0.30844778,0.31625658,0.3240654,0.26159495,0.19522011,0.12884527,0.06637484,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06637484,0.13665408,0.20302892,0.26940376,0.3357786,0.63641757,0.93705654,1.2376955,1.5383345,1.8389735,1.9326792,2.0263848,2.1239948,2.2177005,2.3114061,1.9443923,1.5773785,1.2103647,0.8433509,0.47633708,0.38653582,0.29673457,0.20693332,0.113227665,0.023426414,0.042948425,0.058566034,0.078088045,0.093705654,0.113227665,0.14055848,0.1678893,0.19522011,0.22255093,0.24988174,0.27721256,0.30454338,0.3318742,0.359205,0.38653582,0.3435874,0.30063897,0.26159495,0.21864653,0.1756981,0.14446288,0.113227665,0.08589685,0.05466163,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.078088045,0.12884527,0.1835069,0.23426414,0.28892577,0.47633708,0.6637484,0.8511597,1.038571,1.2259823,1.5969005,1.9639144,2.3348327,2.7057507,3.076669,3.408543,3.7443218,4.0801005,4.415879,4.7516575,5.251421,5.755089,6.2587566,6.75852,7.262188,7.6643414,8.066495,8.468649,8.870802,9.276859,9.296382,9.315904,9.335425,9.354948,9.37447,9.518932,9.659492,9.803954,9.944512,10.088976,9.893755,9.702439,9.511124,9.315904,9.124588,8.862993,8.601398,8.335898,8.074304,7.812709,7.504261,7.195813,6.89127,6.5828223,6.2743745,6.2314262,6.1884775,6.1455293,6.1064854,6.0635366,6.083059,6.1025805,6.1221027,6.141625,6.1611466,6.2860875,6.407124,6.5281606,6.6531014,6.774138,7.1177254,7.461313,7.800996,8.144583,8.488171,9.288573,10.09288,10.893282,11.697589,12.497992,13.228115,13.958238,14.688361,15.418485,16.148607,16.980246,17.811884,18.639616,19.471254,20.298986,20.712854,21.12672,21.536682,21.95055,22.364416,22.590872,22.817327,23.043781,23.274141,23.500597,23.531832,23.559164,23.590399,23.621634,23.648964,24.324427,24.995983,25.66754,26.339098,27.010654,27.838388,28.662216,29.486046,30.31378,31.137608,31.465578,31.793547,32.121517,32.445583,32.773552,32.83602,32.89459,32.953156,33.015625,33.074192,32.863354,32.648613,32.437775,32.22303,32.012196,31.250835,30.485573,29.724215,28.962856,28.201498,25.136541,22.07549,19.010534,15.949483,12.888432,11.826434,10.768341,9.706344,8.648251,7.5862536,7.08649,6.5828223,6.0791545,5.579391,5.0757227,5.0132523,4.950782,4.8883114,4.825841,4.7633705,4.7907014,4.8219366,4.853172,4.884407,4.911738,5.0757227,5.2436123,5.407597,5.571582,5.735567,6.001066,6.266566,6.532065,6.7975645,7.0630636,7.1216297,7.1841,7.2426662,7.3012323,7.363703,7.914223,8.460839,9.01136,9.561881,10.112402,11.318862,12.521418,13.727879,14.934339,16.136894,17.26917,18.401447,19.533724,20.666,21.798277,21.052536,20.306797,19.557152,18.81141,18.061766,18.053955,18.042242,18.034433,18.02272,18.011007,16.839687,15.668366,14.493141,13.32182,12.150499,11.6585455,11.166591,10.670732,10.178777,9.686822,9.019169,8.351517,7.6838636,7.016211,6.348558,6.578918,6.8092775,7.039637,7.269997,7.5003567,8.812236,10.124115,11.435994,12.751778,14.063657,14.446288,14.832824,15.21936,15.601992,15.988527,14.352583,12.716639,11.080693,9.448653,7.812709,8.027451,8.242193,8.456935,8.671678,8.886419,8.55845,8.234385,7.9064145,7.578445,7.250475,6.9732623,6.6960497,6.4188375,6.141625,5.8644123,5.4388323,5.017157,4.5954814,4.173806,3.7482262,3.4007344,3.049338,2.7018464,2.35045,1.999054,1.8389735,1.678893,1.5188124,1.358732,1.1986516,1.2494087,1.2962615,1.3431144,1.3899672,1.43682,1.5149081,1.5929961,1.6710842,1.7491722,1.8233559,1.7218413,1.6164225,1.5110037,1.4055848,1.3001659,1.3743496,1.4485333,1.5266213,1.6008049,1.6749885,1.6906061,1.7062237,1.7218413,1.7335546,1.7491722,1.8741131,1.999054,2.1239948,2.2489357,2.3738766,2.5769055,2.77603,2.9751544,3.174279,3.3734035,3.5608149,3.7443218,3.9317331,4.11524,4.298747,4.4314966,4.560342,4.689187,4.8180323,4.950782,5.024966,5.099149,5.173333,5.251421,5.3256044,5.5832953,5.84489,6.1064854,6.364176,6.6257706,6.8756523,7.1294384,7.3832245,7.633106,7.8868923,8.164105,8.441318,8.718531,8.995743,9.276859,9.823476,10.373997,10.924518,11.475039,12.025558,12.119265,12.209065,12.302772,12.396477,12.486279,12.775204,13.06413,13.349152,13.638077,13.923099,14.512663,15.098324,15.687888,16.273548,16.863113,17.03881,17.210606,17.386303,17.562002,17.7377,17.612759,17.487818,17.362877,17.237936,17.112995,17.206701,17.296501,17.390207,17.483913,17.573715,17.722082,17.87045,18.018816,18.163279,18.311647,18.147661,17.983677,17.815788,17.651802,17.487818,17.183275,16.882635,16.578093,16.277452,15.976814,16.2306,16.48829,16.745981,17.003672,17.261362,17.073952,16.88654,16.69913,16.511717,16.324306,15.8987255,15.469242,15.043662,14.614178,14.188598,14.079274,13.966047,13.856724,13.7474,13.638077,13.122696,12.607315,12.091934,11.576552,11.061172,10.944039,10.826907,10.709775,10.592644,10.475512,9.780528,9.089449,8.398369,7.703386,7.012306,6.9927845,6.9732623,6.9537406,6.9342184,6.910792,6.5828223,6.250948,5.9229784,5.591104,5.263134,5.1108627,4.958591,4.806319,4.6540475,4.5017757,4.415879,4.3299823,4.2440853,4.1581883,4.0761957,3.795079,3.513962,3.2367494,2.9556324,2.6745155,3.0376248,3.4007344,3.7638438,4.123049,4.4861584,4.2011366,3.912211,3.6232853,3.338264,3.049338,3.0337205,3.0141985,2.998581,2.979059,2.9634414,2.8424048,2.7213683,2.6042364,2.4831998,2.3621633,2.4714866,2.5808098,2.6940374,2.803361,2.912684,2.8111696,2.7252727,2.639376,2.5495746,2.463678,2.3738766,2.1513257,1.9248703,1.698415,1.475864,1.2494087,1.0112402,0.77307165,0.5388075,0.30063897,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.08589685,0.113227665,0.13665408,0.1639849,0.18741131,0.19912452,0.21083772,0.22645533,0.23816854,0.24988174,0.27330816,0.30063897,0.3240654,0.3513962,0.37482262,0.38653582,0.39824903,0.41386664,0.42557985,0.43729305,0.47633708,0.5114767,0.5505207,0.58566034,0.62470436,0.6637484,0.698888,0.737932,0.77307165,0.81211567,1.1986516,1.5890918,1.9756275,2.3621633,2.7486992,3.2875066,3.8263142,4.3612175,4.900025,5.4388323,4.950782,4.462732,3.9746814,3.4866312,2.998581,2.87364,2.7486992,2.6237583,2.4988174,2.3738766,2.260649,2.1513257,2.0380979,1.9248703,1.8116426,1.4641509,1.1127546,0.76135844,0.41386664,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10151446,0.14836729,0.19912452,0.24988174,0.27330816,0.30063897,0.3240654,0.3513962,0.37482262,0.30063897,0.22645533,0.14836729,0.07418364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.61299115,0.9136301,1.2142692,1.5110037,1.8116426,1.8506867,1.8858263,1.9248703,1.9639144,1.999054,1.6515622,1.3001659,0.94876975,0.60127795,0.24988174,0.19912452,0.14836729,0.10151446,0.05075723,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.113227665,0.1639849,0.21083772,0.26159495,0.31235218,0.27330816,0.23816854,0.19912452,0.1639849,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10151446,0.19912452,0.30063897,0.39824903,0.4997635,0.8394465,1.175225,1.5110037,1.8506867,2.1864653,2.4480603,2.7135596,2.9751544,3.2367494,3.4983444,3.9863946,4.474445,4.9624953,5.4505453,5.938596,6.2743745,6.6140575,6.949836,7.2856145,7.6252975,7.699481,7.773665,7.8517528,7.9259367,8.00012,8.261715,8.52331,8.78881,9.050405,9.311999,9.175345,9.0386915,8.898132,8.761478,8.624825,8.312472,8.00012,7.687768,7.375416,7.0630636,6.5125427,5.9620223,5.4115014,4.860981,4.3143644,3.951255,3.5881457,3.2250361,2.8619268,2.4988174,2.5495746,2.6003318,2.6510892,2.7018464,2.7486992,2.787743,2.8267872,2.8619268,2.900971,2.9361105,3.2757936,3.611572,3.951255,4.2870336,4.6267166,5.423215,6.223617,7.0240197,7.824422,8.624825,9.6243515,10.6238785,11.623405,12.626837,13.626364,14.825015,16.023666,17.226223,18.424873,19.623526,20.138906,20.650383,21.16186,21.673336,22.188719,22.512783,22.83685,23.160913,23.488884,23.81295,23.87542,23.937891,24.00036,24.062832,24.125301,24.874947,25.624592,26.374237,27.123882,27.873528,28.837915,29.798397,30.762785,31.723269,32.687656,32.960964,33.23818,33.511486,33.788696,34.062004,34.026867,33.987823,33.948776,33.91364,33.874596,33.074192,32.27379,31.473387,30.67689,29.876486,29.46262,29.048752,28.63879,28.224924,27.811058,24.64849,21.485926,18.32336,15.160794,11.998228,10.975275,9.948417,8.925464,7.898606,6.8756523,6.473499,6.0752497,5.6730967,5.2748475,4.8765984,4.860981,4.8492675,4.8375545,4.825841,4.814128,4.8883114,4.9624953,5.036679,5.1108627,5.1889505,5.3997884,5.610626,5.825368,6.036206,6.250948,6.5125427,6.774138,7.0357327,7.3012323,7.562827,7.5120697,7.461313,7.4105554,7.363703,7.3129454,7.9259367,8.538928,9.151918,9.761005,10.373997,11.599979,12.825961,14.051944,15.274021,16.500004,17.823597,19.151093,20.474686,21.798277,23.125774,22.29804,21.474213,20.650383,19.826555,18.998821,19.037865,19.07691,19.11205,19.151093,19.186234,17.964155,16.738173,15.51219,14.286208,13.06413,12.513609,11.963089,11.412568,10.862047,10.311526,9.6243515,8.937177,8.250002,7.562827,6.8756523,7.211431,7.551114,7.8868923,8.226576,8.562354,10.260769,11.963089,13.661504,15.363823,17.062239,17.487818,17.913397,18.338978,18.760653,19.186234,17.24965,15.313066,13.376482,11.435994,9.499411,9.761005,10.0265045,10.2881,10.549695,10.81129,10.350571,9.885946,9.425227,8.960603,8.499884,8.210958,7.9259367,7.6370106,7.348085,7.0630636,6.5125427,5.9620223,5.4115014,4.860981,4.3143644,3.8497405,3.3890212,2.9243972,2.463678,1.999054,1.7999294,1.6008049,1.4016805,1.1986516,0.999527,1.0502841,1.1010414,1.1517987,1.1986516,1.2494087,1.3235924,1.4016805,1.475864,1.5500476,1.6242313,1.475864,1.3235924,1.175225,1.0268579,0.8745861,0.97610056,1.0737107,1.175225,1.2767396,1.3743496,1.4133936,1.4485333,1.4875772,1.5266213,1.5617609,1.6242313,1.6867018,1.7491722,1.8116426,1.8741131,1.9365835,1.999054,2.0615244,2.1239948,2.1864653,2.4519646,2.7135596,2.9751544,3.2367494,3.4983444,3.5256753,3.5491016,3.5764325,3.5998588,3.6232853,3.7247996,3.8263142,3.9239242,4.025439,4.123049,4.4119744,4.7009,4.985922,5.2748475,5.563773,6.0635366,6.5633,7.0630636,7.562827,8.062591,8.324185,8.58578,8.85128,9.112875,9.37447,9.811763,10.249056,10.686349,11.123642,11.560935,11.763964,11.963089,12.162213,12.361338,12.564366,12.67369,12.786918,12.900145,13.013372,13.1266,13.825488,14.524376,15.223265,15.926057,16.624945,16.800642,16.976341,17.148134,17.323833,17.49953,17.362877,17.226223,17.085665,16.94901,16.812357,16.812357,16.812357,16.812357,16.812357,16.812357,17.01148,17.210606,17.413633,17.612759,17.811884,17.788456,17.761126,17.7377,17.714273,17.686943,17.323833,16.960724,16.601519,16.238409,15.875299,16.113468,16.351637,16.585901,16.82407,17.062239,16.72646,16.386776,16.050997,15.711315,15.375536,14.723501,14.07537,13.423335,12.775204,12.123169,12.025558,11.924045,11.826434,11.72492,11.623405,11.100216,10.573121,10.049932,9.526741,8.999647,9.050405,9.101162,9.151918,9.198771,9.249529,8.550641,7.8517528,7.1489606,6.4500723,5.7511845,5.938596,6.126007,6.3134184,6.5008297,6.688241,6.4110284,6.13772,5.8644123,5.5871997,5.3138914,5.099149,4.8883114,4.6735697,4.462732,4.251894,4.138666,4.025439,3.912211,3.7989833,3.6857557,3.3265507,2.9634414,2.6003318,2.2372224,1.8741131,2.4246337,2.9751544,3.5256753,4.0761957,4.6267166,4.3612175,4.0996222,3.8380275,3.5764325,3.310933,3.213323,3.1118085,3.0141985,2.912684,2.8111696,2.787743,2.7643168,2.736986,2.7135596,2.6862288,2.77603,2.8619268,2.951728,3.0376248,3.1235218,2.6862288,2.5612879,2.4324427,2.3035975,2.1786566,2.0498111,1.8389735,1.6281357,1.4212024,1.2103647,0.999527,0.80821127,0.62079996,0.42948425,0.23816854,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.07418364,0.093705654,0.11713207,0.14055848,0.1639849,0.1756981,0.18741131,0.19912452,0.21083772,0.22645533,0.24597734,0.26940376,0.29283017,0.31625658,0.3357786,0.3474918,0.359205,0.3670138,0.37872702,0.38653582,0.43338865,0.47633708,0.5231899,0.5661383,0.61299115,0.6481308,0.6871748,0.7262188,0.76135844,0.80040246,1.1400855,1.4797685,1.8194515,2.1591344,2.4988174,3.0298162,3.5608149,4.0918136,4.618908,5.1499066,4.7516575,4.349504,3.951255,3.5491016,3.1508527,2.9634414,2.7799344,2.5964274,2.4090161,2.2255092,2.077142,1.9287747,1.7843118,1.6359446,1.4875772,1.1986516,0.9136301,0.62470436,0.3357786,0.05075723,0.05075723,0.05466163,0.058566034,0.058566034,0.062470436,0.05075723,0.042948425,0.031235218,0.023426414,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.22645533,0.24988174,0.27330816,0.30063897,0.3240654,0.26549935,0.20693332,0.14446288,0.08589685,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05075723,0.10541886,0.15617609,0.21083772,0.26159495,0.4997635,0.737932,0.97610056,1.2142692,1.4485333,1.4953861,1.5383345,1.5851873,1.6281357,1.6749885,1.3860629,1.0932326,0.80430686,0.5153811,0.22645533,0.1796025,0.13665408,0.08980125,0.046852827,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.08980125,0.12884527,0.1717937,0.21083772,0.24988174,0.21864653,0.19131571,0.16008049,0.12884527,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.078088045,0.16008049,0.23816854,0.32016098,0.39824903,0.6715572,0.94096094,1.2103647,1.4797685,1.7491722,1.9600099,2.1708477,2.3816853,2.5886188,2.7994564,3.193801,3.5881457,3.9863946,4.380739,4.775084,5.040583,5.3060827,5.571582,5.833177,6.098676,6.1611466,6.223617,6.2860875,6.348558,6.4110284,6.6335793,6.852226,7.0708723,7.2934237,7.5120697,7.406651,7.297328,7.1880045,7.082586,6.9732623,6.7702336,6.5633,6.3602715,6.153338,5.950309,5.5950084,5.239708,4.884407,4.5291066,4.173806,3.9629683,3.7482262,3.5373883,3.3265507,3.1118085,3.2094188,3.3031244,3.39683,3.49444,3.5881457,3.5100577,3.4319696,3.3538816,3.2757936,3.2016098,3.455396,3.7091823,3.9668727,4.220659,4.474445,5.153811,5.8292727,6.5086384,7.1841,7.8634663,8.738052,9.612638,10.487225,11.361811,12.236397,13.25935,14.282304,15.305257,16.32821,17.351164,17.921206,18.495153,19.069101,19.639143,20.21309,20.63867,21.068155,21.493734,21.923218,22.348799,22.590872,22.82904,23.071114,23.309282,23.551353,24.273668,24.999887,25.726107,26.448421,27.17464,27.951616,28.724688,29.501663,30.274734,31.051712,31.317211,31.586615,31.852114,32.121517,32.387016,32.289406,32.191795,32.094185,31.996576,31.898966,31.231314,30.559757,29.888199,29.220547,28.548988,27.900858,27.256632,26.608501,25.960371,25.31224,22.602585,19.89293,17.183275,14.473619,11.763964,10.795672,9.82738,8.859089,7.890797,6.9264097,6.6257706,6.329036,6.0323014,5.735567,5.4388323,5.481781,5.520825,5.563773,5.606722,5.64967,5.7668023,5.8800297,5.9932575,6.1103897,6.223617,6.5008297,6.7819467,7.0591593,7.336372,7.6135845,7.8634663,8.117252,8.371038,8.62092,8.874706,8.781001,8.691199,8.597494,8.503788,8.413987,8.859089,9.304191,9.749292,10.194394,10.6355915,11.603884,12.572175,13.540467,14.508759,15.473146,16.683512,17.893875,19.10424,20.314606,21.52497,20.951023,20.37317,19.799223,19.225277,18.651329,18.631807,18.61619,18.596668,18.58105,18.56153,17.48001,16.398489,15.313066,14.231546,13.150026,12.798631,12.4511385,12.099743,11.748346,11.400854,10.783959,10.170968,9.554072,8.941081,8.324185,8.55845,8.78881,9.023073,9.253433,9.487698,10.877665,12.267632,13.657599,15.047566,16.437534,17.124708,17.811884,18.499058,19.186234,19.873407,18.163279,16.449247,14.739119,13.025085,11.311053,11.45942,11.607788,11.756155,11.904523,12.0489855,11.771772,11.49456,11.217348,10.940135,10.662923,10.194394,9.725866,9.261242,8.792714,8.324185,7.703386,7.08649,6.46569,5.84489,5.22409,5.009348,4.794606,4.579864,4.365122,4.1503797,3.7443218,3.338264,2.9361105,2.5300527,2.1239948,2.1083772,2.096664,2.0810463,2.0654287,2.0498111,2.0263848,1.999054,1.9756275,1.9482968,1.9248703,1.7882162,1.6554666,1.5188124,1.3860629,1.2494087,1.2884527,1.3235924,1.3626363,1.4016805,1.43682,1.4641509,1.4875772,1.5110037,1.5383345,1.5617609,1.6047094,1.6476578,1.6906061,1.7335546,1.7765031,1.815547,1.8584955,1.901444,1.9443923,1.9873407,2.2059872,2.4207294,2.639376,2.8580225,3.076669,3.1039999,3.135235,3.1664703,3.193801,3.2250361,3.3070288,3.3890212,3.4710135,3.5569105,3.638903,3.892689,4.1464753,4.4041657,4.657952,4.911738,5.3295093,5.74728,6.165051,6.5828223,7.000593,7.2426662,7.4847393,7.726812,7.968885,8.210958,8.59359,8.972317,9.351044,9.733675,10.112402,10.311526,10.506746,10.705871,10.901091,11.100216,11.186112,11.268105,11.354002,11.4398985,11.525795,12.08803,12.654168,13.220306,13.786445,14.348679,14.458001,14.571229,14.6805525,14.789876,14.899199,14.774258,14.645412,14.516567,14.391626,14.262781,14.254972,14.247164,14.239355,14.231546,14.223738,14.376009,14.528281,14.6805525,14.836729,14.989,14.949956,14.9109125,14.875772,14.836729,14.801589,14.504854,14.208119,13.91529,13.618555,13.325725,13.477997,13.634172,13.790349,13.946525,14.098797,13.821584,13.540467,13.25935,12.978233,12.70102,12.185639,11.6702585,11.154878,10.639496,10.124115,10.03041,9.936704,9.839094,9.745388,9.651682,9.230007,8.8083315,8.39056,7.968885,7.551114,7.590158,7.629202,7.6682463,7.7111945,7.7502384,7.1880045,6.629675,6.0713453,5.5091114,4.950782,5.0913405,5.2358036,5.376362,5.520825,5.661383,5.45445,5.2475166,5.040583,4.83365,4.6267166,4.4978714,4.369026,4.2440853,4.11524,3.9863946,3.9395418,3.892689,3.8458362,3.7989833,3.7482262,3.4124475,3.076669,2.736986,2.4012074,2.0615244,2.592523,3.1235218,3.6506162,4.181615,4.7126136,4.462732,4.21285,3.9629683,3.7130866,3.4632049,3.3655949,3.2679846,3.1703746,3.0727646,2.9751544,2.8892577,2.803361,2.7213683,2.6354716,2.5495746,2.541766,2.5300527,2.5183394,2.5105307,2.4988174,2.5612879,2.3933985,2.2294137,2.0615244,1.893635,1.7257458,1.5305257,1.3353056,1.1400855,0.94486535,0.74964523,0.60908675,0.46462387,0.3240654,0.1796025,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.058566034,0.078088045,0.09761006,0.11713207,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.19912452,0.21864653,0.23816854,0.26159495,0.28111696,0.30063897,0.30844778,0.31625658,0.3240654,0.3318742,0.3357786,0.39044023,0.44119745,0.4958591,0.5466163,0.60127795,0.63641757,0.6754616,0.7106012,0.74964523,0.78868926,1.0815194,1.3743496,1.6632754,1.9561055,2.2489357,2.7721257,3.2953155,3.8185053,4.3416953,4.860981,4.548629,4.2362766,3.9239242,3.611572,3.2992198,3.0532427,2.8111696,2.5651922,2.3192148,2.0732377,1.893635,1.7101282,1.5266213,1.3431144,1.1635119,0.93705654,0.7106012,0.48805028,0.26159495,0.039044023,0.05466163,0.07418364,0.08980125,0.10932326,0.12494087,0.10541886,0.08589685,0.06637484,0.046852827,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.058566034,0.08980125,0.12103647,0.14836729,0.1756981,0.19912452,0.22645533,0.24988174,0.27330816,0.23035973,0.1835069,0.14055848,0.093705654,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.042948425,0.08589685,0.12884527,0.1717937,0.21083772,0.38653582,0.5622339,0.737932,0.9136301,1.0893283,1.1400855,1.1908426,1.2455044,1.2962615,1.3509232,1.1205635,0.8902037,0.659844,0.42948425,0.19912452,0.16008049,0.12103647,0.078088045,0.039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0078088045,0.015617609,0.023426414,0.031235218,0.039044023,0.06637484,0.09761006,0.12884527,0.15617609,0.18741131,0.1639849,0.14055848,0.12103647,0.09761006,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058566034,0.12103647,0.1796025,0.23816854,0.30063897,0.5036679,0.7066968,0.9058213,1.1088502,1.3118792,1.4719596,1.6281357,1.7843118,1.9443923,2.1005683,2.4012074,2.7057507,3.0063896,3.310933,3.611572,3.8067923,3.998108,4.1894236,4.380739,4.575959,4.6267166,4.6735697,4.7243266,4.775084,4.825841,5.001539,5.181142,5.35684,5.5364423,5.7121406,5.6340523,5.5559645,5.481781,5.4036927,5.3256044,5.2279944,5.1303844,5.0327744,4.9351645,4.8375545,4.677474,4.5173936,4.357313,4.1972322,4.037152,3.9746814,3.912211,3.8497405,3.78727,3.7247996,3.8653584,4.0059166,4.1464753,4.283129,4.423688,4.2323723,4.041056,3.8458362,3.6545205,3.4632049,3.6349986,3.8067923,3.978586,4.154284,4.3260775,4.8805027,5.434928,5.989353,6.5437784,7.098203,7.8517528,8.601398,9.351044,10.100689,10.850334,11.693685,12.54094,13.384291,14.231546,15.074897,15.70741,16.339924,16.972437,17.60495,18.237463,18.768461,19.29946,19.826555,20.357553,20.888552,21.306324,21.724094,22.141865,22.555733,22.973503,23.676296,24.375183,25.074072,25.776863,26.475752,27.061413,27.650976,28.236637,28.826202,29.411861,29.673458,29.931149,30.192743,30.454338,30.712029,30.555853,30.395771,30.239595,30.08342,29.92334,29.384531,28.845724,28.306917,27.764204,27.225397,26.343002,25.460608,24.578213,23.695818,22.813423,20.556679,18.296028,16.039284,13.78254,11.525795,10.61607,9.706344,8.796618,7.8868923,6.9732623,6.7780423,6.5867267,6.3915067,6.196286,6.001066,6.098676,6.196286,6.2938967,6.3915067,6.4891167,6.6413884,6.7975645,6.9537406,7.1060123,7.262188,7.605776,7.9493628,8.289046,8.632633,8.976221,9.218294,9.460366,9.702439,9.944512,10.186585,10.053836,9.917182,9.780528,9.647778,9.511124,9.788337,10.065549,10.346666,10.6238785,10.901091,11.611692,12.318389,13.028991,13.739592,14.450192,15.543426,16.640562,17.733795,18.830933,19.924164,19.6001,19.276033,18.95197,18.623999,18.299932,18.22575,18.15547,18.081287,18.011007,17.936825,16.995863,16.058807,15.117846,14.176885,13.235924,13.087557,12.939189,12.786918,12.63855,12.486279,11.943566,11.400854,10.858143,10.319335,9.776623,9.901564,10.03041,10.159255,10.284196,10.413041,11.490656,12.572175,13.653695,14.73131,15.812829,16.761599,17.714273,18.663042,19.611813,20.560583,19.073006,17.589333,16.101755,14.614178,13.1266,13.157836,13.189071,13.224211,13.2554455,13.286681,13.196879,13.103174,13.009468,12.915763,12.825961,12.177831,11.5297,10.881569,10.2334385,9.589212,8.898132,8.207053,7.5159745,6.8287997,6.13772,6.168956,6.2040954,6.2353306,6.266566,6.3017054,5.688714,5.0796275,4.4705405,3.8614538,3.2484627,3.1703746,3.0883822,3.0102942,2.9283018,2.8502135,2.7252727,2.6003318,2.475391,2.35045,2.2255092,2.1044729,1.9834363,1.8663043,1.7452679,1.6242313,1.6008049,1.5734742,1.5500476,1.5266213,1.4992905,1.5110037,1.5266213,1.5383345,1.5500476,1.5617609,1.5851873,1.6086137,1.6281357,1.6515622,1.6749885,1.698415,1.7218413,1.7413634,1.7647898,1.7882162,1.9600099,2.1318035,2.3035975,2.4792955,2.6510892,2.6862288,2.7213683,2.7565079,2.7916477,2.8267872,2.8892577,2.9556324,3.018103,3.084478,3.1508527,3.3734035,3.5959544,3.8185053,4.041056,4.263607,4.5993857,4.93126,5.267039,5.602817,5.938596,6.1611466,6.3836975,6.606249,6.8287997,7.0513506,7.3715115,7.6955767,8.015738,8.339804,8.663869,8.859089,9.054309,9.245625,9.440845,9.636065,9.694631,9.753197,9.811763,9.866425,9.924991,10.354475,10.783959,11.213444,11.6468315,12.076316,12.119265,12.166118,12.209065,12.2559185,12.298867,12.181735,12.064603,11.947471,11.8303385,11.713207,11.697589,11.681972,11.666354,11.650736,11.639023,11.744442,11.845957,11.951375,12.056794,12.162213,12.111456,12.0606985,12.013845,11.963089,11.912332,11.685876,11.45942,11.229061,11.002605,10.77615,10.84643,10.920613,10.990892,11.065076,11.139259,10.916709,10.694158,10.471607,10.249056,10.0265045,9.643873,9.265146,8.886419,8.503788,8.125061,8.03526,7.9454584,7.8556576,7.7658563,7.676055,7.3597984,7.043542,6.7311897,6.4149327,6.098676,6.1299114,6.1611466,6.1884775,6.2197127,6.250948,5.8292727,5.4115014,4.989826,4.5681505,4.1503797,4.2479897,4.3455997,4.4432096,4.5408196,4.6384296,4.4978714,4.357313,4.2167544,4.0761957,3.9356375,3.8965936,3.853645,3.8106966,3.767748,3.7247996,3.7443218,3.7599394,3.775557,3.795079,3.8106966,3.4983444,3.1859922,2.87364,2.5612879,2.2489357,2.7604125,3.2718892,3.7794614,4.290938,4.7985106,4.564246,4.3260775,4.087909,3.8497405,3.611572,3.5178664,3.4241607,3.3265507,3.232845,3.1391394,2.9907722,2.8463092,2.7018464,2.5573835,2.4129205,2.3035975,2.1981785,2.0888553,1.9834363,1.8741131,2.436347,2.2294137,2.0224805,1.815547,1.6086137,1.4016805,1.2181735,1.038571,0.8589685,0.679366,0.4997635,0.40605783,0.30844778,0.21474212,0.12103647,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.042948425,0.058566034,0.078088045,0.093705654,0.113227665,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.19131571,0.21083772,0.22645533,0.24597734,0.26159495,0.26940376,0.27330816,0.27721256,0.28111696,0.28892577,0.3474918,0.40605783,0.46852827,0.5270943,0.58566034,0.62470436,0.6637484,0.698888,0.737932,0.77307165,1.0190489,1.2650263,1.5110037,1.7530766,1.999054,2.514435,3.0298162,3.5451972,4.0605783,4.575959,4.349504,4.126953,3.900498,3.6740425,3.4514916,3.1469483,2.8385005,2.533957,2.2294137,1.9248703,1.7062237,1.4914817,1.2728351,1.0541886,0.8355421,0.6754616,0.5114767,0.3513962,0.18741131,0.023426414,0.058566034,0.08980125,0.12103647,0.15617609,0.18741131,0.15617609,0.12884527,0.09761006,0.06637484,0.039044023,0.031235218,0.023426414,0.015617609,0.0078088045,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.12494087,0.14836729,0.1756981,0.19912452,0.22645533,0.19522011,0.1639849,0.13665408,0.10541886,0.07418364,0.058566034,0.046852827,0.031235218,0.015617609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.031235218,0.06637484,0.09761006,0.12884527,0.1639849,0.27330816,0.38653582,0.4997635,0.61299115,0.7262188,0.78478485,0.8433509,0.9058213,0.96438736,1.0268579,0.8550641,0.6832704,0.5153811,0.3435874,0.1756981,0.14055848,0.10541886,0.07027924,0.03513962,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.011713207,0.015617609,0.019522011,0.023426414,0.046852827,0.06637484,0.08589685,0.10541886,0.12494087,0.10932326,0.093705654,0.078088045,0.06637484,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.039044023,0.078088045,0.12103647,0.16008049,0.19912452,0.3357786,0.46852827,0.60518235,0.7418364,0.8745861,0.98000497,1.0854238,1.1908426,1.2962615,1.4016805,1.6086137,1.8194515,2.0302892,2.241127,2.4480603,2.5690966,2.690133,2.8111696,2.9283018,3.049338,3.0883822,3.1235218,3.1625657,3.2016098,3.2367494,3.3734035,3.506153,3.6428072,3.775557,3.912211,3.8653584,3.8185053,3.7716527,3.7208953,3.6740425,3.6857557,3.6935644,3.7052777,3.7130866,3.7247996,3.7599394,3.795079,3.8302186,3.8653584,3.900498,3.9863946,4.0761957,4.1620927,4.251894,4.337791,4.521298,4.7087092,4.892216,5.0757227,5.263134,4.9546866,4.646239,4.3416953,4.0332475,3.7247996,3.814601,3.9044023,3.9942036,4.084005,4.173806,4.607195,5.040583,5.473972,5.903456,6.336845,6.9615493,7.5862536,8.210958,8.835662,9.464272,10.131924,10.795672,11.4633255,12.130978,12.798631,13.493614,14.184693,14.875772,15.570756,16.261835,16.894348,17.526861,18.159374,18.791887,19.4244,20.021774,20.615244,21.208714,21.806087,22.399555,23.075018,23.750479,24.425941,25.101402,25.776863,26.175114,26.573362,26.975515,27.373764,27.775917,28.025799,28.279585,28.533371,28.783253,29.037039,28.818394,28.603651,28.385004,28.166357,27.951616,27.541653,27.131691,26.72173,26.311768,25.901804,24.78124,23.664581,22.547922,21.431265,20.310701,18.506866,16.703033,14.899199,13.091461,11.287627,10.436467,9.581403,8.730244,7.8790836,7.0240197,6.9342184,6.8405128,6.746807,6.6531014,6.5633,6.715572,6.8678436,7.0201154,7.172387,7.3246584,7.519879,7.715099,7.910319,8.105539,8.300759,8.706817,9.116779,9.522837,9.928895,10.338858,10.569217,10.803481,11.033841,11.268105,11.498465,11.322766,11.143164,10.967466,10.791768,10.612165,10.721489,10.8308115,10.944039,11.053363,11.162686,11.615597,12.068507,12.521418,12.974329,13.423335,14.40334,15.383345,16.36335,17.343355,18.32336,18.249176,18.174992,18.10081,18.026625,17.948538,17.823597,17.694752,17.565907,17.440966,17.31212,16.515621,15.719124,14.918721,14.122223,13.325725,13.376482,13.423335,13.4740925,13.524849,13.575606,13.103174,12.634645,12.166118,11.693685,11.225157,11.248583,11.268105,11.291532,11.314958,11.338385,12.107552,12.8767185,13.645885,14.418958,15.188125,16.398489,17.612759,18.823124,20.037392,21.251661,19.986635,18.725513,17.464392,16.199366,14.938243,14.856251,14.774258,14.688361,14.606369,14.524376,14.618082,14.711788,14.801589,14.895294,14.989,14.161267,13.333533,12.5058,11.678067,10.850334,10.088976,9.331521,8.570163,7.8088045,7.0513506,7.328563,7.60968,7.890797,8.171914,8.449126,7.633106,6.8209906,6.0049706,5.1889505,4.376835,4.2284675,4.084005,3.9395418,3.795079,3.6506162,3.4241607,3.2016098,2.9751544,2.7486992,2.5261483,2.4207294,2.3153105,2.2098918,2.1044729,1.999054,1.9131571,1.8233559,1.737459,1.6515622,1.5617609,1.5617609,1.5617609,1.5617609,1.5617609,1.5617609,1.5656652,1.5656652,1.5695697,1.5734742,1.5734742,1.5773785,1.5812829,1.5812829,1.5851873,1.5890918,1.7140326,1.8428779,1.9717231,2.096664,2.2255092,2.2645533,2.3035975,2.3465457,2.3855898,2.4246337,2.4714866,2.5183394,2.5690966,2.6159496,2.6628022,2.854118,3.0415294,3.232845,3.4241607,3.611572,3.8653584,4.1191444,4.369026,4.6228123,4.8765984,5.0757227,5.278752,5.481781,5.6848097,5.8878384,6.153338,6.4188375,6.6843367,6.9459314,7.211431,7.406651,7.5979667,7.7892823,7.9805984,8.175818,8.203149,8.234385,8.265619,8.296855,8.324185,8.62092,8.913751,9.2104845,9.503315,9.80005,9.780528,9.761005,9.741484,9.718058,9.698535,9.593117,9.483793,9.378374,9.269051,9.163632,9.140205,9.116779,9.093353,9.073831,9.050405,9.108971,9.163632,9.2221985,9.280765,9.339331,9.276859,9.2104845,9.148014,9.085544,9.023073,8.862993,8.706817,8.546737,8.386656,8.226576,8.214863,8.203149,8.19534,8.183627,8.175818,8.011833,7.843944,7.6799593,7.5159745,7.348085,7.1060123,6.860035,6.6140575,6.36808,6.126007,6.04011,5.9542136,5.8683167,5.786324,5.700427,5.4895897,5.278752,5.0718184,4.860981,4.650143,4.6696653,4.689187,4.7087092,4.728231,4.7516575,4.4705405,4.1894236,3.9083066,3.631094,3.349977,3.4007344,3.455396,3.506153,3.5608149,3.611572,3.541293,3.4671092,3.39683,3.3226464,3.2484627,3.2914112,3.3343596,3.377308,3.4202564,3.4632049,3.5451972,3.6271896,3.7091823,3.7911747,3.873167,3.5881457,3.2992198,3.0141985,2.7252727,2.436347,2.9283018,3.416352,3.9083066,4.396357,4.8883114,4.661856,4.4393053,4.21285,3.9863946,3.7638438,3.6701381,3.5764325,3.4866312,3.3929255,3.2992198,3.096191,2.8892577,2.6862288,2.4792955,2.2762666,2.069333,1.8663043,1.6593709,1.456342,1.2494087,2.3114061,2.0654287,1.8194515,1.5695697,1.3235924,1.0737107,0.9097257,0.74574083,0.58175594,0.41386664,0.24988174,0.20302892,0.15617609,0.10932326,0.058566034,0.011713207,0.011713207,0.0078088045,0.0039044023,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.027330816,0.042948425,0.058566034,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.13665408,0.14836729,0.1639849,0.1796025,0.19522011,0.21083772,0.22645533,0.22645533,0.23035973,0.23426414,0.23426414,0.23816854,0.30454338,0.3709182,0.44119745,0.5075723,0.57394713,0.61299115,0.6481308,0.6871748,0.7262188,0.76135844,0.96048295,1.1557031,1.3548276,1.5539521,1.7491722,2.2567444,2.7643168,3.2718892,3.7794614,4.2870336,4.1503797,4.0137253,3.873167,3.736513,3.5998588,3.2367494,2.8697357,2.5066261,2.1396124,1.7765031,1.5227169,1.2689307,1.0190489,0.76526284,0.5114767,0.41386664,0.31235218,0.21083772,0.113227665,0.011713207,0.058566034,0.10932326,0.15617609,0.20302892,0.24988174,0.21083772,0.1717937,0.12884527,0.08980125,0.05075723,0.039044023,0.031235218,0.019522011,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.019522011,0.031235218,0.039044023,0.05075723,0.07418364,0.10151446,0.12494087,0.14836729,0.1756981,0.16008049,0.14446288,0.12884527,0.113227665,0.10151446,0.078088045,0.058566034,0.039044023,0.019522011,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.046852827,0.06637484,0.08980125,0.113227665,0.1639849,0.21083772,0.26159495,0.31235218,0.3631094,0.42948425,0.4958591,0.5661383,0.63251317,0.698888,0.58956474,0.48024148,0.3709182,0.26159495,0.14836729,0.12103647,0.08980125,0.058566034,0.031235218,0.0,0.0,0.0,0.0,0.0,0.0,0.0039044023,0.0039044023,0.0078088045,0.011713207,0.011713207,0.023426414,0.031235218,0.042948425,0.05075723,0.062470436,0.05466163,0.046852827,0.039044023,0.031235218,0.023426414,0.019522011,0.015617609,0.011713207,0.0039044023,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.019522011,0.039044023,0.058566034,0.078088045,0.10151446,0.1678893,0.23426414,0.30063897,0.3709182,0.43729305,0.48805028,0.5427119,0.59346914,0.6481308,0.698888,0.8160201,0.93315214,1.0541886,1.1713207,1.2884527,1.3353056,1.3821584,1.4290112,1.475864,1.5266213,1.5500476,1.5734742,1.6008049,1.6242313,1.6515622,1.7413634,1.8350691,1.9287747,2.018576,2.1122816,2.096664,2.077142,2.0615244,2.0420024,2.0263848,2.1435168,2.260649,2.377781,2.494913,2.612045,2.8424048,3.0727646,3.3031244,3.533484,3.7638438,3.998108,4.2362766,4.474445,4.7126136,4.950782,5.181142,5.4115014,5.6418614,5.8683167,6.098676,5.677001,5.2553253,4.83365,4.40807,3.9863946,3.9942036,4.0020123,4.009821,4.01763,4.025439,4.3338866,4.646239,4.9546866,5.263134,5.575486,6.0752497,6.575013,7.0747766,7.57454,8.074304,8.566258,9.054309,9.546264,10.034314,10.526268,11.275913,12.029464,12.783013,13.536563,14.286208,15.024139,15.758167,16.492195,17.226223,17.964155,18.733322,19.506393,20.279465,21.052536,21.82561,22.47374,23.125774,23.773905,24.425941,25.074072,25.288813,25.499651,25.714394,25.925232,26.136068,26.382046,26.628023,26.874,27.116074,27.362051,27.084839,26.807627,26.530413,26.2532,25.975988,25.694872,25.413754,25.136541,24.855425,24.574308,23.223385,21.868557,20.517633,19.16671,17.811884,16.46096,15.1061325,13.755209,12.404286,11.0494585,10.256865,9.460366,8.663869,7.871275,7.0747766,7.08649,7.094299,7.1060123,7.113821,7.125534,7.3324676,7.5394006,7.746334,7.9532676,8.164105,8.398369,8.632633,8.866898,9.101162,9.339331,9.811763,10.284196,10.756628,11.229061,11.701493,11.924045,12.146595,12.369146,12.591698,12.814248,12.591698,12.373051,12.154405,11.931853,11.713207,11.654641,11.596075,11.541413,11.482847,11.424281,11.619501,11.814721,12.009941,12.205161,12.400381,13.263254,14.130032,14.996809,15.859682,16.72646,16.898252,17.073952,17.24965,17.425346,17.601046,17.417538,17.234032,17.054428,16.870922,16.687416,16.031475,15.37944,14.723501,14.067561,13.411622,13.661504,13.911386,14.161267,14.411149,14.661031,14.2666855,13.868437,13.470188,13.0719385,12.67369,12.591698,12.509705,12.427712,12.34572,12.263727,12.724447,13.181262,13.641981,14.102701,14.56342,16.039284,17.511244,18.987108,20.462973,21.938837,20.900265,19.861694,18.823124,17.788456,16.749886,16.55076,16.355541,16.156416,15.961197,15.762072,16.039284,16.316498,16.59371,16.870922,17.148134,16.140799,15.133463,14.126127,13.118792,12.111456,11.283723,10.452085,9.6243515,8.792714,7.9610763,8.488171,9.019169,9.546264,10.073358,10.600452,9.581403,8.55845,7.5394006,6.520352,5.5013027,5.290465,5.0796275,4.8687897,4.661856,4.4510183,4.123049,3.7989833,3.474918,3.1508527,2.8267872,2.7330816,2.6432803,2.5534792,2.463678,2.3738766,2.2255092,2.0732377,1.9248703,1.7765031,1.6242313,1.6125181,1.6008049,1.5890918,1.5734742,1.5617609,1.5461433,1.5266213,1.5110037,1.4914817,1.475864,1.456342,1.4407244,1.4212024,1.4055848,1.3860629,1.4680552,1.5539521,1.6359446,1.717937,1.7999294,1.8467822,1.8897307,1.9365835,1.979532,2.0263848,2.0537157,2.084951,2.1161861,2.1435168,2.174752,2.330928,2.4910088,2.6471848,2.803361,2.9634414,3.1313305,3.3031244,3.4710135,3.6428072,3.8106966,3.9942036,4.1777105,4.3612175,4.5408196,4.7243266,4.93126,5.138193,5.349031,5.5559645,5.7628975,5.9542136,6.141625,6.3329406,6.524256,6.7116675,6.715572,6.715572,6.719476,6.7233806,6.7233806,6.883461,7.043542,7.2036223,7.363703,7.523783,7.4417906,7.355894,7.269997,7.1841,7.098203,7.000593,6.9068875,6.8092775,6.7116675,6.6140575,6.5828223,6.551587,6.524256,6.493021,6.461786,6.473499,6.481308,6.493021,6.5008297,6.5125427,6.4383593,6.364176,6.2860875,6.211904,6.13772,6.044015,5.9542136,5.860508,5.7668023,5.6730967,5.5832953,5.4895897,5.395884,5.3060827,5.212377,5.1030536,4.997635,4.8883114,4.7828927,4.6735697,4.564246,4.454923,4.3455997,4.2362766,4.123049,4.044961,3.9668727,3.8848803,3.8067923,3.7247996,3.619381,3.513962,3.408543,3.3031244,3.2016098,3.2094188,3.2211318,3.2289407,3.240654,3.2484627,3.1118085,2.97125,2.8306916,2.690133,2.5495746,2.5573835,2.5651922,2.5730011,2.5808098,2.5886188,2.5808098,2.5769055,2.5730011,2.5690966,2.5612879,2.690133,2.8189783,2.9439192,3.0727646,3.2016098,3.3460727,3.49444,3.6428072,3.7911747,3.9356375,3.6740425,3.4124475,3.1508527,2.8892577,2.6237583,3.096191,3.5647192,4.0332475,4.50568,4.9742084,4.7633705,4.548629,4.337791,4.126953,3.912211,3.8224099,3.7326086,3.6428072,3.5530062,3.4632049,3.1977055,2.9322062,2.6667068,2.4012074,2.135708,1.8350691,1.5305257,1.2298868,0.92924774,0.62470436,2.1864653,1.901444,1.6125181,1.3235924,1.038571,0.74964523,0.60127795,0.44900626,0.30063897,0.14836729,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.07418364,0.08589685,0.10151446,0.113227665,0.12494087,0.13665408,0.14836729,0.1639849,0.1756981,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.18741131,0.26159495,0.3357786,0.41386664,0.48805028,0.5622339,0.60127795,0.63641757,0.6754616,0.7106012,0.74964523,0.9019169,1.0502841,1.1986516,1.3509232,1.4992905,1.999054,2.4988174,2.998581,3.4983444,3.998108,3.951255,3.900498,3.8497405,3.7989833,3.7482262,3.3265507,2.900971,2.475391,2.0498111,1.6242313,1.33921,1.0502841,0.76135844,0.47633708,0.18741131,0.14836729,0.113227665,0.07418364,0.039044023,0.0,0.062470436,0.12494087,0.18741131,0.24988174,0.31235218,0.26159495,0.21083772,0.1639849,0.113227665,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.05075723,0.039044023,0.023426414,0.011713207,0.0,0.07418364,0.14836729,0.22645533,0.30063897,0.37482262,0.3240654,0.27330816,0.22645533,0.1756981,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.023426414,0.05075723,0.07418364,0.10151446,0.12494087,0.10151446,0.07418364,0.05075723,0.023426414,0.0,0.011713207,0.023426414,0.039044023,0.05075723,0.062470436,0.113227665,0.1639849,0.21083772,0.26159495,0.31235218,0.3240654,0.3357786,0.3513962,0.3631094,0.37482262,0.60127795,0.8238289,1.0502841,1.2767396,1.4992905,1.9248703,2.35045,2.77603,3.2016098,3.6232853,4.0137253,4.4002614,4.786797,5.173333,5.563773,5.8370814,6.114294,6.387602,6.66091,6.9381227,6.3993154,5.8644123,5.3256044,4.786797,4.251894,4.173806,4.0996222,4.025439,3.951255,3.873167,4.0605783,4.251894,4.4393053,4.6267166,4.814128,5.1889505,5.563773,5.938596,6.3134184,6.688241,7.000593,7.3129454,7.6252975,7.9376497,8.250002,9.062118,9.874233,10.686349,11.498465,12.31058,13.150026,13.985569,14.825015,15.664462,16.500004,17.448774,18.401447,19.350218,20.298986,21.251661,21.876366,22.50107,23.125774,23.750479,24.375183,24.39861,24.425941,24.449368,24.476698,24.500124,24.738293,24.976461,25.210726,25.448895,25.687063,25.351284,25.0116,24.675823,24.33614,24.00036,23.84809,23.699722,23.551353,23.399082,23.250715,21.661623,20.076437,18.487345,16.898252,15.313066,14.411149,13.513136,12.611219,11.713207,10.81129,10.073358,9.339331,8.601398,7.8634663,7.125534,7.238762,7.348085,7.461313,7.57454,7.687768,7.9493628,8.210958,8.476458,8.738052,8.999647,9.276859,9.550168,9.823476,10.100689,10.373997,10.912805,11.4516115,11.986515,12.525322,13.06413,13.274967,13.4858055,13.700547,13.911386,14.126127,13.860628,13.599033,13.337439,13.075843,12.814248,12.587793,12.361338,12.138786,11.912332,11.685876,11.623405,11.560935,11.498465,11.435994,11.373524,12.123169,12.8767185,13.626364,14.376009,15.125654,15.551234,15.976814,16.398489,16.82407,17.24965,17.01148,16.773312,16.539047,16.300879,16.062712,15.551234,15.035853,14.524376,14.012899,13.501423,13.950429,14.399435,14.848442,15.3013525,15.750359,15.426293,15.098324,14.774258,14.450192,14.126127,13.938716,13.751305,13.563893,13.376482,13.189071,13.337439,13.4858055,13.638077,13.786445,13.938716,15.676175,17.413633,19.151093,20.888552,22.62601,21.813896,21.00178,20.18576,19.373644,18.56153,18.249176,17.936825,17.624472,17.31212,16.999767,17.464392,17.92511,18.38583,18.850454,19.311174,18.124235,16.937298,15.750359,14.56342,13.376482,12.4745655,11.576552,10.674636,9.776623,8.874706,9.651682,10.424754,11.20173,11.974802,12.751778,11.525795,10.299813,9.073831,7.8517528,6.6257706,6.348558,6.0752497,5.801942,5.5247293,5.251421,4.825841,4.4002614,3.9746814,3.5491016,3.1235218,3.049338,2.9751544,2.900971,2.8267872,2.7486992,2.5378613,2.3231194,2.1122816,1.901444,1.6867018,1.6632754,1.6359446,1.6125181,1.5890918,1.5617609,1.5266213,1.4875772,1.4485333,1.4133936,1.3743496,1.33921,1.3001659,1.261122,1.2259823,1.1869383,1.2259823,1.261122,1.3001659,1.33921,1.3743496,1.4251068,1.475864,1.5266213,1.5734742,1.6242313,1.6359446,1.6515622,1.6632754,1.6749885,1.6867018,1.8116426,1.9365835,2.0615244,2.1864653,2.3114061,2.4012074,2.4871042,2.5769055,2.6628022,2.7486992,2.912684,3.076669,3.2367494,3.4007344,3.5608149,3.7130866,3.8614538,4.0137253,4.1620927,4.3143644,4.5017757,4.689187,4.8765984,5.0640097,5.251421,5.22409,5.2006636,5.173333,5.1499066,5.12648,5.1499066,5.173333,5.2006636,5.22409,5.251421,5.099149,4.950782,4.7985106,4.650143,4.5017757,4.4119744,4.3260775,4.2362766,4.1503797,4.0605783,4.025439,3.9863946,3.951255,3.912211,3.873167,3.8380275,3.7989833,3.7638438,3.7247996,3.6857557,3.5998588,3.513962,3.4241607,3.338264,3.2484627,3.2250361,3.2016098,3.174279,3.1508527,3.1235218,2.951728,2.77603,2.6003318,2.4246337,2.2489357,2.1981785,2.1513257,2.1005683,2.0498111,1.999054,2.0263848,2.0498111,2.0732377,2.1005683,2.1239948,2.0498111,1.9756275,1.901444,1.8233559,1.7491722,1.7491722,1.7491722,1.7491722,1.7491722,1.7491722,1.7491722,1.7491722,1.7491722,1.7491722,1.7491722,1.7491722,1.7491722,1.7491722,1.7491722,1.7491722,1.7140326,1.6749885,1.6359446,1.6008049,1.5617609,1.6242313,1.6867018,1.7491722,1.8116426,1.8741131,2.0888553,2.2996929,2.514435,2.7252727,2.9361105,3.1508527,3.3616903,3.5764325,3.78727,3.998108,3.7638438,3.5256753,3.2875066,3.049338,2.8111696,3.2640803,3.7130866,4.1620927,4.6110992,5.0640097,4.860981,4.661856,4.462732,4.263607,4.0605783,3.9746814,3.8887846,3.7989833,3.7130866,3.6232853,3.2992198,2.9751544,2.6510892,2.3231194,1.999054,1.6008049,1.1986516,0.80040246,0.39824903,0.0;
 } 
